
module SNPS_CLOCK_GATE_HIGH_avr_pooling_fsm ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKGATETST_X1 latch ( .CK(CLK), .E(EN), .SE(TE), .GCK(ENCLK) );
endmodule


module avr_pooling_unrolled ( clk, rst_fsm, start, done, en, size_1, size_2, 
        pool_sel, d_0, d_1, d_2, d_3, d_4, d_5, d_6, d_7, o_pool_1, o_pool_2, 
        o_pool_3, o_pool_4 );
  input [4:0] size_1;
  input [4:0] size_2;
  input [15:0] d_0;
  input [15:0] d_1;
  input [15:0] d_2;
  input [15:0] d_3;
  input [15:0] d_4;
  input [15:0] d_5;
  input [15:0] d_6;
  input [15:0] d_7;
  output [15:0] o_pool_1;
  output [15:0] o_pool_2;
  output [15:0] o_pool_3;
  output [15:0] o_pool_4;
  input clk, rst_fsm, start, done, en, pool_sel;
  wire   \pool/ld_h , \pool/rst_cnt_r , \pool/rst_cnt_c , \pool/tc ,
         \pool/en_cnt , \pool/rst_cnt , \pool/sync_clr , \pool/sel ,
         \pool/pool/pe_b_o_data[0][43] , \pool/pool/pe_b_o_data[0][42] ,
         \pool/pool/pe_b_o_data[0][41] , \pool/pool/pe_b_o_data[0][40] ,
         \pool/pool/pe_b_o_data[0][39] , \pool/pool/pe_b_o_data[0][38] ,
         \pool/pool/pe_b_o_data[0][37] , \pool/pool/pe_b_o_data[0][36] ,
         \pool/pool/pe_b_o_data[0][35] , \pool/pool/pe_b_o_data[0][34] ,
         \pool/pool/pe_b_o_data[0][33] , \pool/pool/pe_b_o_data[0][32] ,
         \pool/pool/pe_b_o_data[0][31] , \pool/pool/pe_b_o_data[0][30] ,
         \pool/pool/pe_b_o_data[0][29] , \pool/pool/pe_b_o_data[0][28] ,
         \pool/pool/pe_b_o_data[0][27] , \pool/pool/pe_b_o_data[0][26] ,
         \pool/pool/pe_b_o_data[0][25] , \pool/pool/pe_b_o_data[0][24] ,
         \pool/pool/pe_b_o_data[0][23] , \pool/pool/pe_b_o_data[0][22] ,
         \pool/pool/pe_b_o_data[0][21] , \pool/pool/pe_b_o_data[0][20] ,
         \pool/pool/pe_b_o_data[0][19] , \pool/pool/pe_b_o_data[0][18] ,
         \pool/pool/pe_b_o_data[0][17] , \pool/pool/pe_b_o_data[0][16] ,
         \pool/pool/pe_b_o_data[0][15] , \pool/pool/pe_b_o_data[0][14] ,
         \pool/pool/pe_b_o_data[0][13] , \pool/pool/pe_b_o_data[0][12] ,
         \pool/pool/pe_b_o_data[0][11] , \pool/pool/pe_b_o_data[0][10] ,
         \pool/pool/pe_b_o_data[0][9] , \pool/pool/pe_b_o_data[0][8] ,
         \pool/pool/pe_b_o_data[0][7] , \pool/pool/pe_b_o_data[0][6] ,
         \pool/pool/pe_b_o_data[0][5] , \pool/pool/pe_b_o_data[0][4] ,
         \pool/pool/pe_b_o_data[0][3] , \pool/pool/pe_b_o_data[0][2] ,
         \pool/pool/pe_b_o_data[0][1] , \pool/pool/pe_b_o_data[0][0] ,
         \pool/pool/pe_b_o_data[1][43] , \pool/pool/pe_b_o_data[1][42] ,
         \pool/pool/pe_b_o_data[1][41] , \pool/pool/pe_b_o_data[1][40] ,
         \pool/pool/pe_b_o_data[1][39] , \pool/pool/pe_b_o_data[1][38] ,
         \pool/pool/pe_b_o_data[1][37] , \pool/pool/pe_b_o_data[1][36] ,
         \pool/pool/pe_b_o_data[1][35] , \pool/pool/pe_b_o_data[1][34] ,
         \pool/pool/pe_b_o_data[1][33] , \pool/pool/pe_b_o_data[1][32] ,
         \pool/pool/pe_b_o_data[1][31] , \pool/pool/pe_b_o_data[1][30] ,
         \pool/pool/pe_b_o_data[1][29] , \pool/pool/pe_b_o_data[1][28] ,
         \pool/pool/pe_b_o_data[1][27] , \pool/pool/pe_b_o_data[1][26] ,
         \pool/pool/pe_b_o_data[1][25] , \pool/pool/pe_b_o_data[1][24] ,
         \pool/pool/pe_b_o_data[1][23] , \pool/pool/pe_b_o_data[1][22] ,
         \pool/pool/pe_b_o_data[1][21] , \pool/pool/pe_b_o_data[1][20] ,
         \pool/pool/pe_b_o_data[1][19] , \pool/pool/pe_b_o_data[1][18] ,
         \pool/pool/pe_b_o_data[1][17] , \pool/pool/pe_b_o_data[1][16] ,
         \pool/pool/pe_b_o_data[1][15] , \pool/pool/pe_b_o_data[1][14] ,
         \pool/pool/pe_b_o_data[1][13] , \pool/pool/pe_b_o_data[1][12] ,
         \pool/pool/pe_b_o_data[1][11] , \pool/pool/pe_b_o_data[1][10] ,
         \pool/pool/pe_b_o_data[1][9] , \pool/pool/pe_b_o_data[1][8] ,
         \pool/pool/pe_b_o_data[1][7] , \pool/pool/pe_b_o_data[1][6] ,
         \pool/pool/pe_b_o_data[1][5] , \pool/pool/pe_b_o_data[1][4] ,
         \pool/pool/pe_b_o_data[1][3] , \pool/pool/pe_b_o_data[1][2] ,
         \pool/pool/pe_b_o_data[1][1] , \pool/pool/pe_b_o_data[1][0] ,
         \pool/pool/pe_b_o_data[2][43] , \pool/pool/pe_b_o_data[2][42] ,
         \pool/pool/pe_b_o_data[2][41] , \pool/pool/pe_b_o_data[2][40] ,
         \pool/pool/pe_b_o_data[2][39] , \pool/pool/pe_b_o_data[2][38] ,
         \pool/pool/pe_b_o_data[2][37] , \pool/pool/pe_b_o_data[2][36] ,
         \pool/pool/pe_b_o_data[2][35] , \pool/pool/pe_b_o_data[2][34] ,
         \pool/pool/pe_b_o_data[2][33] , \pool/pool/pe_b_o_data[2][32] ,
         \pool/pool/pe_b_o_data[2][31] , \pool/pool/pe_b_o_data[2][30] ,
         \pool/pool/pe_b_o_data[2][29] , \pool/pool/pe_b_o_data[2][28] ,
         \pool/pool/pe_b_o_data[2][27] , \pool/pool/pe_b_o_data[2][26] ,
         \pool/pool/pe_b_o_data[2][25] , \pool/pool/pe_b_o_data[2][24] ,
         \pool/pool/pe_b_o_data[2][23] , \pool/pool/pe_b_o_data[2][22] ,
         \pool/pool/pe_b_o_data[2][21] , \pool/pool/pe_b_o_data[2][20] ,
         \pool/pool/pe_b_o_data[2][19] , \pool/pool/pe_b_o_data[2][18] ,
         \pool/pool/pe_b_o_data[2][17] , \pool/pool/pe_b_o_data[2][16] ,
         \pool/pool/pe_b_o_data[2][15] , \pool/pool/pe_b_o_data[2][14] ,
         \pool/pool/pe_b_o_data[2][13] , \pool/pool/pe_b_o_data[2][12] ,
         \pool/pool/pe_b_o_data[2][11] , \pool/pool/pe_b_o_data[2][10] ,
         \pool/pool/pe_b_o_data[2][9] , \pool/pool/pe_b_o_data[2][8] ,
         \pool/pool/pe_b_o_data[2][7] , \pool/pool/pe_b_o_data[2][6] ,
         \pool/pool/pe_b_o_data[2][5] , \pool/pool/pe_b_o_data[2][4] ,
         \pool/pool/pe_b_o_data[2][3] , \pool/pool/pe_b_o_data[2][2] ,
         \pool/pool/pe_b_o_data[2][1] , \pool/pool/pe_b_o_data[2][0] ,
         \pool/pool/pe_b_o_data[3][43] , \pool/pool/pe_b_o_data[3][42] ,
         \pool/pool/pe_b_o_data[3][41] , \pool/pool/pe_b_o_data[3][40] ,
         \pool/pool/pe_b_o_data[3][39] , \pool/pool/pe_b_o_data[3][38] ,
         \pool/pool/pe_b_o_data[3][37] , \pool/pool/pe_b_o_data[3][36] ,
         \pool/pool/pe_b_o_data[3][35] , \pool/pool/pe_b_o_data[3][34] ,
         \pool/pool/pe_b_o_data[3][33] , \pool/pool/pe_b_o_data[3][32] ,
         \pool/pool/pe_b_o_data[3][31] , \pool/pool/pe_b_o_data[3][30] ,
         \pool/pool/pe_b_o_data[3][29] , \pool/pool/pe_b_o_data[3][28] ,
         \pool/pool/pe_b_o_data[3][27] , \pool/pool/pe_b_o_data[3][26] ,
         \pool/pool/pe_b_o_data[3][25] , \pool/pool/pe_b_o_data[3][24] ,
         \pool/pool/pe_b_o_data[3][23] , \pool/pool/pe_b_o_data[3][22] ,
         \pool/pool/pe_b_o_data[3][21] , \pool/pool/pe_b_o_data[3][20] ,
         \pool/pool/pe_b_o_data[3][19] , \pool/pool/pe_b_o_data[3][18] ,
         \pool/pool/pe_b_o_data[3][17] , \pool/pool/pe_b_o_data[3][16] ,
         \pool/pool/pe_b_o_data[3][15] , \pool/pool/pe_b_o_data[3][14] ,
         \pool/pool/pe_b_o_data[3][13] , \pool/pool/pe_b_o_data[3][12] ,
         \pool/pool/pe_b_o_data[3][11] , \pool/pool/pe_b_o_data[3][10] ,
         \pool/pool/pe_b_o_data[3][9] , \pool/pool/pe_b_o_data[3][8] ,
         \pool/pool/pe_b_o_data[3][7] , \pool/pool/pe_b_o_data[3][6] ,
         \pool/pool/pe_b_o_data[3][5] , \pool/pool/pe_b_o_data[3][4] ,
         \pool/pool/pe_b_o_data[3][3] , \pool/pool/pe_b_o_data[3][2] ,
         \pool/pool/pe_b_o_data[3][1] , \pool/pool/pe_b_o_data[3][0] ,
         \pool/pool/pe_b_i_data[0][15] , \pool/pool/pe_b_i_data[0][14] ,
         \pool/pool/pe_b_i_data[0][13] , \pool/pool/pe_b_i_data[0][12] ,
         \pool/pool/pe_b_i_data[0][11] , \pool/pool/pe_b_i_data[0][10] ,
         \pool/pool/pe_b_i_data[0][9] , \pool/pool/pe_b_i_data[0][8] ,
         \pool/pool/pe_b_i_data[0][7] , \pool/pool/pe_b_i_data[0][6] ,
         \pool/pool/pe_b_i_data[0][5] , \pool/pool/pe_b_i_data[0][4] ,
         \pool/pool/pe_b_i_data[0][3] , \pool/pool/pe_b_i_data[0][2] ,
         \pool/pool/pe_b_i_data[0][1] , \pool/pool/pe_b_i_data[0][0] ,
         \pool/pool/pe_b_i_data[1][15] , \pool/pool/pe_b_i_data[1][14] ,
         \pool/pool/pe_b_i_data[1][13] , \pool/pool/pe_b_i_data[1][12] ,
         \pool/pool/pe_b_i_data[1][11] , \pool/pool/pe_b_i_data[1][10] ,
         \pool/pool/pe_b_i_data[1][9] , \pool/pool/pe_b_i_data[1][8] ,
         \pool/pool/pe_b_i_data[1][7] , \pool/pool/pe_b_i_data[1][6] ,
         \pool/pool/pe_b_i_data[1][5] , \pool/pool/pe_b_i_data[1][4] ,
         \pool/pool/pe_b_i_data[1][3] , \pool/pool/pe_b_i_data[1][2] ,
         \pool/pool/pe_b_i_data[1][1] , \pool/pool/pe_b_i_data[1][0] ,
         \pool/pool/pe_b_i_data[2][15] , \pool/pool/pe_b_i_data[2][14] ,
         \pool/pool/pe_b_i_data[2][13] , \pool/pool/pe_b_i_data[2][12] ,
         \pool/pool/pe_b_i_data[2][11] , \pool/pool/pe_b_i_data[2][10] ,
         \pool/pool/pe_b_i_data[2][9] , \pool/pool/pe_b_i_data[2][8] ,
         \pool/pool/pe_b_i_data[2][7] , \pool/pool/pe_b_i_data[2][6] ,
         \pool/pool/pe_b_i_data[2][5] , \pool/pool/pe_b_i_data[2][4] ,
         \pool/pool/pe_b_i_data[2][3] , \pool/pool/pe_b_i_data[2][2] ,
         \pool/pool/pe_b_i_data[2][1] , \pool/pool/pe_b_i_data[2][0] ,
         \pool/pool/pe_b_i_data[3][15] , \pool/pool/pe_b_i_data[3][14] ,
         \pool/pool/pe_b_i_data[3][13] , \pool/pool/pe_b_i_data[3][12] ,
         \pool/pool/pe_b_i_data[3][11] , \pool/pool/pe_b_i_data[3][10] ,
         \pool/pool/pe_b_i_data[3][9] , \pool/pool/pe_b_i_data[3][8] ,
         \pool/pool/pe_b_i_data[3][7] , \pool/pool/pe_b_i_data[3][6] ,
         \pool/pool/pe_b_i_data[3][5] , \pool/pool/pe_b_i_data[3][4] ,
         \pool/pool/pe_b_i_data[3][3] , \pool/pool/pe_b_i_data[3][2] ,
         \pool/pool/pe_b_i_data[3][1] , \pool/pool/pe_b_i_data[3][0] ,
         \pool/pool/cnt[0] , \pool/pool/cnt[1] ,
         \pool/pool/interface/mux_0/n9 , \pool/pool/interface/mux_0/n8 ,
         \pool/pool/interface/mux_0/n7 , \pool/pool/interface/mux_0/n6 ,
         \pool/pool/interface/mux_0/n5 , \pool/pool/interface/mux_0/n4 ,
         \pool/pool/interface/mux_0/n3 , \pool/pool/interface/mux_0/n2 ,
         \pool/pool/interface/mux_0/n1 , \pool/pool/interface/mux_0/n33 ,
         \pool/pool/interface/mux_0/n32 , \pool/pool/interface/mux_0/n31 ,
         \pool/pool/interface/mux_0/n30 , \pool/pool/interface/mux_0/n29 ,
         \pool/pool/interface/mux_0/n28 , \pool/pool/interface/mux_0/n27 ,
         \pool/pool/interface/mux_0/n26 , \pool/pool/interface/mux_0/n25 ,
         \pool/pool/interface/mux_0/n24 , \pool/pool/interface/mux_0/n23 ,
         \pool/pool/interface/mux_0/n22 , \pool/pool/interface/mux_0/n21 ,
         \pool/pool/interface/mux_0/n20 , \pool/pool/interface/mux_0/n19 ,
         \pool/pool/interface/mux_0/n18 , \pool/pool/interface/mux_1/n33 ,
         \pool/pool/interface/mux_1/n32 , \pool/pool/interface/mux_1/n31 ,
         \pool/pool/interface/mux_1/n30 , \pool/pool/interface/mux_1/n29 ,
         \pool/pool/interface/mux_1/n28 , \pool/pool/interface/mux_1/n27 ,
         \pool/pool/interface/mux_1/n26 , \pool/pool/interface/mux_1/n17 ,
         \pool/pool/interface/mux_1/n16 , \pool/pool/interface/mux_1/n15 ,
         \pool/pool/interface/mux_1/n14 , \pool/pool/interface/mux_1/n13 ,
         \pool/pool/interface/mux_1/n12 , \pool/pool/interface/mux_1/n11 ,
         \pool/pool/interface/mux_1/n10 , \pool/pool/interface/mux_1/n9 ,
         \pool/pool/interface/mux_1/n8 , \pool/pool/interface/mux_1/n7 ,
         \pool/pool/interface/mux_1/n6 , \pool/pool/interface/mux_1/n5 ,
         \pool/pool/interface/mux_1/n4 , \pool/pool/interface/mux_1/n3 ,
         \pool/pool/interface/mux_1/n2 , \pool/pool/interface/mux_1/n1 ,
         \pool/pool/interface/mux_2/n33 , \pool/pool/interface/mux_2/n32 ,
         \pool/pool/interface/mux_2/n31 , \pool/pool/interface/mux_2/n30 ,
         \pool/pool/interface/mux_2/n29 , \pool/pool/interface/mux_2/n28 ,
         \pool/pool/interface/mux_2/n27 , \pool/pool/interface/mux_2/n26 ,
         \pool/pool/interface/mux_2/n17 , \pool/pool/interface/mux_2/n16 ,
         \pool/pool/interface/mux_2/n15 , \pool/pool/interface/mux_2/n14 ,
         \pool/pool/interface/mux_2/n13 , \pool/pool/interface/mux_2/n12 ,
         \pool/pool/interface/mux_2/n11 , \pool/pool/interface/mux_2/n10 ,
         \pool/pool/interface/mux_2/n9 , \pool/pool/interface/mux_2/n8 ,
         \pool/pool/interface/mux_2/n7 , \pool/pool/interface/mux_2/n6 ,
         \pool/pool/interface/mux_2/n5 , \pool/pool/interface/mux_2/n4 ,
         \pool/pool/interface/mux_2/n3 , \pool/pool/interface/mux_2/n2 ,
         \pool/pool/interface/mux_2/n1 , \pool/pool/interface/mux_3/n33 ,
         \pool/pool/interface/mux_3/n32 , \pool/pool/interface/mux_3/n31 ,
         \pool/pool/interface/mux_3/n30 , \pool/pool/interface/mux_3/n29 ,
         \pool/pool/interface/mux_3/n28 , \pool/pool/interface/mux_3/n27 ,
         \pool/pool/interface/mux_3/n26 , \pool/pool/interface/mux_3/n17 ,
         \pool/pool/interface/mux_3/n16 , \pool/pool/interface/mux_3/n15 ,
         \pool/pool/interface/mux_3/n14 , \pool/pool/interface/mux_3/n13 ,
         \pool/pool/interface/mux_3/n12 , \pool/pool/interface/mux_3/n11 ,
         \pool/pool/interface/mux_3/n10 , \pool/pool/interface/mux_3/n9 ,
         \pool/pool/interface/mux_3/n8 , \pool/pool/interface/mux_3/n7 ,
         \pool/pool/interface/mux_3/n6 , \pool/pool/interface/mux_3/n5 ,
         \pool/pool/interface/mux_3/n4 , \pool/pool/interface/mux_3/n3 ,
         \pool/pool/interface/mux_3/n2 , \pool/pool/interface/mux_3/n1 ,
         \pool/pool/pe_b/n7 , \pool/pool/pe_b/n6 , \pool/pool/pe_b/n5 ,
         \pool/pool/pe_b/n4 , \pool/pool/pe_b/n3 , \pool/pool/pe_b/n2 ,
         \pool/pool/pe_b/n1 , \pool/pool/pe_b/int_pe_en[0][0] ,
         \pool/pool/pe_b/int_pe_en[0][1] , \pool/pool/pe_b/int_pe_en[0][2] ,
         \pool/pool/pe_b/int_pe_en[0][3] , \pool/pool/pe_b/int_pe_en[1][0] ,
         \pool/pool/pe_b/int_pe_en[1][1] , \pool/pool/pe_b/int_pe_en[1][2] ,
         \pool/pool/pe_b/int_pe_en[1][3] , \pool/pool/pe_b/int_pe_en[2][0] ,
         \pool/pool/pe_b/int_pe_en[2][1] , \pool/pool/pe_b/int_pe_en[2][2] ,
         \pool/pool/pe_b/int_pe_en[2][3] , \pool/pool/pe_b/int_pe_en[3][0] ,
         \pool/pool/pe_b/int_pe_en[3][1] , \pool/pool/pe_b/int_pe_en[3][2] ,
         \pool/pool/pe_b/int_pe_en[3][3] , \pool/pool/pe_b/peij_0_0/n16 ,
         \pool/pool/pe_b/peij_0_0/n12 , \pool/pool/pe_b/peij_0_0/n11 ,
         \pool/pool/pe_b/peij_0_0/n10 , \pool/pool/pe_b/peij_0_0/n9 ,
         \pool/pool/pe_b/peij_0_0/n8 , \pool/pool/pe_b/peij_0_0/n7 ,
         \pool/pool/pe_b/peij_0_0/n6 , \pool/pool/pe_b/peij_0_0/n5 ,
         \pool/pool/pe_b/peij_0_0/n4 , \pool/pool/pe_b/peij_0_0/n3 ,
         \pool/pool/pe_b/peij_0_0/n2 , \pool/pool/pe_b/peij_0_0/n1 ,
         \pool/pool/pe_b/peij_0_0/n15 , \pool/pool/pe_b/peij_0_0/n14 ,
         \pool/pool/pe_b/peij_0_0/N36 , \pool/pool/pe_b/peij_0_0/N35 ,
         \pool/pool/pe_b/peij_0_0/N34 , \pool/pool/pe_b/peij_0_0/N33 ,
         \pool/pool/pe_b/peij_0_0/q_k , \pool/pool/pe_b/peij_0_0/sgnext_10 ,
         \pool/pool/pe_b/peij_0_0/add/c_out ,
         \pool/pool/pe_b/peij_0_0/add/fai_0/n3 ,
         \pool/pool/pe_b/peij_0_0/add/fai_0/n2 ,
         \pool/pool/pe_b/peij_0_0/add/fai_1/n3 ,
         \pool/pool/pe_b/peij_0_0/add/fai_1/n1 ,
         \pool/pool/pe_b/peij_0_0/add/fai_2/n3 ,
         \pool/pool/pe_b/peij_0_0/add/fai_2/n1 ,
         \pool/pool/pe_b/peij_0_0/add/fai_3/n3 ,
         \pool/pool/pe_b/peij_0_0/add/fai_3/n1 ,
         \pool/pool/pe_b/peij_0_0/add/fai_4/n3 ,
         \pool/pool/pe_b/peij_0_0/add/fai_4/n1 ,
         \pool/pool/pe_b/peij_0_0/add/fai_5/n3 ,
         \pool/pool/pe_b/peij_0_0/add/fai_5/n1 ,
         \pool/pool/pe_b/peij_0_0/add/fai_6/n3 ,
         \pool/pool/pe_b/peij_0_0/add/fai_6/n1 ,
         \pool/pool/pe_b/peij_0_0/add/fai_7/n3 ,
         \pool/pool/pe_b/peij_0_0/add/fai_7/n1 ,
         \pool/pool/pe_b/peij_0_0/add/fai_8/n3 ,
         \pool/pool/pe_b/peij_0_0/add/fai_8/n1 ,
         \pool/pool/pe_b/peij_0_0/add/fai_9/n3 ,
         \pool/pool/pe_b/peij_0_0/add/fai_9/n1 ,
         \pool/pool/pe_b/peij_0_0/add/fai_10/n3 ,
         \pool/pool/pe_b/peij_0_0/add/fai_10/n1 ,
         \pool/pool/pe_b/peij_0_1/n18 , \pool/pool/pe_b/peij_0_1/n17 ,
         \pool/pool/pe_b/peij_0_1/n16 , \pool/pool/pe_b/peij_0_1/n12 ,
         \pool/pool/pe_b/peij_0_1/n11 , \pool/pool/pe_b/peij_0_1/n10 ,
         \pool/pool/pe_b/peij_0_1/n9 , \pool/pool/pe_b/peij_0_1/n8 ,
         \pool/pool/pe_b/peij_0_1/n7 , \pool/pool/pe_b/peij_0_1/n6 ,
         \pool/pool/pe_b/peij_0_1/n5 , \pool/pool/pe_b/peij_0_1/n4 ,
         \pool/pool/pe_b/peij_0_1/n3 , \pool/pool/pe_b/peij_0_1/n2 ,
         \pool/pool/pe_b/peij_0_1/n1 , \pool/pool/pe_b/peij_0_1/N36 ,
         \pool/pool/pe_b/peij_0_1/N35 , \pool/pool/pe_b/peij_0_1/N34 ,
         \pool/pool/pe_b/peij_0_1/N33 , \pool/pool/pe_b/peij_0_1/q_k ,
         \pool/pool/pe_b/peij_0_1/sgnext_10 ,
         \pool/pool/pe_b/peij_0_1/add/c_out ,
         \pool/pool/pe_b/peij_0_1/add/fai_0/n3 ,
         \pool/pool/pe_b/peij_0_1/add/fai_0/n1 ,
         \pool/pool/pe_b/peij_0_1/add/fai_1/n3 ,
         \pool/pool/pe_b/peij_0_1/add/fai_1/n1 ,
         \pool/pool/pe_b/peij_0_1/add/fai_2/n3 ,
         \pool/pool/pe_b/peij_0_1/add/fai_2/n1 ,
         \pool/pool/pe_b/peij_0_1/add/fai_3/n3 ,
         \pool/pool/pe_b/peij_0_1/add/fai_3/n1 ,
         \pool/pool/pe_b/peij_0_1/add/fai_4/n3 ,
         \pool/pool/pe_b/peij_0_1/add/fai_4/n1 ,
         \pool/pool/pe_b/peij_0_1/add/fai_5/n3 ,
         \pool/pool/pe_b/peij_0_1/add/fai_5/n1 ,
         \pool/pool/pe_b/peij_0_1/add/fai_6/n3 ,
         \pool/pool/pe_b/peij_0_1/add/fai_6/n1 ,
         \pool/pool/pe_b/peij_0_1/add/fai_7/n3 ,
         \pool/pool/pe_b/peij_0_1/add/fai_7/n1 ,
         \pool/pool/pe_b/peij_0_1/add/fai_8/n3 ,
         \pool/pool/pe_b/peij_0_1/add/fai_8/n1 ,
         \pool/pool/pe_b/peij_0_1/add/fai_9/n3 ,
         \pool/pool/pe_b/peij_0_1/add/fai_9/n1 ,
         \pool/pool/pe_b/peij_0_1/add/fai_10/n3 ,
         \pool/pool/pe_b/peij_0_1/add/fai_10/n1 ,
         \pool/pool/pe_b/peij_0_2/n18 , \pool/pool/pe_b/peij_0_2/n17 ,
         \pool/pool/pe_b/peij_0_2/n16 , \pool/pool/pe_b/peij_0_2/n12 ,
         \pool/pool/pe_b/peij_0_2/n11 , \pool/pool/pe_b/peij_0_2/n10 ,
         \pool/pool/pe_b/peij_0_2/n9 , \pool/pool/pe_b/peij_0_2/n8 ,
         \pool/pool/pe_b/peij_0_2/n7 , \pool/pool/pe_b/peij_0_2/n6 ,
         \pool/pool/pe_b/peij_0_2/n5 , \pool/pool/pe_b/peij_0_2/n4 ,
         \pool/pool/pe_b/peij_0_2/n3 , \pool/pool/pe_b/peij_0_2/n2 ,
         \pool/pool/pe_b/peij_0_2/n1 , \pool/pool/pe_b/peij_0_2/N36 ,
         \pool/pool/pe_b/peij_0_2/N35 , \pool/pool/pe_b/peij_0_2/N34 ,
         \pool/pool/pe_b/peij_0_2/N33 , \pool/pool/pe_b/peij_0_2/q_k ,
         \pool/pool/pe_b/peij_0_2/sgnext_10 ,
         \pool/pool/pe_b/peij_0_2/add/c_out ,
         \pool/pool/pe_b/peij_0_2/add/fai_0/n3 ,
         \pool/pool/pe_b/peij_0_2/add/fai_0/n1 ,
         \pool/pool/pe_b/peij_0_2/add/fai_1/n3 ,
         \pool/pool/pe_b/peij_0_2/add/fai_1/n1 ,
         \pool/pool/pe_b/peij_0_2/add/fai_2/n3 ,
         \pool/pool/pe_b/peij_0_2/add/fai_2/n1 ,
         \pool/pool/pe_b/peij_0_2/add/fai_3/n3 ,
         \pool/pool/pe_b/peij_0_2/add/fai_3/n1 ,
         \pool/pool/pe_b/peij_0_2/add/fai_4/n3 ,
         \pool/pool/pe_b/peij_0_2/add/fai_4/n1 ,
         \pool/pool/pe_b/peij_0_2/add/fai_5/n3 ,
         \pool/pool/pe_b/peij_0_2/add/fai_5/n1 ,
         \pool/pool/pe_b/peij_0_2/add/fai_6/n3 ,
         \pool/pool/pe_b/peij_0_2/add/fai_6/n1 ,
         \pool/pool/pe_b/peij_0_2/add/fai_7/n3 ,
         \pool/pool/pe_b/peij_0_2/add/fai_7/n1 ,
         \pool/pool/pe_b/peij_0_2/add/fai_8/n3 ,
         \pool/pool/pe_b/peij_0_2/add/fai_8/n1 ,
         \pool/pool/pe_b/peij_0_2/add/fai_9/n3 ,
         \pool/pool/pe_b/peij_0_2/add/fai_9/n1 ,
         \pool/pool/pe_b/peij_0_2/add/fai_10/n3 ,
         \pool/pool/pe_b/peij_0_2/add/fai_10/n1 ,
         \pool/pool/pe_b/peij_0_3/n18 , \pool/pool/pe_b/peij_0_3/n17 ,
         \pool/pool/pe_b/peij_0_3/n16 , \pool/pool/pe_b/peij_0_3/n12 ,
         \pool/pool/pe_b/peij_0_3/n11 , \pool/pool/pe_b/peij_0_3/n10 ,
         \pool/pool/pe_b/peij_0_3/n9 , \pool/pool/pe_b/peij_0_3/n8 ,
         \pool/pool/pe_b/peij_0_3/n7 , \pool/pool/pe_b/peij_0_3/n6 ,
         \pool/pool/pe_b/peij_0_3/n5 , \pool/pool/pe_b/peij_0_3/n4 ,
         \pool/pool/pe_b/peij_0_3/n3 , \pool/pool/pe_b/peij_0_3/n2 ,
         \pool/pool/pe_b/peij_0_3/n1 , \pool/pool/pe_b/peij_0_3/N36 ,
         \pool/pool/pe_b/peij_0_3/N35 , \pool/pool/pe_b/peij_0_3/N34 ,
         \pool/pool/pe_b/peij_0_3/N33 , \pool/pool/pe_b/peij_0_3/q_k ,
         \pool/pool/pe_b/peij_0_3/sgnext_10 ,
         \pool/pool/pe_b/peij_0_3/add/c_out ,
         \pool/pool/pe_b/peij_0_3/add/fai_0/n3 ,
         \pool/pool/pe_b/peij_0_3/add/fai_0/n1 ,
         \pool/pool/pe_b/peij_0_3/add/fai_1/n3 ,
         \pool/pool/pe_b/peij_0_3/add/fai_1/n1 ,
         \pool/pool/pe_b/peij_0_3/add/fai_2/n3 ,
         \pool/pool/pe_b/peij_0_3/add/fai_2/n1 ,
         \pool/pool/pe_b/peij_0_3/add/fai_3/n3 ,
         \pool/pool/pe_b/peij_0_3/add/fai_3/n1 ,
         \pool/pool/pe_b/peij_0_3/add/fai_4/n3 ,
         \pool/pool/pe_b/peij_0_3/add/fai_4/n1 ,
         \pool/pool/pe_b/peij_0_3/add/fai_5/n3 ,
         \pool/pool/pe_b/peij_0_3/add/fai_5/n1 ,
         \pool/pool/pe_b/peij_0_3/add/fai_6/n3 ,
         \pool/pool/pe_b/peij_0_3/add/fai_6/n1 ,
         \pool/pool/pe_b/peij_0_3/add/fai_7/n3 ,
         \pool/pool/pe_b/peij_0_3/add/fai_7/n1 ,
         \pool/pool/pe_b/peij_0_3/add/fai_8/n3 ,
         \pool/pool/pe_b/peij_0_3/add/fai_8/n1 ,
         \pool/pool/pe_b/peij_0_3/add/fai_9/n3 ,
         \pool/pool/pe_b/peij_0_3/add/fai_9/n1 ,
         \pool/pool/pe_b/peij_0_3/add/fai_10/n3 ,
         \pool/pool/pe_b/peij_0_3/add/fai_10/n1 ,
         \pool/pool/pe_b/peij_1_0/n18 , \pool/pool/pe_b/peij_1_0/n17 ,
         \pool/pool/pe_b/peij_1_0/n16 , \pool/pool/pe_b/peij_1_0/n12 ,
         \pool/pool/pe_b/peij_1_0/n11 , \pool/pool/pe_b/peij_1_0/n10 ,
         \pool/pool/pe_b/peij_1_0/n9 , \pool/pool/pe_b/peij_1_0/n8 ,
         \pool/pool/pe_b/peij_1_0/n7 , \pool/pool/pe_b/peij_1_0/n6 ,
         \pool/pool/pe_b/peij_1_0/n5 , \pool/pool/pe_b/peij_1_0/n4 ,
         \pool/pool/pe_b/peij_1_0/n3 , \pool/pool/pe_b/peij_1_0/n2 ,
         \pool/pool/pe_b/peij_1_0/n1 , \pool/pool/pe_b/peij_1_0/N36 ,
         \pool/pool/pe_b/peij_1_0/N35 , \pool/pool/pe_b/peij_1_0/N34 ,
         \pool/pool/pe_b/peij_1_0/N33 , \pool/pool/pe_b/peij_1_0/q_k ,
         \pool/pool/pe_b/peij_1_0/sgnext_10 ,
         \pool/pool/pe_b/peij_1_0/add/c_out ,
         \pool/pool/pe_b/peij_1_0/add/fai_0/n3 ,
         \pool/pool/pe_b/peij_1_0/add/fai_0/n1 ,
         \pool/pool/pe_b/peij_1_0/add/fai_1/n3 ,
         \pool/pool/pe_b/peij_1_0/add/fai_1/n1 ,
         \pool/pool/pe_b/peij_1_0/add/fai_2/n3 ,
         \pool/pool/pe_b/peij_1_0/add/fai_2/n1 ,
         \pool/pool/pe_b/peij_1_0/add/fai_3/n3 ,
         \pool/pool/pe_b/peij_1_0/add/fai_3/n1 ,
         \pool/pool/pe_b/peij_1_0/add/fai_4/n3 ,
         \pool/pool/pe_b/peij_1_0/add/fai_4/n1 ,
         \pool/pool/pe_b/peij_1_0/add/fai_5/n3 ,
         \pool/pool/pe_b/peij_1_0/add/fai_5/n1 ,
         \pool/pool/pe_b/peij_1_0/add/fai_6/n3 ,
         \pool/pool/pe_b/peij_1_0/add/fai_6/n1 ,
         \pool/pool/pe_b/peij_1_0/add/fai_7/n3 ,
         \pool/pool/pe_b/peij_1_0/add/fai_7/n1 ,
         \pool/pool/pe_b/peij_1_0/add/fai_8/n3 ,
         \pool/pool/pe_b/peij_1_0/add/fai_8/n1 ,
         \pool/pool/pe_b/peij_1_0/add/fai_9/n3 ,
         \pool/pool/pe_b/peij_1_0/add/fai_9/n1 ,
         \pool/pool/pe_b/peij_1_0/add/fai_10/n3 ,
         \pool/pool/pe_b/peij_1_0/add/fai_10/n1 ,
         \pool/pool/pe_b/peij_1_1/n18 , \pool/pool/pe_b/peij_1_1/n17 ,
         \pool/pool/pe_b/peij_1_1/n16 , \pool/pool/pe_b/peij_1_1/n12 ,
         \pool/pool/pe_b/peij_1_1/n11 , \pool/pool/pe_b/peij_1_1/n10 ,
         \pool/pool/pe_b/peij_1_1/n9 , \pool/pool/pe_b/peij_1_1/n8 ,
         \pool/pool/pe_b/peij_1_1/n7 , \pool/pool/pe_b/peij_1_1/n6 ,
         \pool/pool/pe_b/peij_1_1/n5 , \pool/pool/pe_b/peij_1_1/n4 ,
         \pool/pool/pe_b/peij_1_1/n3 , \pool/pool/pe_b/peij_1_1/n2 ,
         \pool/pool/pe_b/peij_1_1/n1 , \pool/pool/pe_b/peij_1_1/N36 ,
         \pool/pool/pe_b/peij_1_1/N35 , \pool/pool/pe_b/peij_1_1/N34 ,
         \pool/pool/pe_b/peij_1_1/N33 , \pool/pool/pe_b/peij_1_1/q_k ,
         \pool/pool/pe_b/peij_1_1/sgnext_10 ,
         \pool/pool/pe_b/peij_1_1/add/c_out ,
         \pool/pool/pe_b/peij_1_1/add/fai_0/n3 ,
         \pool/pool/pe_b/peij_1_1/add/fai_0/n1 ,
         \pool/pool/pe_b/peij_1_1/add/fai_1/n3 ,
         \pool/pool/pe_b/peij_1_1/add/fai_1/n1 ,
         \pool/pool/pe_b/peij_1_1/add/fai_2/n3 ,
         \pool/pool/pe_b/peij_1_1/add/fai_2/n1 ,
         \pool/pool/pe_b/peij_1_1/add/fai_3/n3 ,
         \pool/pool/pe_b/peij_1_1/add/fai_3/n1 ,
         \pool/pool/pe_b/peij_1_1/add/fai_4/n3 ,
         \pool/pool/pe_b/peij_1_1/add/fai_4/n1 ,
         \pool/pool/pe_b/peij_1_1/add/fai_5/n3 ,
         \pool/pool/pe_b/peij_1_1/add/fai_5/n1 ,
         \pool/pool/pe_b/peij_1_1/add/fai_6/n3 ,
         \pool/pool/pe_b/peij_1_1/add/fai_6/n1 ,
         \pool/pool/pe_b/peij_1_1/add/fai_7/n3 ,
         \pool/pool/pe_b/peij_1_1/add/fai_7/n1 ,
         \pool/pool/pe_b/peij_1_1/add/fai_8/n3 ,
         \pool/pool/pe_b/peij_1_1/add/fai_8/n1 ,
         \pool/pool/pe_b/peij_1_1/add/fai_9/n3 ,
         \pool/pool/pe_b/peij_1_1/add/fai_9/n1 ,
         \pool/pool/pe_b/peij_1_1/add/fai_10/n3 ,
         \pool/pool/pe_b/peij_1_1/add/fai_10/n1 ,
         \pool/pool/pe_b/peij_1_2/n18 , \pool/pool/pe_b/peij_1_2/n17 ,
         \pool/pool/pe_b/peij_1_2/n16 , \pool/pool/pe_b/peij_1_2/n12 ,
         \pool/pool/pe_b/peij_1_2/n11 , \pool/pool/pe_b/peij_1_2/n10 ,
         \pool/pool/pe_b/peij_1_2/n9 , \pool/pool/pe_b/peij_1_2/n8 ,
         \pool/pool/pe_b/peij_1_2/n7 , \pool/pool/pe_b/peij_1_2/n6 ,
         \pool/pool/pe_b/peij_1_2/n5 , \pool/pool/pe_b/peij_1_2/n4 ,
         \pool/pool/pe_b/peij_1_2/n3 , \pool/pool/pe_b/peij_1_2/n2 ,
         \pool/pool/pe_b/peij_1_2/n1 , \pool/pool/pe_b/peij_1_2/N36 ,
         \pool/pool/pe_b/peij_1_2/N35 , \pool/pool/pe_b/peij_1_2/N34 ,
         \pool/pool/pe_b/peij_1_2/N33 , \pool/pool/pe_b/peij_1_2/q_k ,
         \pool/pool/pe_b/peij_1_2/sgnext_10 ,
         \pool/pool/pe_b/peij_1_2/add/c_out ,
         \pool/pool/pe_b/peij_1_2/add/fai_0/n3 ,
         \pool/pool/pe_b/peij_1_2/add/fai_0/n1 ,
         \pool/pool/pe_b/peij_1_2/add/fai_1/n3 ,
         \pool/pool/pe_b/peij_1_2/add/fai_1/n1 ,
         \pool/pool/pe_b/peij_1_2/add/fai_2/n3 ,
         \pool/pool/pe_b/peij_1_2/add/fai_2/n1 ,
         \pool/pool/pe_b/peij_1_2/add/fai_3/n3 ,
         \pool/pool/pe_b/peij_1_2/add/fai_3/n1 ,
         \pool/pool/pe_b/peij_1_2/add/fai_4/n3 ,
         \pool/pool/pe_b/peij_1_2/add/fai_4/n1 ,
         \pool/pool/pe_b/peij_1_2/add/fai_5/n3 ,
         \pool/pool/pe_b/peij_1_2/add/fai_5/n1 ,
         \pool/pool/pe_b/peij_1_2/add/fai_6/n3 ,
         \pool/pool/pe_b/peij_1_2/add/fai_6/n1 ,
         \pool/pool/pe_b/peij_1_2/add/fai_7/n3 ,
         \pool/pool/pe_b/peij_1_2/add/fai_7/n1 ,
         \pool/pool/pe_b/peij_1_2/add/fai_8/n3 ,
         \pool/pool/pe_b/peij_1_2/add/fai_8/n1 ,
         \pool/pool/pe_b/peij_1_2/add/fai_9/n3 ,
         \pool/pool/pe_b/peij_1_2/add/fai_9/n1 ,
         \pool/pool/pe_b/peij_1_2/add/fai_10/n3 ,
         \pool/pool/pe_b/peij_1_2/add/fai_10/n1 ,
         \pool/pool/pe_b/peij_1_3/n18 , \pool/pool/pe_b/peij_1_3/n17 ,
         \pool/pool/pe_b/peij_1_3/n16 , \pool/pool/pe_b/peij_1_3/n12 ,
         \pool/pool/pe_b/peij_1_3/n11 , \pool/pool/pe_b/peij_1_3/n10 ,
         \pool/pool/pe_b/peij_1_3/n9 , \pool/pool/pe_b/peij_1_3/n8 ,
         \pool/pool/pe_b/peij_1_3/n7 , \pool/pool/pe_b/peij_1_3/n6 ,
         \pool/pool/pe_b/peij_1_3/n5 , \pool/pool/pe_b/peij_1_3/n4 ,
         \pool/pool/pe_b/peij_1_3/n3 , \pool/pool/pe_b/peij_1_3/n2 ,
         \pool/pool/pe_b/peij_1_3/n1 , \pool/pool/pe_b/peij_1_3/N36 ,
         \pool/pool/pe_b/peij_1_3/N35 , \pool/pool/pe_b/peij_1_3/N34 ,
         \pool/pool/pe_b/peij_1_3/N33 , \pool/pool/pe_b/peij_1_3/q_k ,
         \pool/pool/pe_b/peij_1_3/sgnext_10 ,
         \pool/pool/pe_b/peij_1_3/add/c_out ,
         \pool/pool/pe_b/peij_1_3/add/fai_0/n3 ,
         \pool/pool/pe_b/peij_1_3/add/fai_0/n1 ,
         \pool/pool/pe_b/peij_1_3/add/fai_1/n3 ,
         \pool/pool/pe_b/peij_1_3/add/fai_1/n1 ,
         \pool/pool/pe_b/peij_1_3/add/fai_2/n3 ,
         \pool/pool/pe_b/peij_1_3/add/fai_2/n1 ,
         \pool/pool/pe_b/peij_1_3/add/fai_3/n3 ,
         \pool/pool/pe_b/peij_1_3/add/fai_3/n1 ,
         \pool/pool/pe_b/peij_1_3/add/fai_4/n3 ,
         \pool/pool/pe_b/peij_1_3/add/fai_4/n1 ,
         \pool/pool/pe_b/peij_1_3/add/fai_5/n3 ,
         \pool/pool/pe_b/peij_1_3/add/fai_5/n1 ,
         \pool/pool/pe_b/peij_1_3/add/fai_6/n3 ,
         \pool/pool/pe_b/peij_1_3/add/fai_6/n1 ,
         \pool/pool/pe_b/peij_1_3/add/fai_7/n3 ,
         \pool/pool/pe_b/peij_1_3/add/fai_7/n1 ,
         \pool/pool/pe_b/peij_1_3/add/fai_8/n3 ,
         \pool/pool/pe_b/peij_1_3/add/fai_8/n1 ,
         \pool/pool/pe_b/peij_1_3/add/fai_9/n3 ,
         \pool/pool/pe_b/peij_1_3/add/fai_9/n1 ,
         \pool/pool/pe_b/peij_1_3/add/fai_10/n3 ,
         \pool/pool/pe_b/peij_1_3/add/fai_10/n1 ,
         \pool/pool/pe_b/peij_2_0/n18 , \pool/pool/pe_b/peij_2_0/n17 ,
         \pool/pool/pe_b/peij_2_0/n16 , \pool/pool/pe_b/peij_2_0/n12 ,
         \pool/pool/pe_b/peij_2_0/n11 , \pool/pool/pe_b/peij_2_0/n10 ,
         \pool/pool/pe_b/peij_2_0/n9 , \pool/pool/pe_b/peij_2_0/n8 ,
         \pool/pool/pe_b/peij_2_0/n7 , \pool/pool/pe_b/peij_2_0/n6 ,
         \pool/pool/pe_b/peij_2_0/n5 , \pool/pool/pe_b/peij_2_0/n4 ,
         \pool/pool/pe_b/peij_2_0/n3 , \pool/pool/pe_b/peij_2_0/n2 ,
         \pool/pool/pe_b/peij_2_0/n1 , \pool/pool/pe_b/peij_2_0/N36 ,
         \pool/pool/pe_b/peij_2_0/N35 , \pool/pool/pe_b/peij_2_0/N34 ,
         \pool/pool/pe_b/peij_2_0/N33 , \pool/pool/pe_b/peij_2_0/q_k ,
         \pool/pool/pe_b/peij_2_0/sgnext_10 ,
         \pool/pool/pe_b/peij_2_0/add/c_out ,
         \pool/pool/pe_b/peij_2_0/add/fai_0/n3 ,
         \pool/pool/pe_b/peij_2_0/add/fai_0/n1 ,
         \pool/pool/pe_b/peij_2_0/add/fai_1/n3 ,
         \pool/pool/pe_b/peij_2_0/add/fai_1/n1 ,
         \pool/pool/pe_b/peij_2_0/add/fai_2/n3 ,
         \pool/pool/pe_b/peij_2_0/add/fai_2/n1 ,
         \pool/pool/pe_b/peij_2_0/add/fai_3/n3 ,
         \pool/pool/pe_b/peij_2_0/add/fai_3/n1 ,
         \pool/pool/pe_b/peij_2_0/add/fai_4/n3 ,
         \pool/pool/pe_b/peij_2_0/add/fai_4/n1 ,
         \pool/pool/pe_b/peij_2_0/add/fai_5/n3 ,
         \pool/pool/pe_b/peij_2_0/add/fai_5/n1 ,
         \pool/pool/pe_b/peij_2_0/add/fai_6/n3 ,
         \pool/pool/pe_b/peij_2_0/add/fai_6/n1 ,
         \pool/pool/pe_b/peij_2_0/add/fai_7/n3 ,
         \pool/pool/pe_b/peij_2_0/add/fai_7/n1 ,
         \pool/pool/pe_b/peij_2_0/add/fai_8/n3 ,
         \pool/pool/pe_b/peij_2_0/add/fai_8/n1 ,
         \pool/pool/pe_b/peij_2_0/add/fai_9/n3 ,
         \pool/pool/pe_b/peij_2_0/add/fai_9/n1 ,
         \pool/pool/pe_b/peij_2_0/add/fai_10/n3 ,
         \pool/pool/pe_b/peij_2_0/add/fai_10/n1 ,
         \pool/pool/pe_b/peij_2_1/n18 , \pool/pool/pe_b/peij_2_1/n17 ,
         \pool/pool/pe_b/peij_2_1/n16 , \pool/pool/pe_b/peij_2_1/n12 ,
         \pool/pool/pe_b/peij_2_1/n11 , \pool/pool/pe_b/peij_2_1/n10 ,
         \pool/pool/pe_b/peij_2_1/n9 , \pool/pool/pe_b/peij_2_1/n8 ,
         \pool/pool/pe_b/peij_2_1/n7 , \pool/pool/pe_b/peij_2_1/n6 ,
         \pool/pool/pe_b/peij_2_1/n5 , \pool/pool/pe_b/peij_2_1/n4 ,
         \pool/pool/pe_b/peij_2_1/n3 , \pool/pool/pe_b/peij_2_1/n2 ,
         \pool/pool/pe_b/peij_2_1/n1 , \pool/pool/pe_b/peij_2_1/N36 ,
         \pool/pool/pe_b/peij_2_1/N35 , \pool/pool/pe_b/peij_2_1/N34 ,
         \pool/pool/pe_b/peij_2_1/N33 , \pool/pool/pe_b/peij_2_1/q_k ,
         \pool/pool/pe_b/peij_2_1/sgnext_10 ,
         \pool/pool/pe_b/peij_2_1/add/c_out ,
         \pool/pool/pe_b/peij_2_1/add/fai_0/n3 ,
         \pool/pool/pe_b/peij_2_1/add/fai_0/n1 ,
         \pool/pool/pe_b/peij_2_1/add/fai_1/n3 ,
         \pool/pool/pe_b/peij_2_1/add/fai_1/n1 ,
         \pool/pool/pe_b/peij_2_1/add/fai_2/n3 ,
         \pool/pool/pe_b/peij_2_1/add/fai_2/n1 ,
         \pool/pool/pe_b/peij_2_1/add/fai_3/n3 ,
         \pool/pool/pe_b/peij_2_1/add/fai_3/n1 ,
         \pool/pool/pe_b/peij_2_1/add/fai_4/n3 ,
         \pool/pool/pe_b/peij_2_1/add/fai_4/n1 ,
         \pool/pool/pe_b/peij_2_1/add/fai_5/n3 ,
         \pool/pool/pe_b/peij_2_1/add/fai_5/n1 ,
         \pool/pool/pe_b/peij_2_1/add/fai_6/n3 ,
         \pool/pool/pe_b/peij_2_1/add/fai_6/n1 ,
         \pool/pool/pe_b/peij_2_1/add/fai_7/n3 ,
         \pool/pool/pe_b/peij_2_1/add/fai_7/n1 ,
         \pool/pool/pe_b/peij_2_1/add/fai_8/n3 ,
         \pool/pool/pe_b/peij_2_1/add/fai_8/n1 ,
         \pool/pool/pe_b/peij_2_1/add/fai_9/n3 ,
         \pool/pool/pe_b/peij_2_1/add/fai_9/n1 ,
         \pool/pool/pe_b/peij_2_1/add/fai_10/n3 ,
         \pool/pool/pe_b/peij_2_1/add/fai_10/n1 ,
         \pool/pool/pe_b/peij_2_2/n18 , \pool/pool/pe_b/peij_2_2/n17 ,
         \pool/pool/pe_b/peij_2_2/n16 , \pool/pool/pe_b/peij_2_2/n12 ,
         \pool/pool/pe_b/peij_2_2/n11 , \pool/pool/pe_b/peij_2_2/n10 ,
         \pool/pool/pe_b/peij_2_2/n9 , \pool/pool/pe_b/peij_2_2/n8 ,
         \pool/pool/pe_b/peij_2_2/n7 , \pool/pool/pe_b/peij_2_2/n6 ,
         \pool/pool/pe_b/peij_2_2/n5 , \pool/pool/pe_b/peij_2_2/n4 ,
         \pool/pool/pe_b/peij_2_2/n3 , \pool/pool/pe_b/peij_2_2/n2 ,
         \pool/pool/pe_b/peij_2_2/n1 , \pool/pool/pe_b/peij_2_2/N36 ,
         \pool/pool/pe_b/peij_2_2/N35 , \pool/pool/pe_b/peij_2_2/N34 ,
         \pool/pool/pe_b/peij_2_2/N33 , \pool/pool/pe_b/peij_2_2/q_k ,
         \pool/pool/pe_b/peij_2_2/sgnext_10 ,
         \pool/pool/pe_b/peij_2_2/add/c_out ,
         \pool/pool/pe_b/peij_2_2/add/fai_0/n3 ,
         \pool/pool/pe_b/peij_2_2/add/fai_0/n1 ,
         \pool/pool/pe_b/peij_2_2/add/fai_1/n3 ,
         \pool/pool/pe_b/peij_2_2/add/fai_1/n1 ,
         \pool/pool/pe_b/peij_2_2/add/fai_2/n3 ,
         \pool/pool/pe_b/peij_2_2/add/fai_2/n1 ,
         \pool/pool/pe_b/peij_2_2/add/fai_3/n3 ,
         \pool/pool/pe_b/peij_2_2/add/fai_3/n1 ,
         \pool/pool/pe_b/peij_2_2/add/fai_4/n3 ,
         \pool/pool/pe_b/peij_2_2/add/fai_4/n1 ,
         \pool/pool/pe_b/peij_2_2/add/fai_5/n3 ,
         \pool/pool/pe_b/peij_2_2/add/fai_5/n1 ,
         \pool/pool/pe_b/peij_2_2/add/fai_6/n3 ,
         \pool/pool/pe_b/peij_2_2/add/fai_6/n1 ,
         \pool/pool/pe_b/peij_2_2/add/fai_7/n3 ,
         \pool/pool/pe_b/peij_2_2/add/fai_7/n1 ,
         \pool/pool/pe_b/peij_2_2/add/fai_8/n3 ,
         \pool/pool/pe_b/peij_2_2/add/fai_8/n1 ,
         \pool/pool/pe_b/peij_2_2/add/fai_9/n3 ,
         \pool/pool/pe_b/peij_2_2/add/fai_9/n1 ,
         \pool/pool/pe_b/peij_2_2/add/fai_10/n3 ,
         \pool/pool/pe_b/peij_2_2/add/fai_10/n1 ,
         \pool/pool/pe_b/peij_2_3/n18 , \pool/pool/pe_b/peij_2_3/n17 ,
         \pool/pool/pe_b/peij_2_3/n16 , \pool/pool/pe_b/peij_2_3/n12 ,
         \pool/pool/pe_b/peij_2_3/n11 , \pool/pool/pe_b/peij_2_3/n10 ,
         \pool/pool/pe_b/peij_2_3/n9 , \pool/pool/pe_b/peij_2_3/n8 ,
         \pool/pool/pe_b/peij_2_3/n7 , \pool/pool/pe_b/peij_2_3/n6 ,
         \pool/pool/pe_b/peij_2_3/n5 , \pool/pool/pe_b/peij_2_3/n4 ,
         \pool/pool/pe_b/peij_2_3/n3 , \pool/pool/pe_b/peij_2_3/n2 ,
         \pool/pool/pe_b/peij_2_3/n1 , \pool/pool/pe_b/peij_2_3/N36 ,
         \pool/pool/pe_b/peij_2_3/N35 , \pool/pool/pe_b/peij_2_3/N34 ,
         \pool/pool/pe_b/peij_2_3/N33 , \pool/pool/pe_b/peij_2_3/q_k ,
         \pool/pool/pe_b/peij_2_3/sgnext_10 ,
         \pool/pool/pe_b/peij_2_3/add/c_out ,
         \pool/pool/pe_b/peij_2_3/add/fai_0/n3 ,
         \pool/pool/pe_b/peij_2_3/add/fai_0/n1 ,
         \pool/pool/pe_b/peij_2_3/add/fai_1/n3 ,
         \pool/pool/pe_b/peij_2_3/add/fai_1/n1 ,
         \pool/pool/pe_b/peij_2_3/add/fai_2/n3 ,
         \pool/pool/pe_b/peij_2_3/add/fai_2/n1 ,
         \pool/pool/pe_b/peij_2_3/add/fai_3/n3 ,
         \pool/pool/pe_b/peij_2_3/add/fai_3/n1 ,
         \pool/pool/pe_b/peij_2_3/add/fai_4/n3 ,
         \pool/pool/pe_b/peij_2_3/add/fai_4/n1 ,
         \pool/pool/pe_b/peij_2_3/add/fai_5/n3 ,
         \pool/pool/pe_b/peij_2_3/add/fai_5/n1 ,
         \pool/pool/pe_b/peij_2_3/add/fai_6/n3 ,
         \pool/pool/pe_b/peij_2_3/add/fai_6/n1 ,
         \pool/pool/pe_b/peij_2_3/add/fai_7/n3 ,
         \pool/pool/pe_b/peij_2_3/add/fai_7/n1 ,
         \pool/pool/pe_b/peij_2_3/add/fai_8/n3 ,
         \pool/pool/pe_b/peij_2_3/add/fai_8/n1 ,
         \pool/pool/pe_b/peij_2_3/add/fai_9/n3 ,
         \pool/pool/pe_b/peij_2_3/add/fai_9/n1 ,
         \pool/pool/pe_b/peij_2_3/add/fai_10/n3 ,
         \pool/pool/pe_b/peij_2_3/add/fai_10/n1 ,
         \pool/pool/pe_b/peij_3_0/n18 , \pool/pool/pe_b/peij_3_0/n17 ,
         \pool/pool/pe_b/peij_3_0/n16 , \pool/pool/pe_b/peij_3_0/n12 ,
         \pool/pool/pe_b/peij_3_0/n11 , \pool/pool/pe_b/peij_3_0/n10 ,
         \pool/pool/pe_b/peij_3_0/n9 , \pool/pool/pe_b/peij_3_0/n8 ,
         \pool/pool/pe_b/peij_3_0/n7 , \pool/pool/pe_b/peij_3_0/n6 ,
         \pool/pool/pe_b/peij_3_0/n5 , \pool/pool/pe_b/peij_3_0/n4 ,
         \pool/pool/pe_b/peij_3_0/n3 , \pool/pool/pe_b/peij_3_0/n2 ,
         \pool/pool/pe_b/peij_3_0/n1 , \pool/pool/pe_b/peij_3_0/N36 ,
         \pool/pool/pe_b/peij_3_0/N35 , \pool/pool/pe_b/peij_3_0/N34 ,
         \pool/pool/pe_b/peij_3_0/N33 , \pool/pool/pe_b/peij_3_0/q_k ,
         \pool/pool/pe_b/peij_3_0/sgnext_10 ,
         \pool/pool/pe_b/peij_3_0/add/c_out ,
         \pool/pool/pe_b/peij_3_0/add/fai_0/n3 ,
         \pool/pool/pe_b/peij_3_0/add/fai_0/n1 ,
         \pool/pool/pe_b/peij_3_0/add/fai_1/n3 ,
         \pool/pool/pe_b/peij_3_0/add/fai_1/n1 ,
         \pool/pool/pe_b/peij_3_0/add/fai_2/n3 ,
         \pool/pool/pe_b/peij_3_0/add/fai_2/n1 ,
         \pool/pool/pe_b/peij_3_0/add/fai_3/n3 ,
         \pool/pool/pe_b/peij_3_0/add/fai_3/n1 ,
         \pool/pool/pe_b/peij_3_0/add/fai_4/n3 ,
         \pool/pool/pe_b/peij_3_0/add/fai_4/n1 ,
         \pool/pool/pe_b/peij_3_0/add/fai_5/n3 ,
         \pool/pool/pe_b/peij_3_0/add/fai_5/n1 ,
         \pool/pool/pe_b/peij_3_0/add/fai_6/n3 ,
         \pool/pool/pe_b/peij_3_0/add/fai_6/n1 ,
         \pool/pool/pe_b/peij_3_0/add/fai_7/n3 ,
         \pool/pool/pe_b/peij_3_0/add/fai_7/n1 ,
         \pool/pool/pe_b/peij_3_0/add/fai_8/n3 ,
         \pool/pool/pe_b/peij_3_0/add/fai_8/n1 ,
         \pool/pool/pe_b/peij_3_0/add/fai_9/n3 ,
         \pool/pool/pe_b/peij_3_0/add/fai_9/n1 ,
         \pool/pool/pe_b/peij_3_0/add/fai_10/n3 ,
         \pool/pool/pe_b/peij_3_0/add/fai_10/n1 ,
         \pool/pool/pe_b/peij_3_1/n18 , \pool/pool/pe_b/peij_3_1/n17 ,
         \pool/pool/pe_b/peij_3_1/n16 , \pool/pool/pe_b/peij_3_1/n12 ,
         \pool/pool/pe_b/peij_3_1/n11 , \pool/pool/pe_b/peij_3_1/n10 ,
         \pool/pool/pe_b/peij_3_1/n9 , \pool/pool/pe_b/peij_3_1/n8 ,
         \pool/pool/pe_b/peij_3_1/n7 , \pool/pool/pe_b/peij_3_1/n6 ,
         \pool/pool/pe_b/peij_3_1/n5 , \pool/pool/pe_b/peij_3_1/n4 ,
         \pool/pool/pe_b/peij_3_1/n3 , \pool/pool/pe_b/peij_3_1/n2 ,
         \pool/pool/pe_b/peij_3_1/n1 , \pool/pool/pe_b/peij_3_1/N36 ,
         \pool/pool/pe_b/peij_3_1/N35 , \pool/pool/pe_b/peij_3_1/N34 ,
         \pool/pool/pe_b/peij_3_1/N33 , \pool/pool/pe_b/peij_3_1/q_k ,
         \pool/pool/pe_b/peij_3_1/sgnext_10 ,
         \pool/pool/pe_b/peij_3_1/add/c_out ,
         \pool/pool/pe_b/peij_3_1/add/fai_0/n3 ,
         \pool/pool/pe_b/peij_3_1/add/fai_0/n1 ,
         \pool/pool/pe_b/peij_3_1/add/fai_1/n3 ,
         \pool/pool/pe_b/peij_3_1/add/fai_1/n1 ,
         \pool/pool/pe_b/peij_3_1/add/fai_2/n3 ,
         \pool/pool/pe_b/peij_3_1/add/fai_2/n1 ,
         \pool/pool/pe_b/peij_3_1/add/fai_3/n3 ,
         \pool/pool/pe_b/peij_3_1/add/fai_3/n1 ,
         \pool/pool/pe_b/peij_3_1/add/fai_4/n3 ,
         \pool/pool/pe_b/peij_3_1/add/fai_4/n1 ,
         \pool/pool/pe_b/peij_3_1/add/fai_5/n3 ,
         \pool/pool/pe_b/peij_3_1/add/fai_5/n1 ,
         \pool/pool/pe_b/peij_3_1/add/fai_6/n3 ,
         \pool/pool/pe_b/peij_3_1/add/fai_6/n1 ,
         \pool/pool/pe_b/peij_3_1/add/fai_7/n3 ,
         \pool/pool/pe_b/peij_3_1/add/fai_7/n1 ,
         \pool/pool/pe_b/peij_3_1/add/fai_8/n3 ,
         \pool/pool/pe_b/peij_3_1/add/fai_8/n1 ,
         \pool/pool/pe_b/peij_3_1/add/fai_9/n3 ,
         \pool/pool/pe_b/peij_3_1/add/fai_9/n1 ,
         \pool/pool/pe_b/peij_3_1/add/fai_10/n3 ,
         \pool/pool/pe_b/peij_3_1/add/fai_10/n1 ,
         \pool/pool/pe_b/peij_3_2/n19 , \pool/pool/pe_b/peij_3_2/n18 ,
         \pool/pool/pe_b/peij_3_2/n17 , \pool/pool/pe_b/peij_3_2/n16 ,
         \pool/pool/pe_b/peij_3_2/n12 , \pool/pool/pe_b/peij_3_2/n11 ,
         \pool/pool/pe_b/peij_3_2/n10 , \pool/pool/pe_b/peij_3_2/n9 ,
         \pool/pool/pe_b/peij_3_2/n8 , \pool/pool/pe_b/peij_3_2/n7 ,
         \pool/pool/pe_b/peij_3_2/n6 , \pool/pool/pe_b/peij_3_2/n5 ,
         \pool/pool/pe_b/peij_3_2/n4 , \pool/pool/pe_b/peij_3_2/n3 ,
         \pool/pool/pe_b/peij_3_2/n2 , \pool/pool/pe_b/peij_3_2/N36 ,
         \pool/pool/pe_b/peij_3_2/N34 , \pool/pool/pe_b/peij_3_2/N33 ,
         \pool/pool/pe_b/peij_3_2/q_k , \pool/pool/pe_b/peij_3_2/sgnext_10 ,
         \pool/pool/pe_b/peij_3_2/add/c_out ,
         \pool/pool/pe_b/peij_3_2/add/fai_0/n3 ,
         \pool/pool/pe_b/peij_3_2/add/fai_0/n1 ,
         \pool/pool/pe_b/peij_3_2/add/fai_1/n3 ,
         \pool/pool/pe_b/peij_3_2/add/fai_1/n1 ,
         \pool/pool/pe_b/peij_3_2/add/fai_2/n3 ,
         \pool/pool/pe_b/peij_3_2/add/fai_2/n1 ,
         \pool/pool/pe_b/peij_3_2/add/fai_3/n3 ,
         \pool/pool/pe_b/peij_3_2/add/fai_3/n1 ,
         \pool/pool/pe_b/peij_3_2/add/fai_4/n3 ,
         \pool/pool/pe_b/peij_3_2/add/fai_4/n1 ,
         \pool/pool/pe_b/peij_3_2/add/fai_5/n3 ,
         \pool/pool/pe_b/peij_3_2/add/fai_5/n1 ,
         \pool/pool/pe_b/peij_3_2/add/fai_6/n3 ,
         \pool/pool/pe_b/peij_3_2/add/fai_6/n1 ,
         \pool/pool/pe_b/peij_3_2/add/fai_7/n3 ,
         \pool/pool/pe_b/peij_3_2/add/fai_7/n1 ,
         \pool/pool/pe_b/peij_3_2/add/fai_8/n3 ,
         \pool/pool/pe_b/peij_3_2/add/fai_8/n1 ,
         \pool/pool/pe_b/peij_3_2/add/fai_9/n3 ,
         \pool/pool/pe_b/peij_3_2/add/fai_9/n1 ,
         \pool/pool/pe_b/peij_3_2/add/fai_10/n3 ,
         \pool/pool/pe_b/peij_3_2/add/fai_10/n1 ,
         \pool/pool/pe_b/peij_3_3/n18 , \pool/pool/pe_b/peij_3_3/n17 ,
         \pool/pool/pe_b/peij_3_3/n16 , \pool/pool/pe_b/peij_3_3/n12 ,
         \pool/pool/pe_b/peij_3_3/n11 , \pool/pool/pe_b/peij_3_3/n10 ,
         \pool/pool/pe_b/peij_3_3/n9 , \pool/pool/pe_b/peij_3_3/n8 ,
         \pool/pool/pe_b/peij_3_3/n7 , \pool/pool/pe_b/peij_3_3/n6 ,
         \pool/pool/pe_b/peij_3_3/n5 , \pool/pool/pe_b/peij_3_3/n4 ,
         \pool/pool/pe_b/peij_3_3/n3 , \pool/pool/pe_b/peij_3_3/n2 ,
         \pool/pool/pe_b/peij_3_3/n1 , \pool/pool/pe_b/peij_3_3/N36 ,
         \pool/pool/pe_b/peij_3_3/N35 , \pool/pool/pe_b/peij_3_3/N34 ,
         \pool/pool/pe_b/peij_3_3/N33 , \pool/pool/pe_b/peij_3_3/q_k ,
         \pool/pool/pe_b/peij_3_3/sgnext_10 ,
         \pool/pool/pe_b/peij_3_3/add/c_out ,
         \pool/pool/pe_b/peij_3_3/add/fai_0/n3 ,
         \pool/pool/pe_b/peij_3_3/add/fai_0/n1 ,
         \pool/pool/pe_b/peij_3_3/add/fai_1/n3 ,
         \pool/pool/pe_b/peij_3_3/add/fai_1/n1 ,
         \pool/pool/pe_b/peij_3_3/add/fai_2/n3 ,
         \pool/pool/pe_b/peij_3_3/add/fai_2/n1 ,
         \pool/pool/pe_b/peij_3_3/add/fai_3/n3 ,
         \pool/pool/pe_b/peij_3_3/add/fai_3/n1 ,
         \pool/pool/pe_b/peij_3_3/add/fai_4/n3 ,
         \pool/pool/pe_b/peij_3_3/add/fai_4/n1 ,
         \pool/pool/pe_b/peij_3_3/add/fai_5/n3 ,
         \pool/pool/pe_b/peij_3_3/add/fai_5/n1 ,
         \pool/pool/pe_b/peij_3_3/add/fai_6/n3 ,
         \pool/pool/pe_b/peij_3_3/add/fai_6/n1 ,
         \pool/pool/pe_b/peij_3_3/add/fai_7/n3 ,
         \pool/pool/pe_b/peij_3_3/add/fai_7/n1 ,
         \pool/pool/pe_b/peij_3_3/add/fai_8/n3 ,
         \pool/pool/pe_b/peij_3_3/add/fai_8/n1 ,
         \pool/pool/pe_b/peij_3_3/add/fai_9/n3 ,
         \pool/pool/pe_b/peij_3_3/add/fai_9/n1 ,
         \pool/pool/pe_b/peij_3_3/add/fai_10/n3 ,
         \pool/pool/pe_b/peij_3_3/add/fai_10/n1 , \pool/pool/count/n18 ,
         \pool/pool/count/n17 , \pool/pool/count/n16 , \pool/pool/count/n15 ,
         \pool/pool/count/n14 , \pool/pool/count/n13 , \pool/pool/count/n12 ,
         \pool/pool/count/n11 , \pool/pool/count/n10 , \pool/pool/count/n9 ,
         \pool/pool/count/n8 , \pool/pool/count/n7 , \pool/pool/count/n6 ,
         \pool/pool/count/n5 , \pool/pool/count/n4 , \pool/pool/count/n3 ,
         \pool/pool/shift_row0/n12 , \pool/pool/shift_row0/n11 ,
         \pool/pool/shift_row0/n10 , \pool/pool/shift_row0/n9 ,
         \pool/pool/shift_row0/n8 , \pool/pool/shift_row0/n7 ,
         \pool/pool/shift_row0/n6 , \pool/pool/shift_row0/n5 ,
         \pool/pool/shift_row0/n4 , \pool/pool/shift_row0/n3 ,
         \pool/pool/shift_row0/n2 , \pool/pool/shift_row0/n1 ,
         \pool/pool/shift_row1/n24 , \pool/pool/shift_row1/n23 ,
         \pool/pool/shift_row1/n22 , \pool/pool/shift_row1/n21 ,
         \pool/pool/shift_row1/n20 , \pool/pool/shift_row1/n19 ,
         \pool/pool/shift_row1/n18 , \pool/pool/shift_row1/n17 ,
         \pool/pool/shift_row1/n16 , \pool/pool/shift_row1/n15 ,
         \pool/pool/shift_row1/n14 , \pool/pool/shift_row1/n13 ,
         \pool/pool/shift_row2/n24 , \pool/pool/shift_row2/n23 ,
         \pool/pool/shift_row2/n22 , \pool/pool/shift_row2/n21 ,
         \pool/pool/shift_row2/n20 , \pool/pool/shift_row2/n19 ,
         \pool/pool/shift_row2/n18 , \pool/pool/shift_row2/n17 ,
         \pool/pool/shift_row2/n16 , \pool/pool/shift_row2/n15 ,
         \pool/pool/shift_row2/n14 , \pool/pool/shift_row2/n13 ,
         \pool/pool/shift_row3/n24 , \pool/pool/shift_row3/n23 ,
         \pool/pool/shift_row3/n22 , \pool/pool/shift_row3/n21 ,
         \pool/pool/shift_row3/n20 , \pool/pool/shift_row3/n19 ,
         \pool/pool/shift_row3/n18 , \pool/pool/shift_row3/n17 ,
         \pool/pool/shift_row3/n16 , \pool/pool/shift_row3/n15 ,
         \pool/pool/shift_row3/n14 , \pool/pool/shift_row3/n13 ,
         \pool/fsm/n17 , \pool/fsm/n4 , \pool/fsm/n18 , \pool/fsm/n16 ,
         \pool/fsm/n15 , \pool/fsm/n14 , \pool/fsm/n13 , \pool/fsm/n12 ,
         \pool/fsm/n11 , \pool/fsm/n10 , \pool/fsm/n9 , \pool/fsm/n8 ,
         \pool/fsm/n6 , \pool/fsm/n5 , \pool/fsm/n3 , \pool/fsm/n1 ,
         \pool/fsm/net468 , \pool/fsm/N31 , \pool/fsm/N29 , \pool/fsm/N28 ,
         \pool/fsm/N11 , \pool/fsm/current_state[0] ,
         \pool/fsm/current_state[1] , \pool/fsm/current_state[2] ,
         \pool/gate_clk/n32 , \pool/gate_clk/n31 , \pool/gate_clk/n30 ,
         \pool/gate_clk/n14 , \pool/gate_clk/n13 , \pool/gate_clk/n2 ,
         \pool/gate_clk/n1 , \pool/gate_clk/n29 , \pool/gate_clk/n28 ,
         \pool/gate_clk/n27 , \pool/gate_clk/n26 , \pool/gate_clk/n25 ,
         \pool/gate_clk/n24 , \pool/gate_clk/n23 , \pool/gate_clk/n22 ,
         \pool/gate_clk/n21 , \pool/gate_clk/n20 , \pool/gate_clk/n19 ,
         \pool/gate_clk/n18 , \pool/gate_clk/n17 , \pool/gate_clk/n16 ,
         \pool/gate_clk/n15 , \pool/gate_clk/n12 , \pool/gate_clk/n11 ,
         \pool/gate_clk/n10 , \pool/gate_clk/n9 , \pool/gate_clk/n8 ,
         \pool/gate_clk/n7 , \pool/gate_clk/n6 , \pool/gate_clk/n5 ,
         \pool/gate_clk/n4 , \pool/gate_clk/n3 , \pool/gate_clk/del_tc_r_1 ,
         \pool/gate_clk/N45 , \pool/gate_clk/del_tc_r ,
         \pool/gate_clk/cnt_r_out[0] , \pool/gate_clk/cnt_r_out[1] ,
         \pool/gate_clk/tc_c , \pool/gate_clk/cnt_c_out[0] ,
         \pool/gate_clk/cnt_c_out[1] , \pool/gate_clk/del_1_tc ,
         \pool/gate_clk/N21 , \pool/gate_clk/del_0_tc ,
         \pool/gate_clk/dec_out[0] , \pool/gate_clk/dec_out[1] ,
         \pool/gate_clk/dec_out[2] , \pool/gate_clk/pool_size[0] ,
         \pool/gate_clk/pool_size[1] , \pool/gate_clk/pool_size[2] ,
         \pool/gate_clk/pool_size[3] , \pool/gate_clk/pool_size[4] ,
         \pool/gate_clk/mux_pool/n11 , \pool/gate_clk/mux_pool/n10 ,
         \pool/gate_clk/mux_pool/n9 , \pool/gate_clk/mux_pool/n8 ,
         \pool/gate_clk/mux_pool/n7 , \pool/gate_clk/mux_pool/n6 ,
         \pool/gate_clk/mux_cmask/n9 , \pool/gate_clk/mux_cmask/n8 ,
         \pool/gate_clk/mux_cmask/n7 , \pool/gate_clk/mux_cmask/n6 ,
         \pool/gate_clk/mux_cmask/n5 , \pool/gate_clk/mux_rmask/n6 ,
         \pool/gate_clk/mux_rmask/n4 , \pool/gate_clk/mux_rmask/n3 ,
         \pool/gate_clk/mux_rmask/n2 , \pool/gate_clk/mux_rmask/n1 ;
  wire   [3:0] \pool/ckg_cmask ;
  wire   [3:0] \pool/ckg_rmask ;
  wire   [10:0] \pool/pool/pe_b/peij_0_0/d_acc ;
  wire   [2:0] \pool/pool/pe_b/peij_0_0/sgnext ;
  wire   [10:0] \pool/pool/pe_b/peij_0_0/add/notb ;
  wire   [10:1] \pool/pool/pe_b/peij_0_0/add/cprop ;
  wire   [10:0] \pool/pool/pe_b/peij_0_1/d_acc ;
  wire   [2:0] \pool/pool/pe_b/peij_0_1/sgnext ;
  wire   [10:0] \pool/pool/pe_b/peij_0_1/add/notb ;
  wire   [10:1] \pool/pool/pe_b/peij_0_1/add/cprop ;
  wire   [10:0] \pool/pool/pe_b/peij_0_2/d_acc ;
  wire   [2:0] \pool/pool/pe_b/peij_0_2/sgnext ;
  wire   [10:0] \pool/pool/pe_b/peij_0_2/add/notb ;
  wire   [10:1] \pool/pool/pe_b/peij_0_2/add/cprop ;
  wire   [10:0] \pool/pool/pe_b/peij_0_3/d_acc ;
  wire   [2:0] \pool/pool/pe_b/peij_0_3/sgnext ;
  wire   [10:0] \pool/pool/pe_b/peij_0_3/add/notb ;
  wire   [10:1] \pool/pool/pe_b/peij_0_3/add/cprop ;
  wire   [10:0] \pool/pool/pe_b/peij_1_0/d_acc ;
  wire   [2:0] \pool/pool/pe_b/peij_1_0/sgnext ;
  wire   [10:0] \pool/pool/pe_b/peij_1_0/add/notb ;
  wire   [10:1] \pool/pool/pe_b/peij_1_0/add/cprop ;
  wire   [10:0] \pool/pool/pe_b/peij_1_1/d_acc ;
  wire   [2:0] \pool/pool/pe_b/peij_1_1/sgnext ;
  wire   [10:0] \pool/pool/pe_b/peij_1_1/add/notb ;
  wire   [10:1] \pool/pool/pe_b/peij_1_1/add/cprop ;
  wire   [10:0] \pool/pool/pe_b/peij_1_2/d_acc ;
  wire   [2:0] \pool/pool/pe_b/peij_1_2/sgnext ;
  wire   [10:0] \pool/pool/pe_b/peij_1_2/add/notb ;
  wire   [10:1] \pool/pool/pe_b/peij_1_2/add/cprop ;
  wire   [10:0] \pool/pool/pe_b/peij_1_3/d_acc ;
  wire   [2:0] \pool/pool/pe_b/peij_1_3/sgnext ;
  wire   [10:0] \pool/pool/pe_b/peij_1_3/add/notb ;
  wire   [10:1] \pool/pool/pe_b/peij_1_3/add/cprop ;
  wire   [10:0] \pool/pool/pe_b/peij_2_0/d_acc ;
  wire   [2:0] \pool/pool/pe_b/peij_2_0/sgnext ;
  wire   [10:0] \pool/pool/pe_b/peij_2_0/add/notb ;
  wire   [10:1] \pool/pool/pe_b/peij_2_0/add/cprop ;
  wire   [10:0] \pool/pool/pe_b/peij_2_1/d_acc ;
  wire   [2:0] \pool/pool/pe_b/peij_2_1/sgnext ;
  wire   [10:0] \pool/pool/pe_b/peij_2_1/add/notb ;
  wire   [10:1] \pool/pool/pe_b/peij_2_1/add/cprop ;
  wire   [10:0] \pool/pool/pe_b/peij_2_2/d_acc ;
  wire   [2:0] \pool/pool/pe_b/peij_2_2/sgnext ;
  wire   [10:0] \pool/pool/pe_b/peij_2_2/add/notb ;
  wire   [10:1] \pool/pool/pe_b/peij_2_2/add/cprop ;
  wire   [10:0] \pool/pool/pe_b/peij_2_3/d_acc ;
  wire   [2:0] \pool/pool/pe_b/peij_2_3/sgnext ;
  wire   [10:0] \pool/pool/pe_b/peij_2_3/add/notb ;
  wire   [10:1] \pool/pool/pe_b/peij_2_3/add/cprop ;
  wire   [10:0] \pool/pool/pe_b/peij_3_0/d_acc ;
  wire   [2:0] \pool/pool/pe_b/peij_3_0/sgnext ;
  wire   [10:0] \pool/pool/pe_b/peij_3_0/add/notb ;
  wire   [10:1] \pool/pool/pe_b/peij_3_0/add/cprop ;
  wire   [10:0] \pool/pool/pe_b/peij_3_1/d_acc ;
  wire   [2:0] \pool/pool/pe_b/peij_3_1/sgnext ;
  wire   [10:0] \pool/pool/pe_b/peij_3_1/add/notb ;
  wire   [10:1] \pool/pool/pe_b/peij_3_1/add/cprop ;
  wire   [10:0] \pool/pool/pe_b/peij_3_2/d_acc ;
  wire   [2:0] \pool/pool/pe_b/peij_3_2/sgnext ;
  wire   [10:0] \pool/pool/pe_b/peij_3_2/add/notb ;
  wire   [10:1] \pool/pool/pe_b/peij_3_2/add/cprop ;
  wire   [10:0] \pool/pool/pe_b/peij_3_3/d_acc ;
  wire   [2:0] \pool/pool/pe_b/peij_3_3/sgnext ;
  wire   [10:0] \pool/pool/pe_b/peij_3_3/add/notb ;
  wire   [10:1] \pool/pool/pe_b/peij_3_3/add/cprop ;
  wire   [2:0] \pool/fsm/next_state ;
  assign o_pool_2[3] = 1'b0;
  assign o_pool_2[7] = 1'b0;
  assign o_pool_2[11] = 1'b0;
  assign o_pool_2[15] = 1'b0;
  assign o_pool_3[3] = 1'b0;
  assign o_pool_3[7] = 1'b0;
  assign o_pool_3[11] = 1'b0;
  assign o_pool_3[15] = 1'b0;
  assign o_pool_4[3] = 1'b0;
  assign o_pool_4[7] = 1'b0;
  assign o_pool_4[11] = 1'b0;
  assign o_pool_4[15] = 1'b0;
  assign o_pool_1[3] = 1'b0;
  assign o_pool_1[7] = 1'b0;
  assign o_pool_1[11] = 1'b0;
  assign o_pool_1[15] = 1'b0;

  CLKBUF_X3 \pool/pool/interface/mux_0/U41  ( .A(
        \pool/pool/interface/mux_0/n2 ), .Z(\pool/pool/interface/mux_0/n9 ) );
  CLKBUF_X3 \pool/pool/interface/mux_0/U40  ( .A(
        \pool/pool/interface/mux_0/n2 ), .Z(\pool/pool/interface/mux_0/n8 ) );
  CLKBUF_X3 \pool/pool/interface/mux_0/U39  ( .A(
        \pool/pool/interface/mux_0/n1 ), .Z(\pool/pool/interface/mux_0/n7 ) );
  CLKBUF_X3 \pool/pool/interface/mux_0/U38  ( .A(
        \pool/pool/interface/mux_0/n1 ), .Z(\pool/pool/interface/mux_0/n6 ) );
  CLKBUF_X3 \pool/pool/interface/mux_0/U37  ( .A(
        \pool/pool/interface/mux_0/n1 ), .Z(\pool/pool/interface/mux_0/n5 ) );
  INV_X1 \pool/pool/interface/mux_0/U36  ( .A(\pool/pool/interface/mux_0/n9 ), 
        .ZN(\pool/pool/interface/mux_0/n4 ) );
  CLKBUF_X3 \pool/pool/interface/mux_0/U35  ( .A(\pool/sel ), .Z(
        \pool/pool/interface/mux_0/n2 ) );
  CLKBUF_X3 \pool/pool/interface/mux_0/U34  ( .A(\pool/sel ), .Z(
        \pool/pool/interface/mux_0/n1 ) );
  INV_X4 \pool/pool/interface/mux_0/U33  ( .A(\pool/pool/interface/mux_0/n9 ), 
        .ZN(\pool/pool/interface/mux_0/n3 ) );
  INV_X2 \pool/pool/interface/mux_0/U32  ( .A(\pool/pool/interface/mux_0/n33 ), 
        .ZN(\pool/pool/pe_b_i_data[0][0] ) );
  INV_X2 \pool/pool/interface/mux_0/U31  ( .A(\pool/pool/interface/mux_0/n32 ), 
        .ZN(\pool/pool/pe_b_i_data[0][10] ) );
  INV_X2 \pool/pool/interface/mux_0/U30  ( .A(\pool/pool/interface/mux_0/n31 ), 
        .ZN(\pool/pool/pe_b_i_data[0][11] ) );
  INV_X2 \pool/pool/interface/mux_0/U29  ( .A(\pool/pool/interface/mux_0/n30 ), 
        .ZN(\pool/pool/pe_b_i_data[0][12] ) );
  INV_X2 \pool/pool/interface/mux_0/U28  ( .A(\pool/pool/interface/mux_0/n29 ), 
        .ZN(\pool/pool/pe_b_i_data[0][13] ) );
  INV_X2 \pool/pool/interface/mux_0/U27  ( .A(\pool/pool/interface/mux_0/n28 ), 
        .ZN(\pool/pool/pe_b_i_data[0][14] ) );
  INV_X2 \pool/pool/interface/mux_0/U26  ( .A(\pool/pool/interface/mux_0/n27 ), 
        .ZN(\pool/pool/pe_b_i_data[0][15] ) );
  INV_X2 \pool/pool/interface/mux_0/U25  ( .A(\pool/pool/interface/mux_0/n26 ), 
        .ZN(\pool/pool/pe_b_i_data[0][1] ) );
  INV_X2 \pool/pool/interface/mux_0/U24  ( .A(\pool/pool/interface/mux_0/n25 ), 
        .ZN(\pool/pool/pe_b_i_data[0][2] ) );
  INV_X2 \pool/pool/interface/mux_0/U23  ( .A(\pool/pool/interface/mux_0/n24 ), 
        .ZN(\pool/pool/pe_b_i_data[0][3] ) );
  INV_X2 \pool/pool/interface/mux_0/U22  ( .A(\pool/pool/interface/mux_0/n23 ), 
        .ZN(\pool/pool/pe_b_i_data[0][4] ) );
  INV_X2 \pool/pool/interface/mux_0/U21  ( .A(\pool/pool/interface/mux_0/n22 ), 
        .ZN(\pool/pool/pe_b_i_data[0][5] ) );
  INV_X2 \pool/pool/interface/mux_0/U20  ( .A(\pool/pool/interface/mux_0/n21 ), 
        .ZN(\pool/pool/pe_b_i_data[0][6] ) );
  INV_X2 \pool/pool/interface/mux_0/U19  ( .A(\pool/pool/interface/mux_0/n20 ), 
        .ZN(\pool/pool/pe_b_i_data[0][7] ) );
  INV_X2 \pool/pool/interface/mux_0/U18  ( .A(\pool/pool/interface/mux_0/n19 ), 
        .ZN(\pool/pool/pe_b_i_data[0][8] ) );
  INV_X2 \pool/pool/interface/mux_0/U17  ( .A(\pool/pool/interface/mux_0/n18 ), 
        .ZN(\pool/pool/pe_b_i_data[0][9] ) );
  AOI22_X2 \pool/pool/interface/mux_0/U16  ( .A1(d_0[0]), .A2(
        \pool/pool/interface/mux_0/n3 ), .B1(d_4[0]), .B2(
        \pool/pool/interface/mux_0/n8 ), .ZN(\pool/pool/interface/mux_0/n33 )
         );
  AOI22_X2 \pool/pool/interface/mux_0/U15  ( .A1(d_0[10]), .A2(
        \pool/pool/interface/mux_0/n3 ), .B1(d_4[10]), .B2(
        \pool/pool/interface/mux_0/n8 ), .ZN(\pool/pool/interface/mux_0/n32 )
         );
  AOI22_X2 \pool/pool/interface/mux_0/U14  ( .A1(d_0[11]), .A2(
        \pool/pool/interface/mux_0/n3 ), .B1(d_4[11]), .B2(
        \pool/pool/interface/mux_0/n8 ), .ZN(\pool/pool/interface/mux_0/n31 )
         );
  AOI22_X2 \pool/pool/interface/mux_0/U13  ( .A1(d_0[12]), .A2(
        \pool/pool/interface/mux_0/n3 ), .B1(d_4[12]), .B2(
        \pool/pool/interface/mux_0/n7 ), .ZN(\pool/pool/interface/mux_0/n30 )
         );
  AOI22_X2 \pool/pool/interface/mux_0/U12  ( .A1(d_0[13]), .A2(
        \pool/pool/interface/mux_0/n3 ), .B1(d_4[13]), .B2(
        \pool/pool/interface/mux_0/n7 ), .ZN(\pool/pool/interface/mux_0/n29 )
         );
  AOI22_X2 \pool/pool/interface/mux_0/U11  ( .A1(d_0[14]), .A2(
        \pool/pool/interface/mux_0/n3 ), .B1(d_4[14]), .B2(
        \pool/pool/interface/mux_0/n7 ), .ZN(\pool/pool/interface/mux_0/n28 )
         );
  AOI22_X2 \pool/pool/interface/mux_0/U10  ( .A1(d_0[15]), .A2(
        \pool/pool/interface/mux_0/n3 ), .B1(d_4[15]), .B2(
        \pool/pool/interface/mux_0/n6 ), .ZN(\pool/pool/interface/mux_0/n27 )
         );
  AOI22_X2 \pool/pool/interface/mux_0/U9  ( .A1(d_0[1]), .A2(
        \pool/pool/interface/mux_0/n3 ), .B1(d_4[1]), .B2(
        \pool/pool/interface/mux_0/n6 ), .ZN(\pool/pool/interface/mux_0/n26 )
         );
  AOI22_X2 \pool/pool/interface/mux_0/U8  ( .A1(d_0[2]), .A2(
        \pool/pool/interface/mux_0/n3 ), .B1(d_4[2]), .B2(
        \pool/pool/interface/mux_0/n6 ), .ZN(\pool/pool/interface/mux_0/n25 )
         );
  AOI22_X2 \pool/pool/interface/mux_0/U7  ( .A1(d_0[3]), .A2(
        \pool/pool/interface/mux_0/n3 ), .B1(d_4[3]), .B2(
        \pool/pool/interface/mux_0/n6 ), .ZN(\pool/pool/interface/mux_0/n24 )
         );
  AOI22_X2 \pool/pool/interface/mux_0/U6  ( .A1(d_0[4]), .A2(
        \pool/pool/interface/mux_0/n3 ), .B1(d_4[4]), .B2(
        \pool/pool/interface/mux_0/n5 ), .ZN(\pool/pool/interface/mux_0/n23 )
         );
  AOI22_X2 \pool/pool/interface/mux_0/U5  ( .A1(d_0[5]), .A2(
        \pool/pool/interface/mux_0/n3 ), .B1(d_4[5]), .B2(
        \pool/pool/interface/mux_0/n7 ), .ZN(\pool/pool/interface/mux_0/n22 )
         );
  AOI22_X2 \pool/pool/interface/mux_0/U4  ( .A1(d_0[6]), .A2(
        \pool/pool/interface/mux_0/n4 ), .B1(d_4[6]), .B2(
        \pool/pool/interface/mux_0/n5 ), .ZN(\pool/pool/interface/mux_0/n21 )
         );
  AOI22_X2 \pool/pool/interface/mux_0/U3  ( .A1(d_0[7]), .A2(
        \pool/pool/interface/mux_0/n4 ), .B1(d_4[7]), .B2(
        \pool/pool/interface/mux_0/n5 ), .ZN(\pool/pool/interface/mux_0/n20 )
         );
  AOI22_X2 \pool/pool/interface/mux_0/U2  ( .A1(d_0[8]), .A2(
        \pool/pool/interface/mux_0/n4 ), .B1(d_4[8]), .B2(
        \pool/pool/interface/mux_0/n5 ), .ZN(\pool/pool/interface/mux_0/n19 )
         );
  AOI22_X2 \pool/pool/interface/mux_0/U1  ( .A1(d_0[9]), .A2(
        \pool/pool/interface/mux_0/n4 ), .B1(\pool/pool/interface/mux_0/n8 ), 
        .B2(d_4[9]), .ZN(\pool/pool/interface/mux_0/n18 ) );
  CLKBUF_X3 \pool/pool/interface/mux_1/U41  ( .A(
        \pool/pool/interface/mux_1/n2 ), .Z(\pool/pool/interface/mux_1/n9 ) );
  CLKBUF_X3 \pool/pool/interface/mux_1/U40  ( .A(
        \pool/pool/interface/mux_1/n2 ), .Z(\pool/pool/interface/mux_1/n8 ) );
  CLKBUF_X3 \pool/pool/interface/mux_1/U39  ( .A(
        \pool/pool/interface/mux_1/n1 ), .Z(\pool/pool/interface/mux_1/n7 ) );
  CLKBUF_X3 \pool/pool/interface/mux_1/U38  ( .A(
        \pool/pool/interface/mux_1/n1 ), .Z(\pool/pool/interface/mux_1/n6 ) );
  CLKBUF_X3 \pool/pool/interface/mux_1/U37  ( .A(
        \pool/pool/interface/mux_1/n1 ), .Z(\pool/pool/interface/mux_1/n5 ) );
  INV_X1 \pool/pool/interface/mux_1/U36  ( .A(\pool/pool/interface/mux_1/n9 ), 
        .ZN(\pool/pool/interface/mux_1/n4 ) );
  CLKBUF_X3 \pool/pool/interface/mux_1/U35  ( .A(\pool/sel ), .Z(
        \pool/pool/interface/mux_1/n2 ) );
  CLKBUF_X3 \pool/pool/interface/mux_1/U34  ( .A(\pool/sel ), .Z(
        \pool/pool/interface/mux_1/n1 ) );
  INV_X4 \pool/pool/interface/mux_1/U33  ( .A(\pool/pool/interface/mux_1/n9 ), 
        .ZN(\pool/pool/interface/mux_1/n3 ) );
  INV_X2 \pool/pool/interface/mux_1/U32  ( .A(\pool/pool/interface/mux_1/n10 ), 
        .ZN(\pool/pool/pe_b_i_data[1][0] ) );
  INV_X2 \pool/pool/interface/mux_1/U31  ( .A(\pool/pool/interface/mux_1/n11 ), 
        .ZN(\pool/pool/pe_b_i_data[1][10] ) );
  INV_X2 \pool/pool/interface/mux_1/U30  ( .A(\pool/pool/interface/mux_1/n12 ), 
        .ZN(\pool/pool/pe_b_i_data[1][11] ) );
  INV_X2 \pool/pool/interface/mux_1/U29  ( .A(\pool/pool/interface/mux_1/n13 ), 
        .ZN(\pool/pool/pe_b_i_data[1][12] ) );
  INV_X2 \pool/pool/interface/mux_1/U28  ( .A(\pool/pool/interface/mux_1/n14 ), 
        .ZN(\pool/pool/pe_b_i_data[1][13] ) );
  INV_X2 \pool/pool/interface/mux_1/U27  ( .A(\pool/pool/interface/mux_1/n15 ), 
        .ZN(\pool/pool/pe_b_i_data[1][14] ) );
  INV_X2 \pool/pool/interface/mux_1/U26  ( .A(\pool/pool/interface/mux_1/n16 ), 
        .ZN(\pool/pool/pe_b_i_data[1][15] ) );
  INV_X2 \pool/pool/interface/mux_1/U25  ( .A(\pool/pool/interface/mux_1/n17 ), 
        .ZN(\pool/pool/pe_b_i_data[1][1] ) );
  INV_X2 \pool/pool/interface/mux_1/U24  ( .A(\pool/pool/interface/mux_1/n26 ), 
        .ZN(\pool/pool/pe_b_i_data[1][2] ) );
  INV_X2 \pool/pool/interface/mux_1/U23  ( .A(\pool/pool/interface/mux_1/n27 ), 
        .ZN(\pool/pool/pe_b_i_data[1][3] ) );
  INV_X2 \pool/pool/interface/mux_1/U22  ( .A(\pool/pool/interface/mux_1/n28 ), 
        .ZN(\pool/pool/pe_b_i_data[1][4] ) );
  INV_X2 \pool/pool/interface/mux_1/U21  ( .A(\pool/pool/interface/mux_1/n29 ), 
        .ZN(\pool/pool/pe_b_i_data[1][5] ) );
  INV_X2 \pool/pool/interface/mux_1/U20  ( .A(\pool/pool/interface/mux_1/n30 ), 
        .ZN(\pool/pool/pe_b_i_data[1][6] ) );
  INV_X2 \pool/pool/interface/mux_1/U19  ( .A(\pool/pool/interface/mux_1/n31 ), 
        .ZN(\pool/pool/pe_b_i_data[1][7] ) );
  INV_X2 \pool/pool/interface/mux_1/U18  ( .A(\pool/pool/interface/mux_1/n32 ), 
        .ZN(\pool/pool/pe_b_i_data[1][8] ) );
  INV_X2 \pool/pool/interface/mux_1/U17  ( .A(\pool/pool/interface/mux_1/n33 ), 
        .ZN(\pool/pool/pe_b_i_data[1][9] ) );
  AOI22_X2 \pool/pool/interface/mux_1/U16  ( .A1(d_1[0]), .A2(
        \pool/pool/interface/mux_1/n3 ), .B1(d_5[0]), .B2(
        \pool/pool/interface/mux_1/n8 ), .ZN(\pool/pool/interface/mux_1/n10 )
         );
  AOI22_X2 \pool/pool/interface/mux_1/U15  ( .A1(d_1[10]), .A2(
        \pool/pool/interface/mux_1/n3 ), .B1(d_5[10]), .B2(
        \pool/pool/interface/mux_1/n8 ), .ZN(\pool/pool/interface/mux_1/n11 )
         );
  AOI22_X2 \pool/pool/interface/mux_1/U14  ( .A1(d_1[11]), .A2(
        \pool/pool/interface/mux_1/n3 ), .B1(d_5[11]), .B2(
        \pool/pool/interface/mux_1/n8 ), .ZN(\pool/pool/interface/mux_1/n12 )
         );
  AOI22_X2 \pool/pool/interface/mux_1/U13  ( .A1(d_1[12]), .A2(
        \pool/pool/interface/mux_1/n3 ), .B1(d_5[12]), .B2(
        \pool/pool/interface/mux_1/n7 ), .ZN(\pool/pool/interface/mux_1/n13 )
         );
  AOI22_X2 \pool/pool/interface/mux_1/U12  ( .A1(d_1[13]), .A2(
        \pool/pool/interface/mux_1/n3 ), .B1(d_5[13]), .B2(
        \pool/pool/interface/mux_1/n7 ), .ZN(\pool/pool/interface/mux_1/n14 )
         );
  AOI22_X2 \pool/pool/interface/mux_1/U11  ( .A1(d_1[14]), .A2(
        \pool/pool/interface/mux_1/n3 ), .B1(d_5[14]), .B2(
        \pool/pool/interface/mux_1/n7 ), .ZN(\pool/pool/interface/mux_1/n15 )
         );
  AOI22_X2 \pool/pool/interface/mux_1/U10  ( .A1(d_1[15]), .A2(
        \pool/pool/interface/mux_1/n3 ), .B1(d_5[15]), .B2(
        \pool/pool/interface/mux_1/n6 ), .ZN(\pool/pool/interface/mux_1/n16 )
         );
  AOI22_X2 \pool/pool/interface/mux_1/U9  ( .A1(d_1[1]), .A2(
        \pool/pool/interface/mux_1/n3 ), .B1(d_5[1]), .B2(
        \pool/pool/interface/mux_1/n6 ), .ZN(\pool/pool/interface/mux_1/n17 )
         );
  AOI22_X2 \pool/pool/interface/mux_1/U8  ( .A1(d_1[2]), .A2(
        \pool/pool/interface/mux_1/n3 ), .B1(d_5[2]), .B2(
        \pool/pool/interface/mux_1/n6 ), .ZN(\pool/pool/interface/mux_1/n26 )
         );
  AOI22_X2 \pool/pool/interface/mux_1/U7  ( .A1(d_1[3]), .A2(
        \pool/pool/interface/mux_1/n3 ), .B1(d_5[3]), .B2(
        \pool/pool/interface/mux_1/n6 ), .ZN(\pool/pool/interface/mux_1/n27 )
         );
  AOI22_X2 \pool/pool/interface/mux_1/U6  ( .A1(d_1[4]), .A2(
        \pool/pool/interface/mux_1/n3 ), .B1(d_5[4]), .B2(
        \pool/pool/interface/mux_1/n5 ), .ZN(\pool/pool/interface/mux_1/n28 )
         );
  AOI22_X2 \pool/pool/interface/mux_1/U5  ( .A1(d_1[5]), .A2(
        \pool/pool/interface/mux_1/n3 ), .B1(d_5[5]), .B2(
        \pool/pool/interface/mux_1/n7 ), .ZN(\pool/pool/interface/mux_1/n29 )
         );
  AOI22_X2 \pool/pool/interface/mux_1/U4  ( .A1(d_1[6]), .A2(
        \pool/pool/interface/mux_1/n4 ), .B1(d_5[6]), .B2(
        \pool/pool/interface/mux_1/n5 ), .ZN(\pool/pool/interface/mux_1/n30 )
         );
  AOI22_X2 \pool/pool/interface/mux_1/U3  ( .A1(d_1[7]), .A2(
        \pool/pool/interface/mux_1/n4 ), .B1(d_5[7]), .B2(
        \pool/pool/interface/mux_1/n5 ), .ZN(\pool/pool/interface/mux_1/n31 )
         );
  AOI22_X2 \pool/pool/interface/mux_1/U2  ( .A1(d_1[8]), .A2(
        \pool/pool/interface/mux_1/n4 ), .B1(d_5[8]), .B2(
        \pool/pool/interface/mux_1/n5 ), .ZN(\pool/pool/interface/mux_1/n32 )
         );
  AOI22_X2 \pool/pool/interface/mux_1/U1  ( .A1(d_1[9]), .A2(
        \pool/pool/interface/mux_1/n4 ), .B1(\pool/pool/interface/mux_1/n8 ), 
        .B2(d_5[9]), .ZN(\pool/pool/interface/mux_1/n33 ) );
  CLKBUF_X3 \pool/pool/interface/mux_2/U41  ( .A(
        \pool/pool/interface/mux_2/n2 ), .Z(\pool/pool/interface/mux_2/n9 ) );
  CLKBUF_X3 \pool/pool/interface/mux_2/U40  ( .A(
        \pool/pool/interface/mux_2/n2 ), .Z(\pool/pool/interface/mux_2/n8 ) );
  CLKBUF_X3 \pool/pool/interface/mux_2/U39  ( .A(
        \pool/pool/interface/mux_2/n1 ), .Z(\pool/pool/interface/mux_2/n7 ) );
  CLKBUF_X3 \pool/pool/interface/mux_2/U38  ( .A(
        \pool/pool/interface/mux_2/n1 ), .Z(\pool/pool/interface/mux_2/n6 ) );
  CLKBUF_X3 \pool/pool/interface/mux_2/U37  ( .A(
        \pool/pool/interface/mux_2/n1 ), .Z(\pool/pool/interface/mux_2/n5 ) );
  INV_X1 \pool/pool/interface/mux_2/U36  ( .A(\pool/pool/interface/mux_2/n9 ), 
        .ZN(\pool/pool/interface/mux_2/n4 ) );
  CLKBUF_X3 \pool/pool/interface/mux_2/U35  ( .A(\pool/sel ), .Z(
        \pool/pool/interface/mux_2/n2 ) );
  CLKBUF_X3 \pool/pool/interface/mux_2/U34  ( .A(\pool/sel ), .Z(
        \pool/pool/interface/mux_2/n1 ) );
  INV_X4 \pool/pool/interface/mux_2/U33  ( .A(\pool/pool/interface/mux_2/n9 ), 
        .ZN(\pool/pool/interface/mux_2/n3 ) );
  INV_X2 \pool/pool/interface/mux_2/U32  ( .A(\pool/pool/interface/mux_2/n10 ), 
        .ZN(\pool/pool/pe_b_i_data[2][0] ) );
  INV_X2 \pool/pool/interface/mux_2/U31  ( .A(\pool/pool/interface/mux_2/n11 ), 
        .ZN(\pool/pool/pe_b_i_data[2][10] ) );
  INV_X2 \pool/pool/interface/mux_2/U30  ( .A(\pool/pool/interface/mux_2/n12 ), 
        .ZN(\pool/pool/pe_b_i_data[2][11] ) );
  INV_X2 \pool/pool/interface/mux_2/U29  ( .A(\pool/pool/interface/mux_2/n13 ), 
        .ZN(\pool/pool/pe_b_i_data[2][12] ) );
  INV_X2 \pool/pool/interface/mux_2/U28  ( .A(\pool/pool/interface/mux_2/n14 ), 
        .ZN(\pool/pool/pe_b_i_data[2][13] ) );
  INV_X2 \pool/pool/interface/mux_2/U27  ( .A(\pool/pool/interface/mux_2/n15 ), 
        .ZN(\pool/pool/pe_b_i_data[2][14] ) );
  INV_X2 \pool/pool/interface/mux_2/U26  ( .A(\pool/pool/interface/mux_2/n16 ), 
        .ZN(\pool/pool/pe_b_i_data[2][15] ) );
  INV_X2 \pool/pool/interface/mux_2/U25  ( .A(\pool/pool/interface/mux_2/n17 ), 
        .ZN(\pool/pool/pe_b_i_data[2][1] ) );
  INV_X2 \pool/pool/interface/mux_2/U24  ( .A(\pool/pool/interface/mux_2/n26 ), 
        .ZN(\pool/pool/pe_b_i_data[2][2] ) );
  INV_X2 \pool/pool/interface/mux_2/U23  ( .A(\pool/pool/interface/mux_2/n27 ), 
        .ZN(\pool/pool/pe_b_i_data[2][3] ) );
  INV_X2 \pool/pool/interface/mux_2/U22  ( .A(\pool/pool/interface/mux_2/n28 ), 
        .ZN(\pool/pool/pe_b_i_data[2][4] ) );
  INV_X2 \pool/pool/interface/mux_2/U21  ( .A(\pool/pool/interface/mux_2/n29 ), 
        .ZN(\pool/pool/pe_b_i_data[2][5] ) );
  INV_X2 \pool/pool/interface/mux_2/U20  ( .A(\pool/pool/interface/mux_2/n30 ), 
        .ZN(\pool/pool/pe_b_i_data[2][6] ) );
  INV_X2 \pool/pool/interface/mux_2/U19  ( .A(\pool/pool/interface/mux_2/n31 ), 
        .ZN(\pool/pool/pe_b_i_data[2][7] ) );
  INV_X2 \pool/pool/interface/mux_2/U18  ( .A(\pool/pool/interface/mux_2/n32 ), 
        .ZN(\pool/pool/pe_b_i_data[2][8] ) );
  INV_X2 \pool/pool/interface/mux_2/U17  ( .A(\pool/pool/interface/mux_2/n33 ), 
        .ZN(\pool/pool/pe_b_i_data[2][9] ) );
  AOI22_X2 \pool/pool/interface/mux_2/U16  ( .A1(d_2[0]), .A2(
        \pool/pool/interface/mux_2/n3 ), .B1(d_6[0]), .B2(
        \pool/pool/interface/mux_2/n8 ), .ZN(\pool/pool/interface/mux_2/n10 )
         );
  AOI22_X2 \pool/pool/interface/mux_2/U15  ( .A1(d_2[10]), .A2(
        \pool/pool/interface/mux_2/n3 ), .B1(d_6[10]), .B2(
        \pool/pool/interface/mux_2/n8 ), .ZN(\pool/pool/interface/mux_2/n11 )
         );
  AOI22_X2 \pool/pool/interface/mux_2/U14  ( .A1(d_2[11]), .A2(
        \pool/pool/interface/mux_2/n3 ), .B1(d_6[11]), .B2(
        \pool/pool/interface/mux_2/n8 ), .ZN(\pool/pool/interface/mux_2/n12 )
         );
  AOI22_X2 \pool/pool/interface/mux_2/U13  ( .A1(d_2[12]), .A2(
        \pool/pool/interface/mux_2/n3 ), .B1(d_6[12]), .B2(
        \pool/pool/interface/mux_2/n7 ), .ZN(\pool/pool/interface/mux_2/n13 )
         );
  AOI22_X2 \pool/pool/interface/mux_2/U12  ( .A1(d_2[13]), .A2(
        \pool/pool/interface/mux_2/n3 ), .B1(d_6[13]), .B2(
        \pool/pool/interface/mux_2/n7 ), .ZN(\pool/pool/interface/mux_2/n14 )
         );
  AOI22_X2 \pool/pool/interface/mux_2/U11  ( .A1(d_2[14]), .A2(
        \pool/pool/interface/mux_2/n3 ), .B1(d_6[14]), .B2(
        \pool/pool/interface/mux_2/n7 ), .ZN(\pool/pool/interface/mux_2/n15 )
         );
  AOI22_X2 \pool/pool/interface/mux_2/U10  ( .A1(d_2[15]), .A2(
        \pool/pool/interface/mux_2/n3 ), .B1(d_6[15]), .B2(
        \pool/pool/interface/mux_2/n6 ), .ZN(\pool/pool/interface/mux_2/n16 )
         );
  AOI22_X2 \pool/pool/interface/mux_2/U9  ( .A1(d_2[1]), .A2(
        \pool/pool/interface/mux_2/n3 ), .B1(d_6[1]), .B2(
        \pool/pool/interface/mux_2/n6 ), .ZN(\pool/pool/interface/mux_2/n17 )
         );
  AOI22_X2 \pool/pool/interface/mux_2/U8  ( .A1(d_2[2]), .A2(
        \pool/pool/interface/mux_2/n3 ), .B1(d_6[2]), .B2(
        \pool/pool/interface/mux_2/n6 ), .ZN(\pool/pool/interface/mux_2/n26 )
         );
  AOI22_X2 \pool/pool/interface/mux_2/U7  ( .A1(d_2[3]), .A2(
        \pool/pool/interface/mux_2/n3 ), .B1(d_6[3]), .B2(
        \pool/pool/interface/mux_2/n6 ), .ZN(\pool/pool/interface/mux_2/n27 )
         );
  AOI22_X2 \pool/pool/interface/mux_2/U6  ( .A1(d_2[4]), .A2(
        \pool/pool/interface/mux_2/n3 ), .B1(d_6[4]), .B2(
        \pool/pool/interface/mux_2/n5 ), .ZN(\pool/pool/interface/mux_2/n28 )
         );
  AOI22_X2 \pool/pool/interface/mux_2/U5  ( .A1(d_2[5]), .A2(
        \pool/pool/interface/mux_2/n3 ), .B1(d_6[5]), .B2(
        \pool/pool/interface/mux_2/n7 ), .ZN(\pool/pool/interface/mux_2/n29 )
         );
  AOI22_X2 \pool/pool/interface/mux_2/U4  ( .A1(d_2[6]), .A2(
        \pool/pool/interface/mux_2/n4 ), .B1(d_6[6]), .B2(
        \pool/pool/interface/mux_2/n5 ), .ZN(\pool/pool/interface/mux_2/n30 )
         );
  AOI22_X2 \pool/pool/interface/mux_2/U3  ( .A1(d_2[7]), .A2(
        \pool/pool/interface/mux_2/n4 ), .B1(d_6[7]), .B2(
        \pool/pool/interface/mux_2/n5 ), .ZN(\pool/pool/interface/mux_2/n31 )
         );
  AOI22_X2 \pool/pool/interface/mux_2/U2  ( .A1(d_2[8]), .A2(
        \pool/pool/interface/mux_2/n4 ), .B1(d_6[8]), .B2(
        \pool/pool/interface/mux_2/n5 ), .ZN(\pool/pool/interface/mux_2/n32 )
         );
  AOI22_X2 \pool/pool/interface/mux_2/U1  ( .A1(d_2[9]), .A2(
        \pool/pool/interface/mux_2/n4 ), .B1(\pool/pool/interface/mux_2/n8 ), 
        .B2(d_6[9]), .ZN(\pool/pool/interface/mux_2/n33 ) );
  CLKBUF_X3 \pool/pool/interface/mux_3/U41  ( .A(
        \pool/pool/interface/mux_3/n2 ), .Z(\pool/pool/interface/mux_3/n9 ) );
  CLKBUF_X3 \pool/pool/interface/mux_3/U40  ( .A(
        \pool/pool/interface/mux_3/n2 ), .Z(\pool/pool/interface/mux_3/n8 ) );
  CLKBUF_X3 \pool/pool/interface/mux_3/U39  ( .A(
        \pool/pool/interface/mux_3/n1 ), .Z(\pool/pool/interface/mux_3/n7 ) );
  CLKBUF_X3 \pool/pool/interface/mux_3/U38  ( .A(
        \pool/pool/interface/mux_3/n1 ), .Z(\pool/pool/interface/mux_3/n6 ) );
  CLKBUF_X3 \pool/pool/interface/mux_3/U37  ( .A(
        \pool/pool/interface/mux_3/n1 ), .Z(\pool/pool/interface/mux_3/n5 ) );
  INV_X1 \pool/pool/interface/mux_3/U36  ( .A(\pool/pool/interface/mux_3/n9 ), 
        .ZN(\pool/pool/interface/mux_3/n4 ) );
  CLKBUF_X3 \pool/pool/interface/mux_3/U35  ( .A(\pool/sel ), .Z(
        \pool/pool/interface/mux_3/n2 ) );
  CLKBUF_X3 \pool/pool/interface/mux_3/U34  ( .A(\pool/sel ), .Z(
        \pool/pool/interface/mux_3/n1 ) );
  INV_X4 \pool/pool/interface/mux_3/U33  ( .A(\pool/pool/interface/mux_3/n9 ), 
        .ZN(\pool/pool/interface/mux_3/n3 ) );
  INV_X2 \pool/pool/interface/mux_3/U32  ( .A(\pool/pool/interface/mux_3/n10 ), 
        .ZN(\pool/pool/pe_b_i_data[3][0] ) );
  INV_X2 \pool/pool/interface/mux_3/U31  ( .A(\pool/pool/interface/mux_3/n11 ), 
        .ZN(\pool/pool/pe_b_i_data[3][10] ) );
  INV_X2 \pool/pool/interface/mux_3/U30  ( .A(\pool/pool/interface/mux_3/n12 ), 
        .ZN(\pool/pool/pe_b_i_data[3][11] ) );
  INV_X2 \pool/pool/interface/mux_3/U29  ( .A(\pool/pool/interface/mux_3/n13 ), 
        .ZN(\pool/pool/pe_b_i_data[3][12] ) );
  INV_X2 \pool/pool/interface/mux_3/U28  ( .A(\pool/pool/interface/mux_3/n14 ), 
        .ZN(\pool/pool/pe_b_i_data[3][13] ) );
  INV_X2 \pool/pool/interface/mux_3/U27  ( .A(\pool/pool/interface/mux_3/n15 ), 
        .ZN(\pool/pool/pe_b_i_data[3][14] ) );
  INV_X2 \pool/pool/interface/mux_3/U26  ( .A(\pool/pool/interface/mux_3/n16 ), 
        .ZN(\pool/pool/pe_b_i_data[3][15] ) );
  INV_X2 \pool/pool/interface/mux_3/U25  ( .A(\pool/pool/interface/mux_3/n17 ), 
        .ZN(\pool/pool/pe_b_i_data[3][1] ) );
  INV_X2 \pool/pool/interface/mux_3/U24  ( .A(\pool/pool/interface/mux_3/n26 ), 
        .ZN(\pool/pool/pe_b_i_data[3][2] ) );
  INV_X2 \pool/pool/interface/mux_3/U23  ( .A(\pool/pool/interface/mux_3/n27 ), 
        .ZN(\pool/pool/pe_b_i_data[3][3] ) );
  INV_X2 \pool/pool/interface/mux_3/U22  ( .A(\pool/pool/interface/mux_3/n28 ), 
        .ZN(\pool/pool/pe_b_i_data[3][4] ) );
  INV_X2 \pool/pool/interface/mux_3/U21  ( .A(\pool/pool/interface/mux_3/n29 ), 
        .ZN(\pool/pool/pe_b_i_data[3][5] ) );
  INV_X2 \pool/pool/interface/mux_3/U20  ( .A(\pool/pool/interface/mux_3/n30 ), 
        .ZN(\pool/pool/pe_b_i_data[3][6] ) );
  INV_X2 \pool/pool/interface/mux_3/U19  ( .A(\pool/pool/interface/mux_3/n31 ), 
        .ZN(\pool/pool/pe_b_i_data[3][7] ) );
  INV_X2 \pool/pool/interface/mux_3/U18  ( .A(\pool/pool/interface/mux_3/n32 ), 
        .ZN(\pool/pool/pe_b_i_data[3][8] ) );
  INV_X2 \pool/pool/interface/mux_3/U17  ( .A(\pool/pool/interface/mux_3/n33 ), 
        .ZN(\pool/pool/pe_b_i_data[3][9] ) );
  AOI22_X2 \pool/pool/interface/mux_3/U16  ( .A1(d_3[0]), .A2(
        \pool/pool/interface/mux_3/n3 ), .B1(d_7[0]), .B2(
        \pool/pool/interface/mux_3/n8 ), .ZN(\pool/pool/interface/mux_3/n10 )
         );
  AOI22_X2 \pool/pool/interface/mux_3/U15  ( .A1(d_3[10]), .A2(
        \pool/pool/interface/mux_3/n3 ), .B1(d_7[10]), .B2(
        \pool/pool/interface/mux_3/n8 ), .ZN(\pool/pool/interface/mux_3/n11 )
         );
  AOI22_X2 \pool/pool/interface/mux_3/U14  ( .A1(d_3[11]), .A2(
        \pool/pool/interface/mux_3/n3 ), .B1(d_7[11]), .B2(
        \pool/pool/interface/mux_3/n8 ), .ZN(\pool/pool/interface/mux_3/n12 )
         );
  AOI22_X2 \pool/pool/interface/mux_3/U13  ( .A1(d_3[12]), .A2(
        \pool/pool/interface/mux_3/n3 ), .B1(d_7[12]), .B2(
        \pool/pool/interface/mux_3/n7 ), .ZN(\pool/pool/interface/mux_3/n13 )
         );
  AOI22_X2 \pool/pool/interface/mux_3/U12  ( .A1(d_3[13]), .A2(
        \pool/pool/interface/mux_3/n3 ), .B1(d_7[13]), .B2(
        \pool/pool/interface/mux_3/n7 ), .ZN(\pool/pool/interface/mux_3/n14 )
         );
  AOI22_X2 \pool/pool/interface/mux_3/U11  ( .A1(d_3[14]), .A2(
        \pool/pool/interface/mux_3/n3 ), .B1(d_7[14]), .B2(
        \pool/pool/interface/mux_3/n7 ), .ZN(\pool/pool/interface/mux_3/n15 )
         );
  AOI22_X2 \pool/pool/interface/mux_3/U10  ( .A1(d_3[15]), .A2(
        \pool/pool/interface/mux_3/n3 ), .B1(d_7[15]), .B2(
        \pool/pool/interface/mux_3/n6 ), .ZN(\pool/pool/interface/mux_3/n16 )
         );
  AOI22_X2 \pool/pool/interface/mux_3/U9  ( .A1(d_3[1]), .A2(
        \pool/pool/interface/mux_3/n3 ), .B1(d_7[1]), .B2(
        \pool/pool/interface/mux_3/n6 ), .ZN(\pool/pool/interface/mux_3/n17 )
         );
  AOI22_X2 \pool/pool/interface/mux_3/U8  ( .A1(d_3[2]), .A2(
        \pool/pool/interface/mux_3/n3 ), .B1(d_7[2]), .B2(
        \pool/pool/interface/mux_3/n6 ), .ZN(\pool/pool/interface/mux_3/n26 )
         );
  AOI22_X2 \pool/pool/interface/mux_3/U7  ( .A1(d_3[3]), .A2(
        \pool/pool/interface/mux_3/n3 ), .B1(d_7[3]), .B2(
        \pool/pool/interface/mux_3/n6 ), .ZN(\pool/pool/interface/mux_3/n27 )
         );
  AOI22_X2 \pool/pool/interface/mux_3/U6  ( .A1(d_3[4]), .A2(
        \pool/pool/interface/mux_3/n3 ), .B1(d_7[4]), .B2(
        \pool/pool/interface/mux_3/n5 ), .ZN(\pool/pool/interface/mux_3/n28 )
         );
  AOI22_X2 \pool/pool/interface/mux_3/U5  ( .A1(d_3[5]), .A2(
        \pool/pool/interface/mux_3/n3 ), .B1(d_7[5]), .B2(
        \pool/pool/interface/mux_3/n7 ), .ZN(\pool/pool/interface/mux_3/n29 )
         );
  AOI22_X2 \pool/pool/interface/mux_3/U4  ( .A1(d_3[6]), .A2(
        \pool/pool/interface/mux_3/n4 ), .B1(d_7[6]), .B2(
        \pool/pool/interface/mux_3/n5 ), .ZN(\pool/pool/interface/mux_3/n30 )
         );
  AOI22_X2 \pool/pool/interface/mux_3/U3  ( .A1(d_3[7]), .A2(
        \pool/pool/interface/mux_3/n4 ), .B1(d_7[7]), .B2(
        \pool/pool/interface/mux_3/n5 ), .ZN(\pool/pool/interface/mux_3/n31 )
         );
  AOI22_X2 \pool/pool/interface/mux_3/U2  ( .A1(d_3[8]), .A2(
        \pool/pool/interface/mux_3/n4 ), .B1(d_7[8]), .B2(
        \pool/pool/interface/mux_3/n5 ), .ZN(\pool/pool/interface/mux_3/n32 )
         );
  AOI22_X2 \pool/pool/interface/mux_3/U1  ( .A1(d_3[9]), .A2(
        \pool/pool/interface/mux_3/n4 ), .B1(\pool/pool/interface/mux_3/n8 ), 
        .B2(d_7[9]), .ZN(\pool/pool/interface/mux_3/n33 ) );
  CLKBUF_X1 \pool/pool/pe_b/U23  ( .A(\pool/ld_h ), .Z(\pool/pool/pe_b/n7 ) );
  CLKBUF_X3 \pool/pool/pe_b/U22  ( .A(\pool/ld_h ), .Z(\pool/pool/pe_b/n6 ) );
  INV_X2 \pool/pool/pe_b/U21  ( .A(en), .ZN(\pool/pool/pe_b/n1 ) );
  OR2_X2 \pool/pool/pe_b/U20  ( .A1(\pool/ckg_rmask [3]), .A2(
        \pool/pool/pe_b/n1 ), .ZN(\pool/pool/pe_b/n5 ) );
  NOR2_X2 \pool/pool/pe_b/U19  ( .A1(\pool/ckg_cmask [3]), .A2(
        \pool/pool/pe_b/n5 ), .ZN(\pool/pool/pe_b/int_pe_en[0][0] ) );
  NOR2_X2 \pool/pool/pe_b/U18  ( .A1(\pool/ckg_cmask [2]), .A2(
        \pool/pool/pe_b/n5 ), .ZN(\pool/pool/pe_b/int_pe_en[0][1] ) );
  NOR2_X2 \pool/pool/pe_b/U17  ( .A1(\pool/ckg_cmask [1]), .A2(
        \pool/pool/pe_b/n5 ), .ZN(\pool/pool/pe_b/int_pe_en[0][2] ) );
  NOR2_X2 \pool/pool/pe_b/U16  ( .A1(\pool/ckg_cmask [0]), .A2(
        \pool/pool/pe_b/n5 ), .ZN(\pool/pool/pe_b/int_pe_en[0][3] ) );
  OR2_X2 \pool/pool/pe_b/U15  ( .A1(\pool/ckg_rmask [2]), .A2(
        \pool/pool/pe_b/n1 ), .ZN(\pool/pool/pe_b/n4 ) );
  NOR2_X2 \pool/pool/pe_b/U14  ( .A1(\pool/ckg_cmask [3]), .A2(
        \pool/pool/pe_b/n4 ), .ZN(\pool/pool/pe_b/int_pe_en[1][0] ) );
  NOR2_X2 \pool/pool/pe_b/U13  ( .A1(\pool/ckg_cmask [2]), .A2(
        \pool/pool/pe_b/n4 ), .ZN(\pool/pool/pe_b/int_pe_en[1][1] ) );
  NOR2_X2 \pool/pool/pe_b/U12  ( .A1(\pool/ckg_cmask [1]), .A2(
        \pool/pool/pe_b/n4 ), .ZN(\pool/pool/pe_b/int_pe_en[1][2] ) );
  NOR2_X2 \pool/pool/pe_b/U11  ( .A1(\pool/ckg_cmask [0]), .A2(
        \pool/pool/pe_b/n4 ), .ZN(\pool/pool/pe_b/int_pe_en[1][3] ) );
  OR2_X2 \pool/pool/pe_b/U10  ( .A1(\pool/ckg_rmask [1]), .A2(
        \pool/pool/pe_b/n1 ), .ZN(\pool/pool/pe_b/n3 ) );
  NOR2_X2 \pool/pool/pe_b/U9  ( .A1(\pool/ckg_cmask [3]), .A2(
        \pool/pool/pe_b/n3 ), .ZN(\pool/pool/pe_b/int_pe_en[2][0] ) );
  NOR2_X2 \pool/pool/pe_b/U8  ( .A1(\pool/ckg_cmask [2]), .A2(
        \pool/pool/pe_b/n3 ), .ZN(\pool/pool/pe_b/int_pe_en[2][1] ) );
  NOR2_X2 \pool/pool/pe_b/U7  ( .A1(\pool/ckg_cmask [1]), .A2(
        \pool/pool/pe_b/n3 ), .ZN(\pool/pool/pe_b/int_pe_en[2][2] ) );
  NOR2_X2 \pool/pool/pe_b/U6  ( .A1(\pool/ckg_cmask [0]), .A2(
        \pool/pool/pe_b/n3 ), .ZN(\pool/pool/pe_b/int_pe_en[2][3] ) );
  OR2_X2 \pool/pool/pe_b/U5  ( .A1(\pool/ckg_rmask [0]), .A2(
        \pool/pool/pe_b/n1 ), .ZN(\pool/pool/pe_b/n2 ) );
  NOR2_X2 \pool/pool/pe_b/U4  ( .A1(\pool/ckg_cmask [3]), .A2(
        \pool/pool/pe_b/n2 ), .ZN(\pool/pool/pe_b/int_pe_en[3][0] ) );
  NOR2_X2 \pool/pool/pe_b/U3  ( .A1(\pool/ckg_cmask [2]), .A2(
        \pool/pool/pe_b/n2 ), .ZN(\pool/pool/pe_b/int_pe_en[3][1] ) );
  NOR2_X2 \pool/pool/pe_b/U2  ( .A1(\pool/ckg_cmask [1]), .A2(
        \pool/pool/pe_b/n2 ), .ZN(\pool/pool/pe_b/int_pe_en[3][2] ) );
  NOR2_X2 \pool/pool/pe_b/U1  ( .A1(\pool/ckg_cmask [0]), .A2(
        \pool/pool/pe_b/n2 ), .ZN(\pool/pool/pe_b/int_pe_en[3][3] ) );
  INV_X1 \pool/pool/pe_b/peij_0_0/U22  ( .A(\pool/pool/pe_b/n7 ), .ZN(
        \pool/pool/pe_b/peij_0_0/n16 ) );
  INV_X1 \pool/pool/pe_b/peij_0_0/U14  ( .A(\pool/pool/pe_b/n7 ), .ZN(
        \pool/pool/pe_b/peij_0_0/n12 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_0/U13  ( .A1(
        \pool/pool/pe_b/peij_0_0/d_acc [0]), .A2(\pool/pool/pe_b/peij_0_0/n14 ), .ZN(\pool/pool/pe_b/peij_0_0/n11 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_0/U12  ( .A1(
        \pool/pool/pe_b/peij_0_0/d_acc [1]), .A2(\pool/pool/pe_b/peij_0_0/n14 ), .ZN(\pool/pool/pe_b/peij_0_0/n10 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_0/U11  ( .A1(
        \pool/pool/pe_b/peij_0_0/d_acc [2]), .A2(\pool/pool/pe_b/peij_0_0/n14 ), .ZN(\pool/pool/pe_b/peij_0_0/n9 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_0/U10  ( .A1(
        \pool/pool/pe_b/peij_0_0/d_acc [3]), .A2(\pool/pool/pe_b/peij_0_0/n14 ), .ZN(\pool/pool/pe_b/peij_0_0/n8 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_0/U9  ( .A1(
        \pool/pool/pe_b/peij_0_0/d_acc [4]), .A2(\pool/pool/pe_b/peij_0_0/n14 ), .ZN(\pool/pool/pe_b/peij_0_0/n7 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_0/U8  ( .A1(
        \pool/pool/pe_b/peij_0_0/d_acc [5]), .A2(\pool/pool/pe_b/peij_0_0/n14 ), .ZN(\pool/pool/pe_b/peij_0_0/n6 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_0/U7  ( .A1(
        \pool/pool/pe_b/peij_0_0/d_acc [6]), .A2(\pool/pool/pe_b/peij_0_0/n14 ), .ZN(\pool/pool/pe_b/peij_0_0/n5 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_0/U6  ( .A1(
        \pool/pool/pe_b/peij_0_0/d_acc [7]), .A2(\pool/pool/pe_b/peij_0_0/n14 ), .ZN(\pool/pool/pe_b/peij_0_0/n4 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_0/U5  ( .A1(
        \pool/pool/pe_b/peij_0_0/d_acc [8]), .A2(\pool/pool/pe_b/peij_0_0/n14 ), .ZN(\pool/pool/pe_b/peij_0_0/n3 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_0/U4  ( .A1(
        \pool/pool/pe_b/peij_0_0/d_acc [9]), .A2(\pool/pool/pe_b/peij_0_0/n14 ), .ZN(\pool/pool/pe_b/peij_0_0/n2 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_0/U3  ( .A1(
        \pool/pool/pe_b/peij_0_0/d_acc [10]), .A2(
        \pool/pool/pe_b/peij_0_0/n14 ), .ZN(\pool/pool/pe_b/peij_0_0/n1 ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_0/q_im_reg[3]  ( .D(
        \pool/pool/pe_b/peij_0_0/N36 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_0/n16 ), .Q(\pool/pool/pe_b/peij_0_0/sgnext_10 ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_0/q_im_reg[0]  ( .D(
        \pool/pool/pe_b/peij_0_0/N33 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_0/n16 ), .Q(\pool/pool/pe_b/peij_0_0/sgnext [0]) );
  DFFR_X1 \pool/pool/pe_b/peij_0_0/q_im_reg[1]  ( .D(
        \pool/pool/pe_b/peij_0_0/N34 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_0/n16 ), .Q(\pool/pool/pe_b/peij_0_0/sgnext [1]) );
  DFFR_X1 \pool/pool/pe_b/peij_0_0/q_im_reg[2]  ( .D(
        \pool/pool/pe_b/peij_0_0/N35 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_0/n16 ), .Q(\pool/pool/pe_b/peij_0_0/sgnext [2]) );
  DFFR_X1 \pool/pool/pe_b/peij_0_0/q_acc_reg[10]  ( .D(
        \pool/pool/pe_b/peij_0_0/n1 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_0/n16 ), .Q(\pool/pool/pe_b_o_data[0][43] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_0/q_acc_reg[9]  ( .D(
        \pool/pool/pe_b/peij_0_0/n2 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_0/n16 ), .Q(\pool/pool/pe_b_o_data[0][42] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_0/q_acc_reg[8]  ( .D(
        \pool/pool/pe_b/peij_0_0/n3 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_0/n16 ), .Q(\pool/pool/pe_b_o_data[0][41] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_0/q_acc_reg[7]  ( .D(
        \pool/pool/pe_b/peij_0_0/n4 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_0/n16 ), .Q(\pool/pool/pe_b_o_data[0][40] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_0/q_acc_reg[6]  ( .D(
        \pool/pool/pe_b/peij_0_0/n5 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_0/n16 ), .Q(\pool/pool/pe_b_o_data[0][39] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_0/q_acc_reg[5]  ( .D(
        \pool/pool/pe_b/peij_0_0/n6 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_0/n16 ), .Q(\pool/pool/pe_b_o_data[0][38] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_0/q_acc_reg[4]  ( .D(
        \pool/pool/pe_b/peij_0_0/n7 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_0/n16 ), .Q(\pool/pool/pe_b_o_data[0][37] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_0/q_acc_reg[3]  ( .D(
        \pool/pool/pe_b/peij_0_0/n8 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_0/n16 ), .Q(\pool/pool/pe_b_o_data[0][36] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_0/q_acc_reg[2]  ( .D(
        \pool/pool/pe_b/peij_0_0/n9 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_0/n16 ), .Q(\pool/pool/pe_b_o_data[0][35] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_0/q_acc_reg[1]  ( .D(
        \pool/pool/pe_b/peij_0_0/n10 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_0/n16 ), .Q(\pool/pool/pe_b_o_data[0][34] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_0/q_acc_reg[0]  ( .D(
        \pool/pool/pe_b/peij_0_0/n11 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_0/n16 ), .Q(\pool/pool/pe_b_o_data[0][33] ) );
  INV_X2 \pool/pool/pe_b/peij_0_0/U21  ( .A(\pool/sync_clr ), .ZN(
        \pool/pool/pe_b/peij_0_0/n14 ) );
  AND3_X2 \pool/pool/pe_b/peij_0_0/U20  ( .A1(\pool/pool/pe_b/int_pe_en[0][0] ), .A2(\pool/pool/pe_b/peij_0_0/n14 ), .A3(1'b1), .ZN(
        \pool/pool/pe_b/peij_0_0/n15 ) );
  AND2_X2 \pool/pool/pe_b/peij_0_0/U19  ( .A1(\pool/pool/pe_b_i_data[0][12] ), 
        .A2(\pool/pool/pe_b/peij_0_0/n15 ), .ZN(\pool/pool/pe_b/peij_0_0/N33 )
         );
  AND2_X2 \pool/pool/pe_b/peij_0_0/U18  ( .A1(\pool/pool/pe_b_i_data[0][13] ), 
        .A2(\pool/pool/pe_b/peij_0_0/n15 ), .ZN(\pool/pool/pe_b/peij_0_0/N34 )
         );
  AND2_X2 \pool/pool/pe_b/peij_0_0/U17  ( .A1(\pool/pool/pe_b_i_data[0][14] ), 
        .A2(\pool/pool/pe_b/peij_0_0/n15 ), .ZN(\pool/pool/pe_b/peij_0_0/N35 )
         );
  AND4_X4 \pool/pool/pe_b/peij_0_0/U16  ( .A1(1'b1), .A2(
        \pool/pool/pe_b_i_data[0][15] ), .A3(\pool/pool/pe_b/int_pe_en[0][0] ), 
        .A4(\pool/pool/pe_b/peij_0_0/n14 ), .ZN(\pool/pool/pe_b/peij_0_0/N36 )
         );
  SDFFR_X1 \pool/pool/pe_b/peij_0_0/q_k_reg  ( .D(1'b0), .SI(
        \pool/pool/pe_b/peij_0_0/n14 ), .SE(1'b0), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_0/n12 ), .Q(\pool/pool/pe_b/peij_0_0/q_k ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/U11  ( .A(
        \pool/pool/pe_b/peij_0_0/sgnext [0]), .B(\pool/pool/pe_b/peij_0_0/q_k ), .Z(\pool/pool/pe_b/peij_0_0/add/notb [0]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/U10  ( .A(
        \pool/pool/pe_b/peij_0_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_0/q_k ), .Z(\pool/pool/pe_b/peij_0_0/add/notb [10]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/U9  ( .A(
        \pool/pool/pe_b/peij_0_0/sgnext [1]), .B(\pool/pool/pe_b/peij_0_0/q_k ), .Z(\pool/pool/pe_b/peij_0_0/add/notb [1]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/U8  ( .A(
        \pool/pool/pe_b/peij_0_0/sgnext [2]), .B(\pool/pool/pe_b/peij_0_0/q_k ), .Z(\pool/pool/pe_b/peij_0_0/add/notb [2]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/U7  ( .A(
        \pool/pool/pe_b/peij_0_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_0/q_k ), .Z(\pool/pool/pe_b/peij_0_0/add/notb [3]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/U6  ( .A(
        \pool/pool/pe_b/peij_0_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_0/q_k ), .Z(\pool/pool/pe_b/peij_0_0/add/notb [4]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/U5  ( .A(
        \pool/pool/pe_b/peij_0_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_0/q_k ), .Z(\pool/pool/pe_b/peij_0_0/add/notb [5]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/U4  ( .A(
        \pool/pool/pe_b/peij_0_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_0/q_k ), .Z(\pool/pool/pe_b/peij_0_0/add/notb [6]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/U3  ( .A(
        \pool/pool/pe_b/peij_0_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_0/q_k ), .Z(\pool/pool/pe_b/peij_0_0/add/notb [7]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/U2  ( .A(
        \pool/pool/pe_b/peij_0_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_0/q_k ), .Z(\pool/pool/pe_b/peij_0_0/add/notb [8]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/U1  ( .A(
        \pool/pool/pe_b/peij_0_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_0/q_k ), .Z(\pool/pool/pe_b/peij_0_0/add/notb [9]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_0/U4  ( .A(
        \pool/pool/pe_b_o_data[0][33] ), .B(
        \pool/pool/pe_b/peij_0_0/add/notb [0]), .Z(
        \pool/pool/pe_b/peij_0_0/add/fai_0/n2 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_0/U3  ( .A(
        \pool/pool/pe_b/peij_0_0/q_k ), .B(
        \pool/pool/pe_b/peij_0_0/add/fai_0/n2 ), .Z(
        \pool/pool/pe_b/peij_0_0/d_acc [0]) );
  INV_X2 \pool/pool/pe_b/peij_0_0/add/fai_0/U2  ( .A(
        \pool/pool/pe_b/peij_0_0/add/fai_0/n3 ), .ZN(
        \pool/pool/pe_b/peij_0_0/add/cprop [1]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_0/add/fai_0/U1  ( .A1(
        \pool/pool/pe_b/peij_0_0/add/notb [0]), .A2(
        \pool/pool/pe_b_o_data[0][33] ), .B1(
        \pool/pool/pe_b/peij_0_0/add/fai_0/n2 ), .B2(
        \pool/pool/pe_b/peij_0_0/q_k ), .ZN(
        \pool/pool/pe_b/peij_0_0/add/fai_0/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_1/U4  ( .A(
        \pool/pool/pe_b_o_data[0][34] ), .B(
        \pool/pool/pe_b/peij_0_0/add/notb [1]), .Z(
        \pool/pool/pe_b/peij_0_0/add/fai_1/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_1/U3  ( .A(
        \pool/pool/pe_b/peij_0_0/add/cprop [1]), .B(
        \pool/pool/pe_b/peij_0_0/add/fai_1/n3 ), .Z(
        \pool/pool/pe_b/peij_0_0/d_acc [1]) );
  INV_X2 \pool/pool/pe_b/peij_0_0/add/fai_1/U2  ( .A(
        \pool/pool/pe_b/peij_0_0/add/fai_1/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_0/add/cprop [2]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_0/add/fai_1/U1  ( .A1(
        \pool/pool/pe_b/peij_0_0/add/notb [1]), .A2(
        \pool/pool/pe_b_o_data[0][34] ), .B1(
        \pool/pool/pe_b/peij_0_0/add/fai_1/n3 ), .B2(
        \pool/pool/pe_b/peij_0_0/add/cprop [1]), .ZN(
        \pool/pool/pe_b/peij_0_0/add/fai_1/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_2/U4  ( .A(
        \pool/pool/pe_b_o_data[0][35] ), .B(
        \pool/pool/pe_b/peij_0_0/add/notb [2]), .Z(
        \pool/pool/pe_b/peij_0_0/add/fai_2/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_2/U3  ( .A(
        \pool/pool/pe_b/peij_0_0/add/cprop [2]), .B(
        \pool/pool/pe_b/peij_0_0/add/fai_2/n3 ), .Z(
        \pool/pool/pe_b/peij_0_0/d_acc [2]) );
  INV_X2 \pool/pool/pe_b/peij_0_0/add/fai_2/U2  ( .A(
        \pool/pool/pe_b/peij_0_0/add/fai_2/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_0/add/cprop [3]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_0/add/fai_2/U1  ( .A1(
        \pool/pool/pe_b/peij_0_0/add/notb [2]), .A2(
        \pool/pool/pe_b_o_data[0][35] ), .B1(
        \pool/pool/pe_b/peij_0_0/add/fai_2/n3 ), .B2(
        \pool/pool/pe_b/peij_0_0/add/cprop [2]), .ZN(
        \pool/pool/pe_b/peij_0_0/add/fai_2/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_3/U4  ( .A(
        \pool/pool/pe_b_o_data[0][36] ), .B(
        \pool/pool/pe_b/peij_0_0/add/notb [3]), .Z(
        \pool/pool/pe_b/peij_0_0/add/fai_3/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_3/U3  ( .A(
        \pool/pool/pe_b/peij_0_0/add/cprop [3]), .B(
        \pool/pool/pe_b/peij_0_0/add/fai_3/n3 ), .Z(
        \pool/pool/pe_b/peij_0_0/d_acc [3]) );
  INV_X2 \pool/pool/pe_b/peij_0_0/add/fai_3/U2  ( .A(
        \pool/pool/pe_b/peij_0_0/add/fai_3/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_0/add/cprop [4]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_0/add/fai_3/U1  ( .A1(
        \pool/pool/pe_b/peij_0_0/add/notb [3]), .A2(
        \pool/pool/pe_b_o_data[0][36] ), .B1(
        \pool/pool/pe_b/peij_0_0/add/fai_3/n3 ), .B2(
        \pool/pool/pe_b/peij_0_0/add/cprop [3]), .ZN(
        \pool/pool/pe_b/peij_0_0/add/fai_3/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_4/U4  ( .A(
        \pool/pool/pe_b_o_data[0][37] ), .B(
        \pool/pool/pe_b/peij_0_0/add/notb [4]), .Z(
        \pool/pool/pe_b/peij_0_0/add/fai_4/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_4/U3  ( .A(
        \pool/pool/pe_b/peij_0_0/add/cprop [4]), .B(
        \pool/pool/pe_b/peij_0_0/add/fai_4/n3 ), .Z(
        \pool/pool/pe_b/peij_0_0/d_acc [4]) );
  INV_X2 \pool/pool/pe_b/peij_0_0/add/fai_4/U2  ( .A(
        \pool/pool/pe_b/peij_0_0/add/fai_4/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_0/add/cprop [5]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_0/add/fai_4/U1  ( .A1(
        \pool/pool/pe_b/peij_0_0/add/notb [4]), .A2(
        \pool/pool/pe_b_o_data[0][37] ), .B1(
        \pool/pool/pe_b/peij_0_0/add/fai_4/n3 ), .B2(
        \pool/pool/pe_b/peij_0_0/add/cprop [4]), .ZN(
        \pool/pool/pe_b/peij_0_0/add/fai_4/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_5/U4  ( .A(
        \pool/pool/pe_b_o_data[0][38] ), .B(
        \pool/pool/pe_b/peij_0_0/add/notb [5]), .Z(
        \pool/pool/pe_b/peij_0_0/add/fai_5/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_5/U3  ( .A(
        \pool/pool/pe_b/peij_0_0/add/cprop [5]), .B(
        \pool/pool/pe_b/peij_0_0/add/fai_5/n3 ), .Z(
        \pool/pool/pe_b/peij_0_0/d_acc [5]) );
  INV_X2 \pool/pool/pe_b/peij_0_0/add/fai_5/U2  ( .A(
        \pool/pool/pe_b/peij_0_0/add/fai_5/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_0/add/cprop [6]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_0/add/fai_5/U1  ( .A1(
        \pool/pool/pe_b/peij_0_0/add/notb [5]), .A2(
        \pool/pool/pe_b_o_data[0][38] ), .B1(
        \pool/pool/pe_b/peij_0_0/add/fai_5/n3 ), .B2(
        \pool/pool/pe_b/peij_0_0/add/cprop [5]), .ZN(
        \pool/pool/pe_b/peij_0_0/add/fai_5/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_6/U4  ( .A(
        \pool/pool/pe_b_o_data[0][39] ), .B(
        \pool/pool/pe_b/peij_0_0/add/notb [6]), .Z(
        \pool/pool/pe_b/peij_0_0/add/fai_6/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_6/U3  ( .A(
        \pool/pool/pe_b/peij_0_0/add/cprop [6]), .B(
        \pool/pool/pe_b/peij_0_0/add/fai_6/n3 ), .Z(
        \pool/pool/pe_b/peij_0_0/d_acc [6]) );
  INV_X2 \pool/pool/pe_b/peij_0_0/add/fai_6/U2  ( .A(
        \pool/pool/pe_b/peij_0_0/add/fai_6/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_0/add/cprop [7]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_0/add/fai_6/U1  ( .A1(
        \pool/pool/pe_b/peij_0_0/add/notb [6]), .A2(
        \pool/pool/pe_b_o_data[0][39] ), .B1(
        \pool/pool/pe_b/peij_0_0/add/fai_6/n3 ), .B2(
        \pool/pool/pe_b/peij_0_0/add/cprop [6]), .ZN(
        \pool/pool/pe_b/peij_0_0/add/fai_6/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_7/U4  ( .A(
        \pool/pool/pe_b_o_data[0][40] ), .B(
        \pool/pool/pe_b/peij_0_0/add/notb [7]), .Z(
        \pool/pool/pe_b/peij_0_0/add/fai_7/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_7/U3  ( .A(
        \pool/pool/pe_b/peij_0_0/add/cprop [7]), .B(
        \pool/pool/pe_b/peij_0_0/add/fai_7/n3 ), .Z(
        \pool/pool/pe_b/peij_0_0/d_acc [7]) );
  INV_X2 \pool/pool/pe_b/peij_0_0/add/fai_7/U2  ( .A(
        \pool/pool/pe_b/peij_0_0/add/fai_7/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_0/add/cprop [8]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_0/add/fai_7/U1  ( .A1(
        \pool/pool/pe_b/peij_0_0/add/notb [7]), .A2(
        \pool/pool/pe_b_o_data[0][40] ), .B1(
        \pool/pool/pe_b/peij_0_0/add/fai_7/n3 ), .B2(
        \pool/pool/pe_b/peij_0_0/add/cprop [7]), .ZN(
        \pool/pool/pe_b/peij_0_0/add/fai_7/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_8/U4  ( .A(
        \pool/pool/pe_b_o_data[0][41] ), .B(
        \pool/pool/pe_b/peij_0_0/add/notb [8]), .Z(
        \pool/pool/pe_b/peij_0_0/add/fai_8/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_8/U3  ( .A(
        \pool/pool/pe_b/peij_0_0/add/cprop [8]), .B(
        \pool/pool/pe_b/peij_0_0/add/fai_8/n3 ), .Z(
        \pool/pool/pe_b/peij_0_0/d_acc [8]) );
  INV_X2 \pool/pool/pe_b/peij_0_0/add/fai_8/U2  ( .A(
        \pool/pool/pe_b/peij_0_0/add/fai_8/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_0/add/cprop [9]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_0/add/fai_8/U1  ( .A1(
        \pool/pool/pe_b/peij_0_0/add/notb [8]), .A2(
        \pool/pool/pe_b_o_data[0][41] ), .B1(
        \pool/pool/pe_b/peij_0_0/add/fai_8/n3 ), .B2(
        \pool/pool/pe_b/peij_0_0/add/cprop [8]), .ZN(
        \pool/pool/pe_b/peij_0_0/add/fai_8/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_9/U4  ( .A(
        \pool/pool/pe_b_o_data[0][42] ), .B(
        \pool/pool/pe_b/peij_0_0/add/notb [9]), .Z(
        \pool/pool/pe_b/peij_0_0/add/fai_9/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_9/U3  ( .A(
        \pool/pool/pe_b/peij_0_0/add/cprop [9]), .B(
        \pool/pool/pe_b/peij_0_0/add/fai_9/n3 ), .Z(
        \pool/pool/pe_b/peij_0_0/d_acc [9]) );
  INV_X2 \pool/pool/pe_b/peij_0_0/add/fai_9/U2  ( .A(
        \pool/pool/pe_b/peij_0_0/add/fai_9/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_0/add/cprop [10]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_0/add/fai_9/U1  ( .A1(
        \pool/pool/pe_b/peij_0_0/add/notb [9]), .A2(
        \pool/pool/pe_b_o_data[0][42] ), .B1(
        \pool/pool/pe_b/peij_0_0/add/fai_9/n3 ), .B2(
        \pool/pool/pe_b/peij_0_0/add/cprop [9]), .ZN(
        \pool/pool/pe_b/peij_0_0/add/fai_9/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_10/U4  ( .A(
        \pool/pool/pe_b_o_data[0][43] ), .B(
        \pool/pool/pe_b/peij_0_0/add/notb [10]), .Z(
        \pool/pool/pe_b/peij_0_0/add/fai_10/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_0/add/fai_10/U3  ( .A(
        \pool/pool/pe_b/peij_0_0/add/cprop [10]), .B(
        \pool/pool/pe_b/peij_0_0/add/fai_10/n3 ), .Z(
        \pool/pool/pe_b/peij_0_0/d_acc [10]) );
  INV_X2 \pool/pool/pe_b/peij_0_0/add/fai_10/U2  ( .A(
        \pool/pool/pe_b/peij_0_0/add/fai_10/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_0/add/c_out ) );
  AOI22_X2 \pool/pool/pe_b/peij_0_0/add/fai_10/U1  ( .A1(
        \pool/pool/pe_b/peij_0_0/add/notb [10]), .A2(
        \pool/pool/pe_b_o_data[0][43] ), .B1(
        \pool/pool/pe_b/peij_0_0/add/fai_10/n3 ), .B2(
        \pool/pool/pe_b/peij_0_0/add/cprop [10]), .ZN(
        \pool/pool/pe_b/peij_0_0/add/fai_10/n1 ) );
  INV_X1 \pool/pool/pe_b/peij_0_1/U22  ( .A(\pool/pool/pe_b/n6 ), .ZN(
        \pool/pool/pe_b/peij_0_1/n16 ) );
  INV_X1 \pool/pool/pe_b/peij_0_1/U14  ( .A(\pool/pool/pe_b/n6 ), .ZN(
        \pool/pool/pe_b/peij_0_1/n12 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_1/U13  ( .A1(
        \pool/pool/pe_b/peij_0_1/d_acc [0]), .A2(\pool/pool/pe_b/peij_0_1/n18 ), .ZN(\pool/pool/pe_b/peij_0_1/n11 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_1/U12  ( .A1(
        \pool/pool/pe_b/peij_0_1/d_acc [1]), .A2(\pool/pool/pe_b/peij_0_1/n18 ), .ZN(\pool/pool/pe_b/peij_0_1/n10 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_1/U11  ( .A1(
        \pool/pool/pe_b/peij_0_1/d_acc [2]), .A2(\pool/pool/pe_b/peij_0_1/n18 ), .ZN(\pool/pool/pe_b/peij_0_1/n9 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_1/U10  ( .A1(
        \pool/pool/pe_b/peij_0_1/d_acc [3]), .A2(\pool/pool/pe_b/peij_0_1/n18 ), .ZN(\pool/pool/pe_b/peij_0_1/n8 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_1/U9  ( .A1(
        \pool/pool/pe_b/peij_0_1/d_acc [4]), .A2(\pool/pool/pe_b/peij_0_1/n18 ), .ZN(\pool/pool/pe_b/peij_0_1/n7 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_1/U8  ( .A1(
        \pool/pool/pe_b/peij_0_1/d_acc [5]), .A2(\pool/pool/pe_b/peij_0_1/n18 ), .ZN(\pool/pool/pe_b/peij_0_1/n6 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_1/U7  ( .A1(
        \pool/pool/pe_b/peij_0_1/d_acc [6]), .A2(\pool/pool/pe_b/peij_0_1/n18 ), .ZN(\pool/pool/pe_b/peij_0_1/n5 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_1/U6  ( .A1(
        \pool/pool/pe_b/peij_0_1/d_acc [7]), .A2(\pool/pool/pe_b/peij_0_1/n18 ), .ZN(\pool/pool/pe_b/peij_0_1/n4 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_1/U5  ( .A1(
        \pool/pool/pe_b/peij_0_1/d_acc [8]), .A2(\pool/pool/pe_b/peij_0_1/n18 ), .ZN(\pool/pool/pe_b/peij_0_1/n3 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_1/U4  ( .A1(
        \pool/pool/pe_b/peij_0_1/d_acc [9]), .A2(\pool/pool/pe_b/peij_0_1/n18 ), .ZN(\pool/pool/pe_b/peij_0_1/n2 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_1/U3  ( .A1(
        \pool/pool/pe_b/peij_0_1/d_acc [10]), .A2(
        \pool/pool/pe_b/peij_0_1/n18 ), .ZN(\pool/pool/pe_b/peij_0_1/n1 ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_1/q_acc_reg[10]  ( .D(
        \pool/pool/pe_b/peij_0_1/n1 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_1/n16 ), .Q(\pool/pool/pe_b_o_data[0][32] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_1/q_acc_reg[9]  ( .D(
        \pool/pool/pe_b/peij_0_1/n2 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_1/n16 ), .Q(\pool/pool/pe_b_o_data[0][31] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_1/q_acc_reg[8]  ( .D(
        \pool/pool/pe_b/peij_0_1/n3 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_1/n16 ), .Q(\pool/pool/pe_b_o_data[0][30] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_1/q_acc_reg[7]  ( .D(
        \pool/pool/pe_b/peij_0_1/n4 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_1/n16 ), .Q(\pool/pool/pe_b_o_data[0][29] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_1/q_acc_reg[6]  ( .D(
        \pool/pool/pe_b/peij_0_1/n5 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_1/n16 ), .Q(\pool/pool/pe_b_o_data[0][28] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_1/q_acc_reg[5]  ( .D(
        \pool/pool/pe_b/peij_0_1/n6 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_1/n16 ), .Q(\pool/pool/pe_b_o_data[0][27] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_1/q_acc_reg[4]  ( .D(
        \pool/pool/pe_b/peij_0_1/n7 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_1/n16 ), .Q(\pool/pool/pe_b_o_data[0][26] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_1/q_acc_reg[3]  ( .D(
        \pool/pool/pe_b/peij_0_1/n8 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_1/n16 ), .Q(\pool/pool/pe_b_o_data[0][25] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_1/q_acc_reg[2]  ( .D(
        \pool/pool/pe_b/peij_0_1/n9 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_1/n16 ), .Q(\pool/pool/pe_b_o_data[0][24] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_1/q_acc_reg[1]  ( .D(
        \pool/pool/pe_b/peij_0_1/n10 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_1/n16 ), .Q(\pool/pool/pe_b_o_data[0][23] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_1/q_acc_reg[0]  ( .D(
        \pool/pool/pe_b/peij_0_1/n11 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_1/n16 ), .Q(\pool/pool/pe_b_o_data[0][22] ) );
  INV_X2 \pool/pool/pe_b/peij_0_1/U21  ( .A(\pool/sync_clr ), .ZN(
        \pool/pool/pe_b/peij_0_1/n18 ) );
  AND3_X2 \pool/pool/pe_b/peij_0_1/U20  ( .A1(\pool/pool/pe_b/int_pe_en[0][1] ), .A2(\pool/pool/pe_b/peij_0_1/n18 ), .A3(1'b1), .ZN(
        \pool/pool/pe_b/peij_0_1/n17 ) );
  AND2_X2 \pool/pool/pe_b/peij_0_1/U19  ( .A1(\pool/pool/pe_b_i_data[0][8] ), 
        .A2(\pool/pool/pe_b/peij_0_1/n17 ), .ZN(\pool/pool/pe_b/peij_0_1/N33 )
         );
  AND2_X2 \pool/pool/pe_b/peij_0_1/U18  ( .A1(\pool/pool/pe_b_i_data[0][9] ), 
        .A2(\pool/pool/pe_b/peij_0_1/n17 ), .ZN(\pool/pool/pe_b/peij_0_1/N34 )
         );
  AND2_X2 \pool/pool/pe_b/peij_0_1/U17  ( .A1(\pool/pool/pe_b_i_data[0][10] ), 
        .A2(\pool/pool/pe_b/peij_0_1/n17 ), .ZN(\pool/pool/pe_b/peij_0_1/N35 )
         );
  AND4_X4 \pool/pool/pe_b/peij_0_1/U16  ( .A1(1'b1), .A2(
        \pool/pool/pe_b_i_data[0][11] ), .A3(\pool/pool/pe_b/int_pe_en[0][1] ), 
        .A4(\pool/pool/pe_b/peij_0_1/n18 ), .ZN(\pool/pool/pe_b/peij_0_1/N36 )
         );
  DFFR_X1 \pool/pool/pe_b/peij_0_1/q_im_reg[0]  ( .D(
        \pool/pool/pe_b/peij_0_1/N33 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_1/n12 ), .Q(\pool/pool/pe_b/peij_0_1/sgnext [0]) );
  DFFR_X1 \pool/pool/pe_b/peij_0_1/q_im_reg[1]  ( .D(
        \pool/pool/pe_b/peij_0_1/N34 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_1/n12 ), .Q(\pool/pool/pe_b/peij_0_1/sgnext [1]) );
  DFFR_X1 \pool/pool/pe_b/peij_0_1/q_im_reg[2]  ( .D(
        \pool/pool/pe_b/peij_0_1/N35 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_1/n12 ), .Q(\pool/pool/pe_b/peij_0_1/sgnext [2]) );
  DFFR_X1 \pool/pool/pe_b/peij_0_1/q_im_reg[3]  ( .D(
        \pool/pool/pe_b/peij_0_1/N36 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_1/n12 ), .Q(\pool/pool/pe_b/peij_0_1/sgnext_10 ) );
  SDFFR_X1 \pool/pool/pe_b/peij_0_1/q_k_reg  ( .D(1'b0), .SI(
        \pool/pool/pe_b/peij_0_1/n18 ), .SE(1'b0), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_1/n12 ), .Q(\pool/pool/pe_b/peij_0_1/q_k ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/U11  ( .A(
        \pool/pool/pe_b/peij_0_1/sgnext [0]), .B(\pool/pool/pe_b/peij_0_1/q_k ), .Z(\pool/pool/pe_b/peij_0_1/add/notb [0]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/U10  ( .A(
        \pool/pool/pe_b/peij_0_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_1/q_k ), .Z(\pool/pool/pe_b/peij_0_1/add/notb [10]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/U9  ( .A(
        \pool/pool/pe_b/peij_0_1/sgnext [1]), .B(\pool/pool/pe_b/peij_0_1/q_k ), .Z(\pool/pool/pe_b/peij_0_1/add/notb [1]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/U8  ( .A(
        \pool/pool/pe_b/peij_0_1/sgnext [2]), .B(\pool/pool/pe_b/peij_0_1/q_k ), .Z(\pool/pool/pe_b/peij_0_1/add/notb [2]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/U7  ( .A(
        \pool/pool/pe_b/peij_0_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_1/q_k ), .Z(\pool/pool/pe_b/peij_0_1/add/notb [3]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/U6  ( .A(
        \pool/pool/pe_b/peij_0_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_1/q_k ), .Z(\pool/pool/pe_b/peij_0_1/add/notb [4]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/U5  ( .A(
        \pool/pool/pe_b/peij_0_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_1/q_k ), .Z(\pool/pool/pe_b/peij_0_1/add/notb [5]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/U4  ( .A(
        \pool/pool/pe_b/peij_0_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_1/q_k ), .Z(\pool/pool/pe_b/peij_0_1/add/notb [6]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/U3  ( .A(
        \pool/pool/pe_b/peij_0_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_1/q_k ), .Z(\pool/pool/pe_b/peij_0_1/add/notb [7]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/U2  ( .A(
        \pool/pool/pe_b/peij_0_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_1/q_k ), .Z(\pool/pool/pe_b/peij_0_1/add/notb [8]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/U1  ( .A(
        \pool/pool/pe_b/peij_0_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_1/q_k ), .Z(\pool/pool/pe_b/peij_0_1/add/notb [9]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_0/U4  ( .A(
        \pool/pool/pe_b_o_data[0][22] ), .B(
        \pool/pool/pe_b/peij_0_1/add/notb [0]), .Z(
        \pool/pool/pe_b/peij_0_1/add/fai_0/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_0/U3  ( .A(
        \pool/pool/pe_b/peij_0_1/q_k ), .B(
        \pool/pool/pe_b/peij_0_1/add/fai_0/n3 ), .Z(
        \pool/pool/pe_b/peij_0_1/d_acc [0]) );
  INV_X2 \pool/pool/pe_b/peij_0_1/add/fai_0/U2  ( .A(
        \pool/pool/pe_b/peij_0_1/add/fai_0/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_1/add/cprop [1]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_1/add/fai_0/U1  ( .A1(
        \pool/pool/pe_b/peij_0_1/add/notb [0]), .A2(
        \pool/pool/pe_b_o_data[0][22] ), .B1(
        \pool/pool/pe_b/peij_0_1/add/fai_0/n3 ), .B2(
        \pool/pool/pe_b/peij_0_1/q_k ), .ZN(
        \pool/pool/pe_b/peij_0_1/add/fai_0/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_1/U4  ( .A(
        \pool/pool/pe_b_o_data[0][23] ), .B(
        \pool/pool/pe_b/peij_0_1/add/notb [1]), .Z(
        \pool/pool/pe_b/peij_0_1/add/fai_1/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_1/U3  ( .A(
        \pool/pool/pe_b/peij_0_1/add/cprop [1]), .B(
        \pool/pool/pe_b/peij_0_1/add/fai_1/n3 ), .Z(
        \pool/pool/pe_b/peij_0_1/d_acc [1]) );
  INV_X2 \pool/pool/pe_b/peij_0_1/add/fai_1/U2  ( .A(
        \pool/pool/pe_b/peij_0_1/add/fai_1/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_1/add/cprop [2]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_1/add/fai_1/U1  ( .A1(
        \pool/pool/pe_b/peij_0_1/add/notb [1]), .A2(
        \pool/pool/pe_b_o_data[0][23] ), .B1(
        \pool/pool/pe_b/peij_0_1/add/fai_1/n3 ), .B2(
        \pool/pool/pe_b/peij_0_1/add/cprop [1]), .ZN(
        \pool/pool/pe_b/peij_0_1/add/fai_1/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_2/U4  ( .A(
        \pool/pool/pe_b_o_data[0][24] ), .B(
        \pool/pool/pe_b/peij_0_1/add/notb [2]), .Z(
        \pool/pool/pe_b/peij_0_1/add/fai_2/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_2/U3  ( .A(
        \pool/pool/pe_b/peij_0_1/add/cprop [2]), .B(
        \pool/pool/pe_b/peij_0_1/add/fai_2/n3 ), .Z(
        \pool/pool/pe_b/peij_0_1/d_acc [2]) );
  INV_X2 \pool/pool/pe_b/peij_0_1/add/fai_2/U2  ( .A(
        \pool/pool/pe_b/peij_0_1/add/fai_2/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_1/add/cprop [3]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_1/add/fai_2/U1  ( .A1(
        \pool/pool/pe_b/peij_0_1/add/notb [2]), .A2(
        \pool/pool/pe_b_o_data[0][24] ), .B1(
        \pool/pool/pe_b/peij_0_1/add/fai_2/n3 ), .B2(
        \pool/pool/pe_b/peij_0_1/add/cprop [2]), .ZN(
        \pool/pool/pe_b/peij_0_1/add/fai_2/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_3/U4  ( .A(
        \pool/pool/pe_b_o_data[0][25] ), .B(
        \pool/pool/pe_b/peij_0_1/add/notb [3]), .Z(
        \pool/pool/pe_b/peij_0_1/add/fai_3/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_3/U3  ( .A(
        \pool/pool/pe_b/peij_0_1/add/cprop [3]), .B(
        \pool/pool/pe_b/peij_0_1/add/fai_3/n3 ), .Z(
        \pool/pool/pe_b/peij_0_1/d_acc [3]) );
  INV_X2 \pool/pool/pe_b/peij_0_1/add/fai_3/U2  ( .A(
        \pool/pool/pe_b/peij_0_1/add/fai_3/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_1/add/cprop [4]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_1/add/fai_3/U1  ( .A1(
        \pool/pool/pe_b/peij_0_1/add/notb [3]), .A2(
        \pool/pool/pe_b_o_data[0][25] ), .B1(
        \pool/pool/pe_b/peij_0_1/add/fai_3/n3 ), .B2(
        \pool/pool/pe_b/peij_0_1/add/cprop [3]), .ZN(
        \pool/pool/pe_b/peij_0_1/add/fai_3/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_4/U4  ( .A(
        \pool/pool/pe_b_o_data[0][26] ), .B(
        \pool/pool/pe_b/peij_0_1/add/notb [4]), .Z(
        \pool/pool/pe_b/peij_0_1/add/fai_4/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_4/U3  ( .A(
        \pool/pool/pe_b/peij_0_1/add/cprop [4]), .B(
        \pool/pool/pe_b/peij_0_1/add/fai_4/n3 ), .Z(
        \pool/pool/pe_b/peij_0_1/d_acc [4]) );
  INV_X2 \pool/pool/pe_b/peij_0_1/add/fai_4/U2  ( .A(
        \pool/pool/pe_b/peij_0_1/add/fai_4/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_1/add/cprop [5]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_1/add/fai_4/U1  ( .A1(
        \pool/pool/pe_b/peij_0_1/add/notb [4]), .A2(
        \pool/pool/pe_b_o_data[0][26] ), .B1(
        \pool/pool/pe_b/peij_0_1/add/fai_4/n3 ), .B2(
        \pool/pool/pe_b/peij_0_1/add/cprop [4]), .ZN(
        \pool/pool/pe_b/peij_0_1/add/fai_4/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_5/U4  ( .A(
        \pool/pool/pe_b_o_data[0][27] ), .B(
        \pool/pool/pe_b/peij_0_1/add/notb [5]), .Z(
        \pool/pool/pe_b/peij_0_1/add/fai_5/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_5/U3  ( .A(
        \pool/pool/pe_b/peij_0_1/add/cprop [5]), .B(
        \pool/pool/pe_b/peij_0_1/add/fai_5/n3 ), .Z(
        \pool/pool/pe_b/peij_0_1/d_acc [5]) );
  INV_X2 \pool/pool/pe_b/peij_0_1/add/fai_5/U2  ( .A(
        \pool/pool/pe_b/peij_0_1/add/fai_5/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_1/add/cprop [6]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_1/add/fai_5/U1  ( .A1(
        \pool/pool/pe_b/peij_0_1/add/notb [5]), .A2(
        \pool/pool/pe_b_o_data[0][27] ), .B1(
        \pool/pool/pe_b/peij_0_1/add/fai_5/n3 ), .B2(
        \pool/pool/pe_b/peij_0_1/add/cprop [5]), .ZN(
        \pool/pool/pe_b/peij_0_1/add/fai_5/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_6/U4  ( .A(
        \pool/pool/pe_b_o_data[0][28] ), .B(
        \pool/pool/pe_b/peij_0_1/add/notb [6]), .Z(
        \pool/pool/pe_b/peij_0_1/add/fai_6/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_6/U3  ( .A(
        \pool/pool/pe_b/peij_0_1/add/cprop [6]), .B(
        \pool/pool/pe_b/peij_0_1/add/fai_6/n3 ), .Z(
        \pool/pool/pe_b/peij_0_1/d_acc [6]) );
  INV_X2 \pool/pool/pe_b/peij_0_1/add/fai_6/U2  ( .A(
        \pool/pool/pe_b/peij_0_1/add/fai_6/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_1/add/cprop [7]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_1/add/fai_6/U1  ( .A1(
        \pool/pool/pe_b/peij_0_1/add/notb [6]), .A2(
        \pool/pool/pe_b_o_data[0][28] ), .B1(
        \pool/pool/pe_b/peij_0_1/add/fai_6/n3 ), .B2(
        \pool/pool/pe_b/peij_0_1/add/cprop [6]), .ZN(
        \pool/pool/pe_b/peij_0_1/add/fai_6/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_7/U4  ( .A(
        \pool/pool/pe_b_o_data[0][29] ), .B(
        \pool/pool/pe_b/peij_0_1/add/notb [7]), .Z(
        \pool/pool/pe_b/peij_0_1/add/fai_7/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_7/U3  ( .A(
        \pool/pool/pe_b/peij_0_1/add/cprop [7]), .B(
        \pool/pool/pe_b/peij_0_1/add/fai_7/n3 ), .Z(
        \pool/pool/pe_b/peij_0_1/d_acc [7]) );
  INV_X2 \pool/pool/pe_b/peij_0_1/add/fai_7/U2  ( .A(
        \pool/pool/pe_b/peij_0_1/add/fai_7/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_1/add/cprop [8]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_1/add/fai_7/U1  ( .A1(
        \pool/pool/pe_b/peij_0_1/add/notb [7]), .A2(
        \pool/pool/pe_b_o_data[0][29] ), .B1(
        \pool/pool/pe_b/peij_0_1/add/fai_7/n3 ), .B2(
        \pool/pool/pe_b/peij_0_1/add/cprop [7]), .ZN(
        \pool/pool/pe_b/peij_0_1/add/fai_7/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_8/U4  ( .A(
        \pool/pool/pe_b_o_data[0][30] ), .B(
        \pool/pool/pe_b/peij_0_1/add/notb [8]), .Z(
        \pool/pool/pe_b/peij_0_1/add/fai_8/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_8/U3  ( .A(
        \pool/pool/pe_b/peij_0_1/add/cprop [8]), .B(
        \pool/pool/pe_b/peij_0_1/add/fai_8/n3 ), .Z(
        \pool/pool/pe_b/peij_0_1/d_acc [8]) );
  INV_X2 \pool/pool/pe_b/peij_0_1/add/fai_8/U2  ( .A(
        \pool/pool/pe_b/peij_0_1/add/fai_8/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_1/add/cprop [9]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_1/add/fai_8/U1  ( .A1(
        \pool/pool/pe_b/peij_0_1/add/notb [8]), .A2(
        \pool/pool/pe_b_o_data[0][30] ), .B1(
        \pool/pool/pe_b/peij_0_1/add/fai_8/n3 ), .B2(
        \pool/pool/pe_b/peij_0_1/add/cprop [8]), .ZN(
        \pool/pool/pe_b/peij_0_1/add/fai_8/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_9/U4  ( .A(
        \pool/pool/pe_b_o_data[0][31] ), .B(
        \pool/pool/pe_b/peij_0_1/add/notb [9]), .Z(
        \pool/pool/pe_b/peij_0_1/add/fai_9/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_9/U3  ( .A(
        \pool/pool/pe_b/peij_0_1/add/cprop [9]), .B(
        \pool/pool/pe_b/peij_0_1/add/fai_9/n3 ), .Z(
        \pool/pool/pe_b/peij_0_1/d_acc [9]) );
  INV_X2 \pool/pool/pe_b/peij_0_1/add/fai_9/U2  ( .A(
        \pool/pool/pe_b/peij_0_1/add/fai_9/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_1/add/cprop [10]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_1/add/fai_9/U1  ( .A1(
        \pool/pool/pe_b/peij_0_1/add/notb [9]), .A2(
        \pool/pool/pe_b_o_data[0][31] ), .B1(
        \pool/pool/pe_b/peij_0_1/add/fai_9/n3 ), .B2(
        \pool/pool/pe_b/peij_0_1/add/cprop [9]), .ZN(
        \pool/pool/pe_b/peij_0_1/add/fai_9/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_10/U4  ( .A(
        \pool/pool/pe_b_o_data[0][32] ), .B(
        \pool/pool/pe_b/peij_0_1/add/notb [10]), .Z(
        \pool/pool/pe_b/peij_0_1/add/fai_10/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_1/add/fai_10/U3  ( .A(
        \pool/pool/pe_b/peij_0_1/add/cprop [10]), .B(
        \pool/pool/pe_b/peij_0_1/add/fai_10/n3 ), .Z(
        \pool/pool/pe_b/peij_0_1/d_acc [10]) );
  INV_X2 \pool/pool/pe_b/peij_0_1/add/fai_10/U2  ( .A(
        \pool/pool/pe_b/peij_0_1/add/fai_10/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_1/add/c_out ) );
  AOI22_X2 \pool/pool/pe_b/peij_0_1/add/fai_10/U1  ( .A1(
        \pool/pool/pe_b/peij_0_1/add/notb [10]), .A2(
        \pool/pool/pe_b_o_data[0][32] ), .B1(
        \pool/pool/pe_b/peij_0_1/add/fai_10/n3 ), .B2(
        \pool/pool/pe_b/peij_0_1/add/cprop [10]), .ZN(
        \pool/pool/pe_b/peij_0_1/add/fai_10/n1 ) );
  INV_X1 \pool/pool/pe_b/peij_0_2/U22  ( .A(\pool/pool/pe_b/n6 ), .ZN(
        \pool/pool/pe_b/peij_0_2/n16 ) );
  INV_X1 \pool/pool/pe_b/peij_0_2/U14  ( .A(\pool/pool/pe_b/n6 ), .ZN(
        \pool/pool/pe_b/peij_0_2/n12 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_2/U13  ( .A1(
        \pool/pool/pe_b/peij_0_2/d_acc [0]), .A2(\pool/pool/pe_b/peij_0_2/n18 ), .ZN(\pool/pool/pe_b/peij_0_2/n11 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_2/U12  ( .A1(
        \pool/pool/pe_b/peij_0_2/d_acc [1]), .A2(\pool/pool/pe_b/peij_0_2/n18 ), .ZN(\pool/pool/pe_b/peij_0_2/n10 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_2/U11  ( .A1(
        \pool/pool/pe_b/peij_0_2/d_acc [2]), .A2(\pool/pool/pe_b/peij_0_2/n18 ), .ZN(\pool/pool/pe_b/peij_0_2/n9 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_2/U10  ( .A1(
        \pool/pool/pe_b/peij_0_2/d_acc [3]), .A2(\pool/pool/pe_b/peij_0_2/n18 ), .ZN(\pool/pool/pe_b/peij_0_2/n8 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_2/U9  ( .A1(
        \pool/pool/pe_b/peij_0_2/d_acc [4]), .A2(\pool/pool/pe_b/peij_0_2/n18 ), .ZN(\pool/pool/pe_b/peij_0_2/n7 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_2/U8  ( .A1(
        \pool/pool/pe_b/peij_0_2/d_acc [5]), .A2(\pool/pool/pe_b/peij_0_2/n18 ), .ZN(\pool/pool/pe_b/peij_0_2/n6 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_2/U7  ( .A1(
        \pool/pool/pe_b/peij_0_2/d_acc [6]), .A2(\pool/pool/pe_b/peij_0_2/n18 ), .ZN(\pool/pool/pe_b/peij_0_2/n5 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_2/U6  ( .A1(
        \pool/pool/pe_b/peij_0_2/d_acc [7]), .A2(\pool/pool/pe_b/peij_0_2/n18 ), .ZN(\pool/pool/pe_b/peij_0_2/n4 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_2/U5  ( .A1(
        \pool/pool/pe_b/peij_0_2/d_acc [8]), .A2(\pool/pool/pe_b/peij_0_2/n18 ), .ZN(\pool/pool/pe_b/peij_0_2/n3 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_2/U4  ( .A1(
        \pool/pool/pe_b/peij_0_2/d_acc [9]), .A2(\pool/pool/pe_b/peij_0_2/n18 ), .ZN(\pool/pool/pe_b/peij_0_2/n2 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_2/U3  ( .A1(
        \pool/pool/pe_b/peij_0_2/d_acc [10]), .A2(
        \pool/pool/pe_b/peij_0_2/n18 ), .ZN(\pool/pool/pe_b/peij_0_2/n1 ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_2/q_acc_reg[10]  ( .D(
        \pool/pool/pe_b/peij_0_2/n1 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_2/n16 ), .Q(\pool/pool/pe_b_o_data[0][21] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_2/q_acc_reg[9]  ( .D(
        \pool/pool/pe_b/peij_0_2/n2 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_2/n16 ), .Q(\pool/pool/pe_b_o_data[0][20] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_2/q_acc_reg[8]  ( .D(
        \pool/pool/pe_b/peij_0_2/n3 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_2/n16 ), .Q(\pool/pool/pe_b_o_data[0][19] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_2/q_acc_reg[7]  ( .D(
        \pool/pool/pe_b/peij_0_2/n4 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_2/n16 ), .Q(\pool/pool/pe_b_o_data[0][18] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_2/q_acc_reg[6]  ( .D(
        \pool/pool/pe_b/peij_0_2/n5 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_2/n16 ), .Q(\pool/pool/pe_b_o_data[0][17] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_2/q_acc_reg[5]  ( .D(
        \pool/pool/pe_b/peij_0_2/n6 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_2/n16 ), .Q(\pool/pool/pe_b_o_data[0][16] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_2/q_acc_reg[4]  ( .D(
        \pool/pool/pe_b/peij_0_2/n7 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_2/n16 ), .Q(\pool/pool/pe_b_o_data[0][15] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_2/q_acc_reg[3]  ( .D(
        \pool/pool/pe_b/peij_0_2/n8 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_2/n16 ), .Q(\pool/pool/pe_b_o_data[0][14] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_2/q_acc_reg[2]  ( .D(
        \pool/pool/pe_b/peij_0_2/n9 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_2/n16 ), .Q(\pool/pool/pe_b_o_data[0][13] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_2/q_acc_reg[1]  ( .D(
        \pool/pool/pe_b/peij_0_2/n10 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_2/n16 ), .Q(\pool/pool/pe_b_o_data[0][12] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_2/q_acc_reg[0]  ( .D(
        \pool/pool/pe_b/peij_0_2/n11 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_2/n16 ), .Q(\pool/pool/pe_b_o_data[0][11] ) );
  INV_X2 \pool/pool/pe_b/peij_0_2/U21  ( .A(\pool/sync_clr ), .ZN(
        \pool/pool/pe_b/peij_0_2/n18 ) );
  AND3_X2 \pool/pool/pe_b/peij_0_2/U20  ( .A1(\pool/pool/pe_b/int_pe_en[0][2] ), .A2(\pool/pool/pe_b/peij_0_2/n18 ), .A3(1'b1), .ZN(
        \pool/pool/pe_b/peij_0_2/n17 ) );
  AND2_X2 \pool/pool/pe_b/peij_0_2/U19  ( .A1(\pool/pool/pe_b_i_data[0][4] ), 
        .A2(\pool/pool/pe_b/peij_0_2/n17 ), .ZN(\pool/pool/pe_b/peij_0_2/N33 )
         );
  AND2_X2 \pool/pool/pe_b/peij_0_2/U18  ( .A1(\pool/pool/pe_b_i_data[0][5] ), 
        .A2(\pool/pool/pe_b/peij_0_2/n17 ), .ZN(\pool/pool/pe_b/peij_0_2/N34 )
         );
  AND2_X2 \pool/pool/pe_b/peij_0_2/U17  ( .A1(\pool/pool/pe_b_i_data[0][6] ), 
        .A2(\pool/pool/pe_b/peij_0_2/n17 ), .ZN(\pool/pool/pe_b/peij_0_2/N35 )
         );
  AND4_X4 \pool/pool/pe_b/peij_0_2/U16  ( .A1(1'b1), .A2(
        \pool/pool/pe_b_i_data[0][7] ), .A3(\pool/pool/pe_b/int_pe_en[0][2] ), 
        .A4(\pool/pool/pe_b/peij_0_2/n18 ), .ZN(\pool/pool/pe_b/peij_0_2/N36 )
         );
  DFFR_X1 \pool/pool/pe_b/peij_0_2/q_im_reg[0]  ( .D(
        \pool/pool/pe_b/peij_0_2/N33 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_2/n12 ), .Q(\pool/pool/pe_b/peij_0_2/sgnext [0]) );
  DFFR_X1 \pool/pool/pe_b/peij_0_2/q_im_reg[1]  ( .D(
        \pool/pool/pe_b/peij_0_2/N34 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_2/n12 ), .Q(\pool/pool/pe_b/peij_0_2/sgnext [1]) );
  DFFR_X1 \pool/pool/pe_b/peij_0_2/q_im_reg[2]  ( .D(
        \pool/pool/pe_b/peij_0_2/N35 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_2/n12 ), .Q(\pool/pool/pe_b/peij_0_2/sgnext [2]) );
  DFFR_X1 \pool/pool/pe_b/peij_0_2/q_im_reg[3]  ( .D(
        \pool/pool/pe_b/peij_0_2/N36 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_2/n12 ), .Q(\pool/pool/pe_b/peij_0_2/sgnext_10 ) );
  SDFFR_X1 \pool/pool/pe_b/peij_0_2/q_k_reg  ( .D(1'b0), .SI(
        \pool/pool/pe_b/peij_0_2/n18 ), .SE(1'b0), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_2/n12 ), .Q(\pool/pool/pe_b/peij_0_2/q_k ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/U11  ( .A(
        \pool/pool/pe_b/peij_0_2/sgnext [0]), .B(\pool/pool/pe_b/peij_0_2/q_k ), .Z(\pool/pool/pe_b/peij_0_2/add/notb [0]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/U10  ( .A(
        \pool/pool/pe_b/peij_0_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_2/q_k ), .Z(\pool/pool/pe_b/peij_0_2/add/notb [10]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/U9  ( .A(
        \pool/pool/pe_b/peij_0_2/sgnext [1]), .B(\pool/pool/pe_b/peij_0_2/q_k ), .Z(\pool/pool/pe_b/peij_0_2/add/notb [1]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/U8  ( .A(
        \pool/pool/pe_b/peij_0_2/sgnext [2]), .B(\pool/pool/pe_b/peij_0_2/q_k ), .Z(\pool/pool/pe_b/peij_0_2/add/notb [2]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/U7  ( .A(
        \pool/pool/pe_b/peij_0_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_2/q_k ), .Z(\pool/pool/pe_b/peij_0_2/add/notb [3]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/U6  ( .A(
        \pool/pool/pe_b/peij_0_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_2/q_k ), .Z(\pool/pool/pe_b/peij_0_2/add/notb [4]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/U5  ( .A(
        \pool/pool/pe_b/peij_0_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_2/q_k ), .Z(\pool/pool/pe_b/peij_0_2/add/notb [5]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/U4  ( .A(
        \pool/pool/pe_b/peij_0_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_2/q_k ), .Z(\pool/pool/pe_b/peij_0_2/add/notb [6]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/U3  ( .A(
        \pool/pool/pe_b/peij_0_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_2/q_k ), .Z(\pool/pool/pe_b/peij_0_2/add/notb [7]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/U2  ( .A(
        \pool/pool/pe_b/peij_0_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_2/q_k ), .Z(\pool/pool/pe_b/peij_0_2/add/notb [8]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/U1  ( .A(
        \pool/pool/pe_b/peij_0_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_2/q_k ), .Z(\pool/pool/pe_b/peij_0_2/add/notb [9]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_0/U4  ( .A(
        \pool/pool/pe_b_o_data[0][11] ), .B(
        \pool/pool/pe_b/peij_0_2/add/notb [0]), .Z(
        \pool/pool/pe_b/peij_0_2/add/fai_0/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_0/U3  ( .A(
        \pool/pool/pe_b/peij_0_2/q_k ), .B(
        \pool/pool/pe_b/peij_0_2/add/fai_0/n3 ), .Z(
        \pool/pool/pe_b/peij_0_2/d_acc [0]) );
  INV_X2 \pool/pool/pe_b/peij_0_2/add/fai_0/U2  ( .A(
        \pool/pool/pe_b/peij_0_2/add/fai_0/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_2/add/cprop [1]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_2/add/fai_0/U1  ( .A1(
        \pool/pool/pe_b/peij_0_2/add/notb [0]), .A2(
        \pool/pool/pe_b_o_data[0][11] ), .B1(
        \pool/pool/pe_b/peij_0_2/add/fai_0/n3 ), .B2(
        \pool/pool/pe_b/peij_0_2/q_k ), .ZN(
        \pool/pool/pe_b/peij_0_2/add/fai_0/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_1/U4  ( .A(
        \pool/pool/pe_b_o_data[0][12] ), .B(
        \pool/pool/pe_b/peij_0_2/add/notb [1]), .Z(
        \pool/pool/pe_b/peij_0_2/add/fai_1/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_1/U3  ( .A(
        \pool/pool/pe_b/peij_0_2/add/cprop [1]), .B(
        \pool/pool/pe_b/peij_0_2/add/fai_1/n3 ), .Z(
        \pool/pool/pe_b/peij_0_2/d_acc [1]) );
  INV_X2 \pool/pool/pe_b/peij_0_2/add/fai_1/U2  ( .A(
        \pool/pool/pe_b/peij_0_2/add/fai_1/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_2/add/cprop [2]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_2/add/fai_1/U1  ( .A1(
        \pool/pool/pe_b/peij_0_2/add/notb [1]), .A2(
        \pool/pool/pe_b_o_data[0][12] ), .B1(
        \pool/pool/pe_b/peij_0_2/add/fai_1/n3 ), .B2(
        \pool/pool/pe_b/peij_0_2/add/cprop [1]), .ZN(
        \pool/pool/pe_b/peij_0_2/add/fai_1/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_2/U4  ( .A(
        \pool/pool/pe_b_o_data[0][13] ), .B(
        \pool/pool/pe_b/peij_0_2/add/notb [2]), .Z(
        \pool/pool/pe_b/peij_0_2/add/fai_2/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_2/U3  ( .A(
        \pool/pool/pe_b/peij_0_2/add/cprop [2]), .B(
        \pool/pool/pe_b/peij_0_2/add/fai_2/n3 ), .Z(
        \pool/pool/pe_b/peij_0_2/d_acc [2]) );
  INV_X2 \pool/pool/pe_b/peij_0_2/add/fai_2/U2  ( .A(
        \pool/pool/pe_b/peij_0_2/add/fai_2/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_2/add/cprop [3]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_2/add/fai_2/U1  ( .A1(
        \pool/pool/pe_b/peij_0_2/add/notb [2]), .A2(
        \pool/pool/pe_b_o_data[0][13] ), .B1(
        \pool/pool/pe_b/peij_0_2/add/fai_2/n3 ), .B2(
        \pool/pool/pe_b/peij_0_2/add/cprop [2]), .ZN(
        \pool/pool/pe_b/peij_0_2/add/fai_2/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_3/U4  ( .A(
        \pool/pool/pe_b_o_data[0][14] ), .B(
        \pool/pool/pe_b/peij_0_2/add/notb [3]), .Z(
        \pool/pool/pe_b/peij_0_2/add/fai_3/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_3/U3  ( .A(
        \pool/pool/pe_b/peij_0_2/add/cprop [3]), .B(
        \pool/pool/pe_b/peij_0_2/add/fai_3/n3 ), .Z(
        \pool/pool/pe_b/peij_0_2/d_acc [3]) );
  INV_X2 \pool/pool/pe_b/peij_0_2/add/fai_3/U2  ( .A(
        \pool/pool/pe_b/peij_0_2/add/fai_3/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_2/add/cprop [4]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_2/add/fai_3/U1  ( .A1(
        \pool/pool/pe_b/peij_0_2/add/notb [3]), .A2(
        \pool/pool/pe_b_o_data[0][14] ), .B1(
        \pool/pool/pe_b/peij_0_2/add/fai_3/n3 ), .B2(
        \pool/pool/pe_b/peij_0_2/add/cprop [3]), .ZN(
        \pool/pool/pe_b/peij_0_2/add/fai_3/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_4/U4  ( .A(
        \pool/pool/pe_b_o_data[0][15] ), .B(
        \pool/pool/pe_b/peij_0_2/add/notb [4]), .Z(
        \pool/pool/pe_b/peij_0_2/add/fai_4/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_4/U3  ( .A(
        \pool/pool/pe_b/peij_0_2/add/cprop [4]), .B(
        \pool/pool/pe_b/peij_0_2/add/fai_4/n3 ), .Z(
        \pool/pool/pe_b/peij_0_2/d_acc [4]) );
  INV_X2 \pool/pool/pe_b/peij_0_2/add/fai_4/U2  ( .A(
        \pool/pool/pe_b/peij_0_2/add/fai_4/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_2/add/cprop [5]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_2/add/fai_4/U1  ( .A1(
        \pool/pool/pe_b/peij_0_2/add/notb [4]), .A2(
        \pool/pool/pe_b_o_data[0][15] ), .B1(
        \pool/pool/pe_b/peij_0_2/add/fai_4/n3 ), .B2(
        \pool/pool/pe_b/peij_0_2/add/cprop [4]), .ZN(
        \pool/pool/pe_b/peij_0_2/add/fai_4/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_5/U4  ( .A(
        \pool/pool/pe_b_o_data[0][16] ), .B(
        \pool/pool/pe_b/peij_0_2/add/notb [5]), .Z(
        \pool/pool/pe_b/peij_0_2/add/fai_5/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_5/U3  ( .A(
        \pool/pool/pe_b/peij_0_2/add/cprop [5]), .B(
        \pool/pool/pe_b/peij_0_2/add/fai_5/n3 ), .Z(
        \pool/pool/pe_b/peij_0_2/d_acc [5]) );
  INV_X2 \pool/pool/pe_b/peij_0_2/add/fai_5/U2  ( .A(
        \pool/pool/pe_b/peij_0_2/add/fai_5/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_2/add/cprop [6]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_2/add/fai_5/U1  ( .A1(
        \pool/pool/pe_b/peij_0_2/add/notb [5]), .A2(
        \pool/pool/pe_b_o_data[0][16] ), .B1(
        \pool/pool/pe_b/peij_0_2/add/fai_5/n3 ), .B2(
        \pool/pool/pe_b/peij_0_2/add/cprop [5]), .ZN(
        \pool/pool/pe_b/peij_0_2/add/fai_5/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_6/U4  ( .A(
        \pool/pool/pe_b_o_data[0][17] ), .B(
        \pool/pool/pe_b/peij_0_2/add/notb [6]), .Z(
        \pool/pool/pe_b/peij_0_2/add/fai_6/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_6/U3  ( .A(
        \pool/pool/pe_b/peij_0_2/add/cprop [6]), .B(
        \pool/pool/pe_b/peij_0_2/add/fai_6/n3 ), .Z(
        \pool/pool/pe_b/peij_0_2/d_acc [6]) );
  INV_X2 \pool/pool/pe_b/peij_0_2/add/fai_6/U2  ( .A(
        \pool/pool/pe_b/peij_0_2/add/fai_6/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_2/add/cprop [7]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_2/add/fai_6/U1  ( .A1(
        \pool/pool/pe_b/peij_0_2/add/notb [6]), .A2(
        \pool/pool/pe_b_o_data[0][17] ), .B1(
        \pool/pool/pe_b/peij_0_2/add/fai_6/n3 ), .B2(
        \pool/pool/pe_b/peij_0_2/add/cprop [6]), .ZN(
        \pool/pool/pe_b/peij_0_2/add/fai_6/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_7/U4  ( .A(
        \pool/pool/pe_b_o_data[0][18] ), .B(
        \pool/pool/pe_b/peij_0_2/add/notb [7]), .Z(
        \pool/pool/pe_b/peij_0_2/add/fai_7/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_7/U3  ( .A(
        \pool/pool/pe_b/peij_0_2/add/cprop [7]), .B(
        \pool/pool/pe_b/peij_0_2/add/fai_7/n3 ), .Z(
        \pool/pool/pe_b/peij_0_2/d_acc [7]) );
  INV_X2 \pool/pool/pe_b/peij_0_2/add/fai_7/U2  ( .A(
        \pool/pool/pe_b/peij_0_2/add/fai_7/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_2/add/cprop [8]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_2/add/fai_7/U1  ( .A1(
        \pool/pool/pe_b/peij_0_2/add/notb [7]), .A2(
        \pool/pool/pe_b_o_data[0][18] ), .B1(
        \pool/pool/pe_b/peij_0_2/add/fai_7/n3 ), .B2(
        \pool/pool/pe_b/peij_0_2/add/cprop [7]), .ZN(
        \pool/pool/pe_b/peij_0_2/add/fai_7/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_8/U4  ( .A(
        \pool/pool/pe_b_o_data[0][19] ), .B(
        \pool/pool/pe_b/peij_0_2/add/notb [8]), .Z(
        \pool/pool/pe_b/peij_0_2/add/fai_8/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_8/U3  ( .A(
        \pool/pool/pe_b/peij_0_2/add/cprop [8]), .B(
        \pool/pool/pe_b/peij_0_2/add/fai_8/n3 ), .Z(
        \pool/pool/pe_b/peij_0_2/d_acc [8]) );
  INV_X2 \pool/pool/pe_b/peij_0_2/add/fai_8/U2  ( .A(
        \pool/pool/pe_b/peij_0_2/add/fai_8/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_2/add/cprop [9]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_2/add/fai_8/U1  ( .A1(
        \pool/pool/pe_b/peij_0_2/add/notb [8]), .A2(
        \pool/pool/pe_b_o_data[0][19] ), .B1(
        \pool/pool/pe_b/peij_0_2/add/fai_8/n3 ), .B2(
        \pool/pool/pe_b/peij_0_2/add/cprop [8]), .ZN(
        \pool/pool/pe_b/peij_0_2/add/fai_8/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_9/U4  ( .A(
        \pool/pool/pe_b_o_data[0][20] ), .B(
        \pool/pool/pe_b/peij_0_2/add/notb [9]), .Z(
        \pool/pool/pe_b/peij_0_2/add/fai_9/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_9/U3  ( .A(
        \pool/pool/pe_b/peij_0_2/add/cprop [9]), .B(
        \pool/pool/pe_b/peij_0_2/add/fai_9/n3 ), .Z(
        \pool/pool/pe_b/peij_0_2/d_acc [9]) );
  INV_X2 \pool/pool/pe_b/peij_0_2/add/fai_9/U2  ( .A(
        \pool/pool/pe_b/peij_0_2/add/fai_9/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_2/add/cprop [10]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_2/add/fai_9/U1  ( .A1(
        \pool/pool/pe_b/peij_0_2/add/notb [9]), .A2(
        \pool/pool/pe_b_o_data[0][20] ), .B1(
        \pool/pool/pe_b/peij_0_2/add/fai_9/n3 ), .B2(
        \pool/pool/pe_b/peij_0_2/add/cprop [9]), .ZN(
        \pool/pool/pe_b/peij_0_2/add/fai_9/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_10/U4  ( .A(
        \pool/pool/pe_b_o_data[0][21] ), .B(
        \pool/pool/pe_b/peij_0_2/add/notb [10]), .Z(
        \pool/pool/pe_b/peij_0_2/add/fai_10/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_2/add/fai_10/U3  ( .A(
        \pool/pool/pe_b/peij_0_2/add/cprop [10]), .B(
        \pool/pool/pe_b/peij_0_2/add/fai_10/n3 ), .Z(
        \pool/pool/pe_b/peij_0_2/d_acc [10]) );
  INV_X2 \pool/pool/pe_b/peij_0_2/add/fai_10/U2  ( .A(
        \pool/pool/pe_b/peij_0_2/add/fai_10/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_2/add/c_out ) );
  AOI22_X2 \pool/pool/pe_b/peij_0_2/add/fai_10/U1  ( .A1(
        \pool/pool/pe_b/peij_0_2/add/notb [10]), .A2(
        \pool/pool/pe_b_o_data[0][21] ), .B1(
        \pool/pool/pe_b/peij_0_2/add/fai_10/n3 ), .B2(
        \pool/pool/pe_b/peij_0_2/add/cprop [10]), .ZN(
        \pool/pool/pe_b/peij_0_2/add/fai_10/n1 ) );
  INV_X1 \pool/pool/pe_b/peij_0_3/U22  ( .A(\pool/pool/pe_b/n6 ), .ZN(
        \pool/pool/pe_b/peij_0_3/n16 ) );
  INV_X1 \pool/pool/pe_b/peij_0_3/U14  ( .A(\pool/pool/pe_b/n6 ), .ZN(
        \pool/pool/pe_b/peij_0_3/n12 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_3/U13  ( .A1(
        \pool/pool/pe_b/peij_0_3/d_acc [0]), .A2(\pool/pool/pe_b/peij_0_3/n18 ), .ZN(\pool/pool/pe_b/peij_0_3/n11 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_3/U12  ( .A1(
        \pool/pool/pe_b/peij_0_3/d_acc [1]), .A2(\pool/pool/pe_b/peij_0_3/n18 ), .ZN(\pool/pool/pe_b/peij_0_3/n10 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_3/U11  ( .A1(
        \pool/pool/pe_b/peij_0_3/d_acc [2]), .A2(\pool/pool/pe_b/peij_0_3/n18 ), .ZN(\pool/pool/pe_b/peij_0_3/n9 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_3/U10  ( .A1(
        \pool/pool/pe_b/peij_0_3/d_acc [3]), .A2(\pool/pool/pe_b/peij_0_3/n18 ), .ZN(\pool/pool/pe_b/peij_0_3/n8 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_3/U9  ( .A1(
        \pool/pool/pe_b/peij_0_3/d_acc [4]), .A2(\pool/pool/pe_b/peij_0_3/n18 ), .ZN(\pool/pool/pe_b/peij_0_3/n7 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_3/U8  ( .A1(
        \pool/pool/pe_b/peij_0_3/d_acc [5]), .A2(\pool/pool/pe_b/peij_0_3/n18 ), .ZN(\pool/pool/pe_b/peij_0_3/n6 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_3/U7  ( .A1(
        \pool/pool/pe_b/peij_0_3/d_acc [6]), .A2(\pool/pool/pe_b/peij_0_3/n18 ), .ZN(\pool/pool/pe_b/peij_0_3/n5 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_3/U6  ( .A1(
        \pool/pool/pe_b/peij_0_3/d_acc [7]), .A2(\pool/pool/pe_b/peij_0_3/n18 ), .ZN(\pool/pool/pe_b/peij_0_3/n4 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_3/U5  ( .A1(
        \pool/pool/pe_b/peij_0_3/d_acc [8]), .A2(\pool/pool/pe_b/peij_0_3/n18 ), .ZN(\pool/pool/pe_b/peij_0_3/n3 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_3/U4  ( .A1(
        \pool/pool/pe_b/peij_0_3/d_acc [9]), .A2(\pool/pool/pe_b/peij_0_3/n18 ), .ZN(\pool/pool/pe_b/peij_0_3/n2 ) );
  AND2_X1 \pool/pool/pe_b/peij_0_3/U3  ( .A1(
        \pool/pool/pe_b/peij_0_3/d_acc [10]), .A2(
        \pool/pool/pe_b/peij_0_3/n18 ), .ZN(\pool/pool/pe_b/peij_0_3/n1 ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_3/q_acc_reg[10]  ( .D(
        \pool/pool/pe_b/peij_0_3/n1 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_3/n16 ), .Q(\pool/pool/pe_b_o_data[0][10] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_3/q_acc_reg[9]  ( .D(
        \pool/pool/pe_b/peij_0_3/n2 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_3/n16 ), .Q(\pool/pool/pe_b_o_data[0][9] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_3/q_acc_reg[8]  ( .D(
        \pool/pool/pe_b/peij_0_3/n3 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_3/n16 ), .Q(\pool/pool/pe_b_o_data[0][8] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_3/q_acc_reg[7]  ( .D(
        \pool/pool/pe_b/peij_0_3/n4 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_3/n16 ), .Q(\pool/pool/pe_b_o_data[0][7] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_3/q_acc_reg[6]  ( .D(
        \pool/pool/pe_b/peij_0_3/n5 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_3/n16 ), .Q(\pool/pool/pe_b_o_data[0][6] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_3/q_acc_reg[5]  ( .D(
        \pool/pool/pe_b/peij_0_3/n6 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_3/n16 ), .Q(\pool/pool/pe_b_o_data[0][5] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_3/q_acc_reg[4]  ( .D(
        \pool/pool/pe_b/peij_0_3/n7 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_3/n16 ), .Q(\pool/pool/pe_b_o_data[0][4] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_3/q_acc_reg[3]  ( .D(
        \pool/pool/pe_b/peij_0_3/n8 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_3/n16 ), .Q(\pool/pool/pe_b_o_data[0][3] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_3/q_acc_reg[2]  ( .D(
        \pool/pool/pe_b/peij_0_3/n9 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_3/n16 ), .Q(\pool/pool/pe_b_o_data[0][2] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_3/q_acc_reg[1]  ( .D(
        \pool/pool/pe_b/peij_0_3/n10 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_3/n16 ), .Q(\pool/pool/pe_b_o_data[0][1] ) );
  DFFR_X1 \pool/pool/pe_b/peij_0_3/q_acc_reg[0]  ( .D(
        \pool/pool/pe_b/peij_0_3/n11 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_3/n16 ), .Q(\pool/pool/pe_b_o_data[0][0] ) );
  INV_X2 \pool/pool/pe_b/peij_0_3/U21  ( .A(\pool/sync_clr ), .ZN(
        \pool/pool/pe_b/peij_0_3/n18 ) );
  AND3_X2 \pool/pool/pe_b/peij_0_3/U20  ( .A1(\pool/pool/pe_b/int_pe_en[0][3] ), .A2(\pool/pool/pe_b/peij_0_3/n18 ), .A3(1'b1), .ZN(
        \pool/pool/pe_b/peij_0_3/n17 ) );
  AND2_X2 \pool/pool/pe_b/peij_0_3/U19  ( .A1(\pool/pool/pe_b_i_data[0][0] ), 
        .A2(\pool/pool/pe_b/peij_0_3/n17 ), .ZN(\pool/pool/pe_b/peij_0_3/N33 )
         );
  AND2_X2 \pool/pool/pe_b/peij_0_3/U18  ( .A1(\pool/pool/pe_b_i_data[0][1] ), 
        .A2(\pool/pool/pe_b/peij_0_3/n17 ), .ZN(\pool/pool/pe_b/peij_0_3/N34 )
         );
  AND2_X2 \pool/pool/pe_b/peij_0_3/U17  ( .A1(\pool/pool/pe_b_i_data[0][2] ), 
        .A2(\pool/pool/pe_b/peij_0_3/n17 ), .ZN(\pool/pool/pe_b/peij_0_3/N35 )
         );
  AND4_X4 \pool/pool/pe_b/peij_0_3/U16  ( .A1(1'b1), .A2(
        \pool/pool/pe_b_i_data[0][3] ), .A3(\pool/pool/pe_b/int_pe_en[0][3] ), 
        .A4(\pool/pool/pe_b/peij_0_3/n18 ), .ZN(\pool/pool/pe_b/peij_0_3/N36 )
         );
  DFFR_X1 \pool/pool/pe_b/peij_0_3/q_im_reg[0]  ( .D(
        \pool/pool/pe_b/peij_0_3/N33 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_3/n12 ), .Q(\pool/pool/pe_b/peij_0_3/sgnext [0]) );
  DFFR_X1 \pool/pool/pe_b/peij_0_3/q_im_reg[1]  ( .D(
        \pool/pool/pe_b/peij_0_3/N34 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_3/n12 ), .Q(\pool/pool/pe_b/peij_0_3/sgnext [1]) );
  DFFR_X1 \pool/pool/pe_b/peij_0_3/q_im_reg[2]  ( .D(
        \pool/pool/pe_b/peij_0_3/N35 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_3/n12 ), .Q(\pool/pool/pe_b/peij_0_3/sgnext [2]) );
  DFFR_X1 \pool/pool/pe_b/peij_0_3/q_im_reg[3]  ( .D(
        \pool/pool/pe_b/peij_0_3/N36 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_3/n12 ), .Q(\pool/pool/pe_b/peij_0_3/sgnext_10 ) );
  SDFFR_X1 \pool/pool/pe_b/peij_0_3/q_k_reg  ( .D(1'b0), .SI(
        \pool/pool/pe_b/peij_0_3/n18 ), .SE(1'b0), .CK(clk), .RN(
        \pool/pool/pe_b/peij_0_3/n12 ), .Q(\pool/pool/pe_b/peij_0_3/q_k ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/U11  ( .A(
        \pool/pool/pe_b/peij_0_3/sgnext [0]), .B(\pool/pool/pe_b/peij_0_3/q_k ), .Z(\pool/pool/pe_b/peij_0_3/add/notb [0]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/U10  ( .A(
        \pool/pool/pe_b/peij_0_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_3/q_k ), .Z(\pool/pool/pe_b/peij_0_3/add/notb [10]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/U9  ( .A(
        \pool/pool/pe_b/peij_0_3/sgnext [1]), .B(\pool/pool/pe_b/peij_0_3/q_k ), .Z(\pool/pool/pe_b/peij_0_3/add/notb [1]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/U8  ( .A(
        \pool/pool/pe_b/peij_0_3/sgnext [2]), .B(\pool/pool/pe_b/peij_0_3/q_k ), .Z(\pool/pool/pe_b/peij_0_3/add/notb [2]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/U7  ( .A(
        \pool/pool/pe_b/peij_0_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_3/q_k ), .Z(\pool/pool/pe_b/peij_0_3/add/notb [3]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/U6  ( .A(
        \pool/pool/pe_b/peij_0_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_3/q_k ), .Z(\pool/pool/pe_b/peij_0_3/add/notb [4]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/U5  ( .A(
        \pool/pool/pe_b/peij_0_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_3/q_k ), .Z(\pool/pool/pe_b/peij_0_3/add/notb [5]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/U4  ( .A(
        \pool/pool/pe_b/peij_0_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_3/q_k ), .Z(\pool/pool/pe_b/peij_0_3/add/notb [6]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/U3  ( .A(
        \pool/pool/pe_b/peij_0_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_3/q_k ), .Z(\pool/pool/pe_b/peij_0_3/add/notb [7]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/U2  ( .A(
        \pool/pool/pe_b/peij_0_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_3/q_k ), .Z(\pool/pool/pe_b/peij_0_3/add/notb [8]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/U1  ( .A(
        \pool/pool/pe_b/peij_0_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_0_3/q_k ), .Z(\pool/pool/pe_b/peij_0_3/add/notb [9]) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_0/U4  ( .A(
        \pool/pool/pe_b_o_data[0][0] ), .B(
        \pool/pool/pe_b/peij_0_3/add/notb [0]), .Z(
        \pool/pool/pe_b/peij_0_3/add/fai_0/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_0/U3  ( .A(
        \pool/pool/pe_b/peij_0_3/q_k ), .B(
        \pool/pool/pe_b/peij_0_3/add/fai_0/n3 ), .Z(
        \pool/pool/pe_b/peij_0_3/d_acc [0]) );
  INV_X2 \pool/pool/pe_b/peij_0_3/add/fai_0/U2  ( .A(
        \pool/pool/pe_b/peij_0_3/add/fai_0/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_3/add/cprop [1]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_3/add/fai_0/U1  ( .A1(
        \pool/pool/pe_b/peij_0_3/add/notb [0]), .A2(
        \pool/pool/pe_b_o_data[0][0] ), .B1(
        \pool/pool/pe_b/peij_0_3/add/fai_0/n3 ), .B2(
        \pool/pool/pe_b/peij_0_3/q_k ), .ZN(
        \pool/pool/pe_b/peij_0_3/add/fai_0/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_1/U4  ( .A(
        \pool/pool/pe_b_o_data[0][1] ), .B(
        \pool/pool/pe_b/peij_0_3/add/notb [1]), .Z(
        \pool/pool/pe_b/peij_0_3/add/fai_1/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_1/U3  ( .A(
        \pool/pool/pe_b/peij_0_3/add/cprop [1]), .B(
        \pool/pool/pe_b/peij_0_3/add/fai_1/n3 ), .Z(
        \pool/pool/pe_b/peij_0_3/d_acc [1]) );
  INV_X2 \pool/pool/pe_b/peij_0_3/add/fai_1/U2  ( .A(
        \pool/pool/pe_b/peij_0_3/add/fai_1/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_3/add/cprop [2]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_3/add/fai_1/U1  ( .A1(
        \pool/pool/pe_b/peij_0_3/add/notb [1]), .A2(
        \pool/pool/pe_b_o_data[0][1] ), .B1(
        \pool/pool/pe_b/peij_0_3/add/fai_1/n3 ), .B2(
        \pool/pool/pe_b/peij_0_3/add/cprop [1]), .ZN(
        \pool/pool/pe_b/peij_0_3/add/fai_1/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_2/U4  ( .A(
        \pool/pool/pe_b_o_data[0][2] ), .B(
        \pool/pool/pe_b/peij_0_3/add/notb [2]), .Z(
        \pool/pool/pe_b/peij_0_3/add/fai_2/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_2/U3  ( .A(
        \pool/pool/pe_b/peij_0_3/add/cprop [2]), .B(
        \pool/pool/pe_b/peij_0_3/add/fai_2/n3 ), .Z(
        \pool/pool/pe_b/peij_0_3/d_acc [2]) );
  INV_X2 \pool/pool/pe_b/peij_0_3/add/fai_2/U2  ( .A(
        \pool/pool/pe_b/peij_0_3/add/fai_2/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_3/add/cprop [3]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_3/add/fai_2/U1  ( .A1(
        \pool/pool/pe_b/peij_0_3/add/notb [2]), .A2(
        \pool/pool/pe_b_o_data[0][2] ), .B1(
        \pool/pool/pe_b/peij_0_3/add/fai_2/n3 ), .B2(
        \pool/pool/pe_b/peij_0_3/add/cprop [2]), .ZN(
        \pool/pool/pe_b/peij_0_3/add/fai_2/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_3/U4  ( .A(
        \pool/pool/pe_b_o_data[0][3] ), .B(
        \pool/pool/pe_b/peij_0_3/add/notb [3]), .Z(
        \pool/pool/pe_b/peij_0_3/add/fai_3/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_3/U3  ( .A(
        \pool/pool/pe_b/peij_0_3/add/cprop [3]), .B(
        \pool/pool/pe_b/peij_0_3/add/fai_3/n3 ), .Z(
        \pool/pool/pe_b/peij_0_3/d_acc [3]) );
  INV_X2 \pool/pool/pe_b/peij_0_3/add/fai_3/U2  ( .A(
        \pool/pool/pe_b/peij_0_3/add/fai_3/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_3/add/cprop [4]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_3/add/fai_3/U1  ( .A1(
        \pool/pool/pe_b/peij_0_3/add/notb [3]), .A2(
        \pool/pool/pe_b_o_data[0][3] ), .B1(
        \pool/pool/pe_b/peij_0_3/add/fai_3/n3 ), .B2(
        \pool/pool/pe_b/peij_0_3/add/cprop [3]), .ZN(
        \pool/pool/pe_b/peij_0_3/add/fai_3/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_4/U4  ( .A(
        \pool/pool/pe_b_o_data[0][4] ), .B(
        \pool/pool/pe_b/peij_0_3/add/notb [4]), .Z(
        \pool/pool/pe_b/peij_0_3/add/fai_4/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_4/U3  ( .A(
        \pool/pool/pe_b/peij_0_3/add/cprop [4]), .B(
        \pool/pool/pe_b/peij_0_3/add/fai_4/n3 ), .Z(
        \pool/pool/pe_b/peij_0_3/d_acc [4]) );
  INV_X2 \pool/pool/pe_b/peij_0_3/add/fai_4/U2  ( .A(
        \pool/pool/pe_b/peij_0_3/add/fai_4/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_3/add/cprop [5]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_3/add/fai_4/U1  ( .A1(
        \pool/pool/pe_b/peij_0_3/add/notb [4]), .A2(
        \pool/pool/pe_b_o_data[0][4] ), .B1(
        \pool/pool/pe_b/peij_0_3/add/fai_4/n3 ), .B2(
        \pool/pool/pe_b/peij_0_3/add/cprop [4]), .ZN(
        \pool/pool/pe_b/peij_0_3/add/fai_4/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_5/U4  ( .A(
        \pool/pool/pe_b_o_data[0][5] ), .B(
        \pool/pool/pe_b/peij_0_3/add/notb [5]), .Z(
        \pool/pool/pe_b/peij_0_3/add/fai_5/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_5/U3  ( .A(
        \pool/pool/pe_b/peij_0_3/add/cprop [5]), .B(
        \pool/pool/pe_b/peij_0_3/add/fai_5/n3 ), .Z(
        \pool/pool/pe_b/peij_0_3/d_acc [5]) );
  INV_X2 \pool/pool/pe_b/peij_0_3/add/fai_5/U2  ( .A(
        \pool/pool/pe_b/peij_0_3/add/fai_5/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_3/add/cprop [6]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_3/add/fai_5/U1  ( .A1(
        \pool/pool/pe_b/peij_0_3/add/notb [5]), .A2(
        \pool/pool/pe_b_o_data[0][5] ), .B1(
        \pool/pool/pe_b/peij_0_3/add/fai_5/n3 ), .B2(
        \pool/pool/pe_b/peij_0_3/add/cprop [5]), .ZN(
        \pool/pool/pe_b/peij_0_3/add/fai_5/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_6/U4  ( .A(
        \pool/pool/pe_b_o_data[0][6] ), .B(
        \pool/pool/pe_b/peij_0_3/add/notb [6]), .Z(
        \pool/pool/pe_b/peij_0_3/add/fai_6/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_6/U3  ( .A(
        \pool/pool/pe_b/peij_0_3/add/cprop [6]), .B(
        \pool/pool/pe_b/peij_0_3/add/fai_6/n3 ), .Z(
        \pool/pool/pe_b/peij_0_3/d_acc [6]) );
  INV_X2 \pool/pool/pe_b/peij_0_3/add/fai_6/U2  ( .A(
        \pool/pool/pe_b/peij_0_3/add/fai_6/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_3/add/cprop [7]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_3/add/fai_6/U1  ( .A1(
        \pool/pool/pe_b/peij_0_3/add/notb [6]), .A2(
        \pool/pool/pe_b_o_data[0][6] ), .B1(
        \pool/pool/pe_b/peij_0_3/add/fai_6/n3 ), .B2(
        \pool/pool/pe_b/peij_0_3/add/cprop [6]), .ZN(
        \pool/pool/pe_b/peij_0_3/add/fai_6/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_7/U4  ( .A(
        \pool/pool/pe_b_o_data[0][7] ), .B(
        \pool/pool/pe_b/peij_0_3/add/notb [7]), .Z(
        \pool/pool/pe_b/peij_0_3/add/fai_7/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_7/U3  ( .A(
        \pool/pool/pe_b/peij_0_3/add/cprop [7]), .B(
        \pool/pool/pe_b/peij_0_3/add/fai_7/n3 ), .Z(
        \pool/pool/pe_b/peij_0_3/d_acc [7]) );
  INV_X2 \pool/pool/pe_b/peij_0_3/add/fai_7/U2  ( .A(
        \pool/pool/pe_b/peij_0_3/add/fai_7/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_3/add/cprop [8]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_3/add/fai_7/U1  ( .A1(
        \pool/pool/pe_b/peij_0_3/add/notb [7]), .A2(
        \pool/pool/pe_b_o_data[0][7] ), .B1(
        \pool/pool/pe_b/peij_0_3/add/fai_7/n3 ), .B2(
        \pool/pool/pe_b/peij_0_3/add/cprop [7]), .ZN(
        \pool/pool/pe_b/peij_0_3/add/fai_7/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_8/U4  ( .A(
        \pool/pool/pe_b_o_data[0][8] ), .B(
        \pool/pool/pe_b/peij_0_3/add/notb [8]), .Z(
        \pool/pool/pe_b/peij_0_3/add/fai_8/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_8/U3  ( .A(
        \pool/pool/pe_b/peij_0_3/add/cprop [8]), .B(
        \pool/pool/pe_b/peij_0_3/add/fai_8/n3 ), .Z(
        \pool/pool/pe_b/peij_0_3/d_acc [8]) );
  INV_X2 \pool/pool/pe_b/peij_0_3/add/fai_8/U2  ( .A(
        \pool/pool/pe_b/peij_0_3/add/fai_8/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_3/add/cprop [9]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_3/add/fai_8/U1  ( .A1(
        \pool/pool/pe_b/peij_0_3/add/notb [8]), .A2(
        \pool/pool/pe_b_o_data[0][8] ), .B1(
        \pool/pool/pe_b/peij_0_3/add/fai_8/n3 ), .B2(
        \pool/pool/pe_b/peij_0_3/add/cprop [8]), .ZN(
        \pool/pool/pe_b/peij_0_3/add/fai_8/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_9/U4  ( .A(
        \pool/pool/pe_b_o_data[0][9] ), .B(
        \pool/pool/pe_b/peij_0_3/add/notb [9]), .Z(
        \pool/pool/pe_b/peij_0_3/add/fai_9/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_9/U3  ( .A(
        \pool/pool/pe_b/peij_0_3/add/cprop [9]), .B(
        \pool/pool/pe_b/peij_0_3/add/fai_9/n3 ), .Z(
        \pool/pool/pe_b/peij_0_3/d_acc [9]) );
  INV_X2 \pool/pool/pe_b/peij_0_3/add/fai_9/U2  ( .A(
        \pool/pool/pe_b/peij_0_3/add/fai_9/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_3/add/cprop [10]) );
  AOI22_X2 \pool/pool/pe_b/peij_0_3/add/fai_9/U1  ( .A1(
        \pool/pool/pe_b/peij_0_3/add/notb [9]), .A2(
        \pool/pool/pe_b_o_data[0][9] ), .B1(
        \pool/pool/pe_b/peij_0_3/add/fai_9/n3 ), .B2(
        \pool/pool/pe_b/peij_0_3/add/cprop [9]), .ZN(
        \pool/pool/pe_b/peij_0_3/add/fai_9/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_10/U4  ( .A(
        \pool/pool/pe_b_o_data[0][10] ), .B(
        \pool/pool/pe_b/peij_0_3/add/notb [10]), .Z(
        \pool/pool/pe_b/peij_0_3/add/fai_10/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_0_3/add/fai_10/U3  ( .A(
        \pool/pool/pe_b/peij_0_3/add/cprop [10]), .B(
        \pool/pool/pe_b/peij_0_3/add/fai_10/n3 ), .Z(
        \pool/pool/pe_b/peij_0_3/d_acc [10]) );
  INV_X2 \pool/pool/pe_b/peij_0_3/add/fai_10/U2  ( .A(
        \pool/pool/pe_b/peij_0_3/add/fai_10/n1 ), .ZN(
        \pool/pool/pe_b/peij_0_3/add/c_out ) );
  AOI22_X2 \pool/pool/pe_b/peij_0_3/add/fai_10/U1  ( .A1(
        \pool/pool/pe_b/peij_0_3/add/notb [10]), .A2(
        \pool/pool/pe_b_o_data[0][10] ), .B1(
        \pool/pool/pe_b/peij_0_3/add/fai_10/n3 ), .B2(
        \pool/pool/pe_b/peij_0_3/add/cprop [10]), .ZN(
        \pool/pool/pe_b/peij_0_3/add/fai_10/n1 ) );
  INV_X1 \pool/pool/pe_b/peij_1_0/U22  ( .A(\pool/pool/pe_b/n6 ), .ZN(
        \pool/pool/pe_b/peij_1_0/n16 ) );
  INV_X1 \pool/pool/pe_b/peij_1_0/U14  ( .A(\pool/pool/pe_b/n6 ), .ZN(
        \pool/pool/pe_b/peij_1_0/n12 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_0/U13  ( .A1(
        \pool/pool/pe_b/peij_1_0/d_acc [0]), .A2(\pool/pool/pe_b/peij_1_0/n18 ), .ZN(\pool/pool/pe_b/peij_1_0/n11 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_0/U12  ( .A1(
        \pool/pool/pe_b/peij_1_0/d_acc [1]), .A2(\pool/pool/pe_b/peij_1_0/n18 ), .ZN(\pool/pool/pe_b/peij_1_0/n10 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_0/U11  ( .A1(
        \pool/pool/pe_b/peij_1_0/d_acc [2]), .A2(\pool/pool/pe_b/peij_1_0/n18 ), .ZN(\pool/pool/pe_b/peij_1_0/n9 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_0/U10  ( .A1(
        \pool/pool/pe_b/peij_1_0/d_acc [3]), .A2(\pool/pool/pe_b/peij_1_0/n18 ), .ZN(\pool/pool/pe_b/peij_1_0/n8 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_0/U9  ( .A1(
        \pool/pool/pe_b/peij_1_0/d_acc [4]), .A2(\pool/pool/pe_b/peij_1_0/n18 ), .ZN(\pool/pool/pe_b/peij_1_0/n7 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_0/U8  ( .A1(
        \pool/pool/pe_b/peij_1_0/d_acc [5]), .A2(\pool/pool/pe_b/peij_1_0/n18 ), .ZN(\pool/pool/pe_b/peij_1_0/n6 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_0/U7  ( .A1(
        \pool/pool/pe_b/peij_1_0/d_acc [6]), .A2(\pool/pool/pe_b/peij_1_0/n18 ), .ZN(\pool/pool/pe_b/peij_1_0/n5 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_0/U6  ( .A1(
        \pool/pool/pe_b/peij_1_0/d_acc [7]), .A2(\pool/pool/pe_b/peij_1_0/n18 ), .ZN(\pool/pool/pe_b/peij_1_0/n4 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_0/U5  ( .A1(
        \pool/pool/pe_b/peij_1_0/d_acc [8]), .A2(\pool/pool/pe_b/peij_1_0/n18 ), .ZN(\pool/pool/pe_b/peij_1_0/n3 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_0/U4  ( .A1(
        \pool/pool/pe_b/peij_1_0/d_acc [9]), .A2(\pool/pool/pe_b/peij_1_0/n18 ), .ZN(\pool/pool/pe_b/peij_1_0/n2 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_0/U3  ( .A1(
        \pool/pool/pe_b/peij_1_0/d_acc [10]), .A2(
        \pool/pool/pe_b/peij_1_0/n18 ), .ZN(\pool/pool/pe_b/peij_1_0/n1 ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_0/q_acc_reg[10]  ( .D(
        \pool/pool/pe_b/peij_1_0/n1 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_0/n16 ), .Q(\pool/pool/pe_b_o_data[1][43] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_0/q_acc_reg[9]  ( .D(
        \pool/pool/pe_b/peij_1_0/n2 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_0/n16 ), .Q(\pool/pool/pe_b_o_data[1][42] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_0/q_acc_reg[8]  ( .D(
        \pool/pool/pe_b/peij_1_0/n3 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_0/n16 ), .Q(\pool/pool/pe_b_o_data[1][41] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_0/q_acc_reg[7]  ( .D(
        \pool/pool/pe_b/peij_1_0/n4 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_0/n16 ), .Q(\pool/pool/pe_b_o_data[1][40] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_0/q_acc_reg[6]  ( .D(
        \pool/pool/pe_b/peij_1_0/n5 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_0/n16 ), .Q(\pool/pool/pe_b_o_data[1][39] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_0/q_acc_reg[5]  ( .D(
        \pool/pool/pe_b/peij_1_0/n6 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_0/n16 ), .Q(\pool/pool/pe_b_o_data[1][38] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_0/q_acc_reg[4]  ( .D(
        \pool/pool/pe_b/peij_1_0/n7 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_0/n16 ), .Q(\pool/pool/pe_b_o_data[1][37] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_0/q_acc_reg[3]  ( .D(
        \pool/pool/pe_b/peij_1_0/n8 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_0/n16 ), .Q(\pool/pool/pe_b_o_data[1][36] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_0/q_acc_reg[2]  ( .D(
        \pool/pool/pe_b/peij_1_0/n9 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_0/n16 ), .Q(\pool/pool/pe_b_o_data[1][35] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_0/q_acc_reg[1]  ( .D(
        \pool/pool/pe_b/peij_1_0/n10 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_0/n16 ), .Q(\pool/pool/pe_b_o_data[1][34] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_0/q_acc_reg[0]  ( .D(
        \pool/pool/pe_b/peij_1_0/n11 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_0/n16 ), .Q(\pool/pool/pe_b_o_data[1][33] ) );
  INV_X2 \pool/pool/pe_b/peij_1_0/U21  ( .A(\pool/sync_clr ), .ZN(
        \pool/pool/pe_b/peij_1_0/n18 ) );
  AND3_X2 \pool/pool/pe_b/peij_1_0/U20  ( .A1(\pool/pool/pe_b/int_pe_en[1][0] ), .A2(\pool/pool/pe_b/peij_1_0/n18 ), .A3(1'b1), .ZN(
        \pool/pool/pe_b/peij_1_0/n17 ) );
  AND2_X2 \pool/pool/pe_b/peij_1_0/U19  ( .A1(\pool/pool/pe_b_i_data[1][12] ), 
        .A2(\pool/pool/pe_b/peij_1_0/n17 ), .ZN(\pool/pool/pe_b/peij_1_0/N33 )
         );
  AND2_X2 \pool/pool/pe_b/peij_1_0/U18  ( .A1(\pool/pool/pe_b_i_data[1][13] ), 
        .A2(\pool/pool/pe_b/peij_1_0/n17 ), .ZN(\pool/pool/pe_b/peij_1_0/N34 )
         );
  AND2_X2 \pool/pool/pe_b/peij_1_0/U17  ( .A1(\pool/pool/pe_b_i_data[1][14] ), 
        .A2(\pool/pool/pe_b/peij_1_0/n17 ), .ZN(\pool/pool/pe_b/peij_1_0/N35 )
         );
  AND4_X4 \pool/pool/pe_b/peij_1_0/U16  ( .A1(1'b1), .A2(
        \pool/pool/pe_b_i_data[1][15] ), .A3(\pool/pool/pe_b/int_pe_en[1][0] ), 
        .A4(\pool/pool/pe_b/peij_1_0/n18 ), .ZN(\pool/pool/pe_b/peij_1_0/N36 )
         );
  DFFR_X1 \pool/pool/pe_b/peij_1_0/q_im_reg[0]  ( .D(
        \pool/pool/pe_b/peij_1_0/N33 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_0/n12 ), .Q(\pool/pool/pe_b/peij_1_0/sgnext [0]) );
  DFFR_X1 \pool/pool/pe_b/peij_1_0/q_im_reg[1]  ( .D(
        \pool/pool/pe_b/peij_1_0/N34 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_0/n12 ), .Q(\pool/pool/pe_b/peij_1_0/sgnext [1]) );
  DFFR_X1 \pool/pool/pe_b/peij_1_0/q_im_reg[2]  ( .D(
        \pool/pool/pe_b/peij_1_0/N35 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_0/n12 ), .Q(\pool/pool/pe_b/peij_1_0/sgnext [2]) );
  DFFR_X1 \pool/pool/pe_b/peij_1_0/q_im_reg[3]  ( .D(
        \pool/pool/pe_b/peij_1_0/N36 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_0/n12 ), .Q(\pool/pool/pe_b/peij_1_0/sgnext_10 ) );
  SDFFR_X1 \pool/pool/pe_b/peij_1_0/q_k_reg  ( .D(1'b0), .SI(
        \pool/pool/pe_b/peij_1_0/n18 ), .SE(1'b0), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_0/n12 ), .Q(\pool/pool/pe_b/peij_1_0/q_k ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/U11  ( .A(
        \pool/pool/pe_b/peij_1_0/sgnext [0]), .B(\pool/pool/pe_b/peij_1_0/q_k ), .Z(\pool/pool/pe_b/peij_1_0/add/notb [0]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/U10  ( .A(
        \pool/pool/pe_b/peij_1_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_0/q_k ), .Z(\pool/pool/pe_b/peij_1_0/add/notb [10]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/U9  ( .A(
        \pool/pool/pe_b/peij_1_0/sgnext [1]), .B(\pool/pool/pe_b/peij_1_0/q_k ), .Z(\pool/pool/pe_b/peij_1_0/add/notb [1]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/U8  ( .A(
        \pool/pool/pe_b/peij_1_0/sgnext [2]), .B(\pool/pool/pe_b/peij_1_0/q_k ), .Z(\pool/pool/pe_b/peij_1_0/add/notb [2]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/U7  ( .A(
        \pool/pool/pe_b/peij_1_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_0/q_k ), .Z(\pool/pool/pe_b/peij_1_0/add/notb [3]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/U6  ( .A(
        \pool/pool/pe_b/peij_1_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_0/q_k ), .Z(\pool/pool/pe_b/peij_1_0/add/notb [4]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/U5  ( .A(
        \pool/pool/pe_b/peij_1_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_0/q_k ), .Z(\pool/pool/pe_b/peij_1_0/add/notb [5]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/U4  ( .A(
        \pool/pool/pe_b/peij_1_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_0/q_k ), .Z(\pool/pool/pe_b/peij_1_0/add/notb [6]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/U3  ( .A(
        \pool/pool/pe_b/peij_1_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_0/q_k ), .Z(\pool/pool/pe_b/peij_1_0/add/notb [7]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/U2  ( .A(
        \pool/pool/pe_b/peij_1_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_0/q_k ), .Z(\pool/pool/pe_b/peij_1_0/add/notb [8]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/U1  ( .A(
        \pool/pool/pe_b/peij_1_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_0/q_k ), .Z(\pool/pool/pe_b/peij_1_0/add/notb [9]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_0/U4  ( .A(
        \pool/pool/pe_b_o_data[1][33] ), .B(
        \pool/pool/pe_b/peij_1_0/add/notb [0]), .Z(
        \pool/pool/pe_b/peij_1_0/add/fai_0/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_0/U3  ( .A(
        \pool/pool/pe_b/peij_1_0/q_k ), .B(
        \pool/pool/pe_b/peij_1_0/add/fai_0/n3 ), .Z(
        \pool/pool/pe_b/peij_1_0/d_acc [0]) );
  INV_X2 \pool/pool/pe_b/peij_1_0/add/fai_0/U2  ( .A(
        \pool/pool/pe_b/peij_1_0/add/fai_0/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_0/add/cprop [1]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_0/add/fai_0/U1  ( .A1(
        \pool/pool/pe_b/peij_1_0/add/notb [0]), .A2(
        \pool/pool/pe_b_o_data[1][33] ), .B1(
        \pool/pool/pe_b/peij_1_0/add/fai_0/n3 ), .B2(
        \pool/pool/pe_b/peij_1_0/q_k ), .ZN(
        \pool/pool/pe_b/peij_1_0/add/fai_0/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_1/U4  ( .A(
        \pool/pool/pe_b_o_data[1][34] ), .B(
        \pool/pool/pe_b/peij_1_0/add/notb [1]), .Z(
        \pool/pool/pe_b/peij_1_0/add/fai_1/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_1/U3  ( .A(
        \pool/pool/pe_b/peij_1_0/add/cprop [1]), .B(
        \pool/pool/pe_b/peij_1_0/add/fai_1/n3 ), .Z(
        \pool/pool/pe_b/peij_1_0/d_acc [1]) );
  INV_X2 \pool/pool/pe_b/peij_1_0/add/fai_1/U2  ( .A(
        \pool/pool/pe_b/peij_1_0/add/fai_1/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_0/add/cprop [2]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_0/add/fai_1/U1  ( .A1(
        \pool/pool/pe_b/peij_1_0/add/notb [1]), .A2(
        \pool/pool/pe_b_o_data[1][34] ), .B1(
        \pool/pool/pe_b/peij_1_0/add/fai_1/n3 ), .B2(
        \pool/pool/pe_b/peij_1_0/add/cprop [1]), .ZN(
        \pool/pool/pe_b/peij_1_0/add/fai_1/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_2/U4  ( .A(
        \pool/pool/pe_b_o_data[1][35] ), .B(
        \pool/pool/pe_b/peij_1_0/add/notb [2]), .Z(
        \pool/pool/pe_b/peij_1_0/add/fai_2/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_2/U3  ( .A(
        \pool/pool/pe_b/peij_1_0/add/cprop [2]), .B(
        \pool/pool/pe_b/peij_1_0/add/fai_2/n3 ), .Z(
        \pool/pool/pe_b/peij_1_0/d_acc [2]) );
  INV_X2 \pool/pool/pe_b/peij_1_0/add/fai_2/U2  ( .A(
        \pool/pool/pe_b/peij_1_0/add/fai_2/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_0/add/cprop [3]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_0/add/fai_2/U1  ( .A1(
        \pool/pool/pe_b/peij_1_0/add/notb [2]), .A2(
        \pool/pool/pe_b_o_data[1][35] ), .B1(
        \pool/pool/pe_b/peij_1_0/add/fai_2/n3 ), .B2(
        \pool/pool/pe_b/peij_1_0/add/cprop [2]), .ZN(
        \pool/pool/pe_b/peij_1_0/add/fai_2/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_3/U4  ( .A(
        \pool/pool/pe_b_o_data[1][36] ), .B(
        \pool/pool/pe_b/peij_1_0/add/notb [3]), .Z(
        \pool/pool/pe_b/peij_1_0/add/fai_3/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_3/U3  ( .A(
        \pool/pool/pe_b/peij_1_0/add/cprop [3]), .B(
        \pool/pool/pe_b/peij_1_0/add/fai_3/n3 ), .Z(
        \pool/pool/pe_b/peij_1_0/d_acc [3]) );
  INV_X2 \pool/pool/pe_b/peij_1_0/add/fai_3/U2  ( .A(
        \pool/pool/pe_b/peij_1_0/add/fai_3/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_0/add/cprop [4]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_0/add/fai_3/U1  ( .A1(
        \pool/pool/pe_b/peij_1_0/add/notb [3]), .A2(
        \pool/pool/pe_b_o_data[1][36] ), .B1(
        \pool/pool/pe_b/peij_1_0/add/fai_3/n3 ), .B2(
        \pool/pool/pe_b/peij_1_0/add/cprop [3]), .ZN(
        \pool/pool/pe_b/peij_1_0/add/fai_3/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_4/U4  ( .A(
        \pool/pool/pe_b_o_data[1][37] ), .B(
        \pool/pool/pe_b/peij_1_0/add/notb [4]), .Z(
        \pool/pool/pe_b/peij_1_0/add/fai_4/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_4/U3  ( .A(
        \pool/pool/pe_b/peij_1_0/add/cprop [4]), .B(
        \pool/pool/pe_b/peij_1_0/add/fai_4/n3 ), .Z(
        \pool/pool/pe_b/peij_1_0/d_acc [4]) );
  INV_X2 \pool/pool/pe_b/peij_1_0/add/fai_4/U2  ( .A(
        \pool/pool/pe_b/peij_1_0/add/fai_4/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_0/add/cprop [5]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_0/add/fai_4/U1  ( .A1(
        \pool/pool/pe_b/peij_1_0/add/notb [4]), .A2(
        \pool/pool/pe_b_o_data[1][37] ), .B1(
        \pool/pool/pe_b/peij_1_0/add/fai_4/n3 ), .B2(
        \pool/pool/pe_b/peij_1_0/add/cprop [4]), .ZN(
        \pool/pool/pe_b/peij_1_0/add/fai_4/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_5/U4  ( .A(
        \pool/pool/pe_b_o_data[1][38] ), .B(
        \pool/pool/pe_b/peij_1_0/add/notb [5]), .Z(
        \pool/pool/pe_b/peij_1_0/add/fai_5/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_5/U3  ( .A(
        \pool/pool/pe_b/peij_1_0/add/cprop [5]), .B(
        \pool/pool/pe_b/peij_1_0/add/fai_5/n3 ), .Z(
        \pool/pool/pe_b/peij_1_0/d_acc [5]) );
  INV_X2 \pool/pool/pe_b/peij_1_0/add/fai_5/U2  ( .A(
        \pool/pool/pe_b/peij_1_0/add/fai_5/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_0/add/cprop [6]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_0/add/fai_5/U1  ( .A1(
        \pool/pool/pe_b/peij_1_0/add/notb [5]), .A2(
        \pool/pool/pe_b_o_data[1][38] ), .B1(
        \pool/pool/pe_b/peij_1_0/add/fai_5/n3 ), .B2(
        \pool/pool/pe_b/peij_1_0/add/cprop [5]), .ZN(
        \pool/pool/pe_b/peij_1_0/add/fai_5/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_6/U4  ( .A(
        \pool/pool/pe_b_o_data[1][39] ), .B(
        \pool/pool/pe_b/peij_1_0/add/notb [6]), .Z(
        \pool/pool/pe_b/peij_1_0/add/fai_6/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_6/U3  ( .A(
        \pool/pool/pe_b/peij_1_0/add/cprop [6]), .B(
        \pool/pool/pe_b/peij_1_0/add/fai_6/n3 ), .Z(
        \pool/pool/pe_b/peij_1_0/d_acc [6]) );
  INV_X2 \pool/pool/pe_b/peij_1_0/add/fai_6/U2  ( .A(
        \pool/pool/pe_b/peij_1_0/add/fai_6/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_0/add/cprop [7]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_0/add/fai_6/U1  ( .A1(
        \pool/pool/pe_b/peij_1_0/add/notb [6]), .A2(
        \pool/pool/pe_b_o_data[1][39] ), .B1(
        \pool/pool/pe_b/peij_1_0/add/fai_6/n3 ), .B2(
        \pool/pool/pe_b/peij_1_0/add/cprop [6]), .ZN(
        \pool/pool/pe_b/peij_1_0/add/fai_6/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_7/U4  ( .A(
        \pool/pool/pe_b_o_data[1][40] ), .B(
        \pool/pool/pe_b/peij_1_0/add/notb [7]), .Z(
        \pool/pool/pe_b/peij_1_0/add/fai_7/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_7/U3  ( .A(
        \pool/pool/pe_b/peij_1_0/add/cprop [7]), .B(
        \pool/pool/pe_b/peij_1_0/add/fai_7/n3 ), .Z(
        \pool/pool/pe_b/peij_1_0/d_acc [7]) );
  INV_X2 \pool/pool/pe_b/peij_1_0/add/fai_7/U2  ( .A(
        \pool/pool/pe_b/peij_1_0/add/fai_7/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_0/add/cprop [8]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_0/add/fai_7/U1  ( .A1(
        \pool/pool/pe_b/peij_1_0/add/notb [7]), .A2(
        \pool/pool/pe_b_o_data[1][40] ), .B1(
        \pool/pool/pe_b/peij_1_0/add/fai_7/n3 ), .B2(
        \pool/pool/pe_b/peij_1_0/add/cprop [7]), .ZN(
        \pool/pool/pe_b/peij_1_0/add/fai_7/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_8/U4  ( .A(
        \pool/pool/pe_b_o_data[1][41] ), .B(
        \pool/pool/pe_b/peij_1_0/add/notb [8]), .Z(
        \pool/pool/pe_b/peij_1_0/add/fai_8/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_8/U3  ( .A(
        \pool/pool/pe_b/peij_1_0/add/cprop [8]), .B(
        \pool/pool/pe_b/peij_1_0/add/fai_8/n3 ), .Z(
        \pool/pool/pe_b/peij_1_0/d_acc [8]) );
  INV_X2 \pool/pool/pe_b/peij_1_0/add/fai_8/U2  ( .A(
        \pool/pool/pe_b/peij_1_0/add/fai_8/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_0/add/cprop [9]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_0/add/fai_8/U1  ( .A1(
        \pool/pool/pe_b/peij_1_0/add/notb [8]), .A2(
        \pool/pool/pe_b_o_data[1][41] ), .B1(
        \pool/pool/pe_b/peij_1_0/add/fai_8/n3 ), .B2(
        \pool/pool/pe_b/peij_1_0/add/cprop [8]), .ZN(
        \pool/pool/pe_b/peij_1_0/add/fai_8/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_9/U4  ( .A(
        \pool/pool/pe_b_o_data[1][42] ), .B(
        \pool/pool/pe_b/peij_1_0/add/notb [9]), .Z(
        \pool/pool/pe_b/peij_1_0/add/fai_9/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_9/U3  ( .A(
        \pool/pool/pe_b/peij_1_0/add/cprop [9]), .B(
        \pool/pool/pe_b/peij_1_0/add/fai_9/n3 ), .Z(
        \pool/pool/pe_b/peij_1_0/d_acc [9]) );
  INV_X2 \pool/pool/pe_b/peij_1_0/add/fai_9/U2  ( .A(
        \pool/pool/pe_b/peij_1_0/add/fai_9/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_0/add/cprop [10]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_0/add/fai_9/U1  ( .A1(
        \pool/pool/pe_b/peij_1_0/add/notb [9]), .A2(
        \pool/pool/pe_b_o_data[1][42] ), .B1(
        \pool/pool/pe_b/peij_1_0/add/fai_9/n3 ), .B2(
        \pool/pool/pe_b/peij_1_0/add/cprop [9]), .ZN(
        \pool/pool/pe_b/peij_1_0/add/fai_9/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_10/U4  ( .A(
        \pool/pool/pe_b_o_data[1][43] ), .B(
        \pool/pool/pe_b/peij_1_0/add/notb [10]), .Z(
        \pool/pool/pe_b/peij_1_0/add/fai_10/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_0/add/fai_10/U3  ( .A(
        \pool/pool/pe_b/peij_1_0/add/cprop [10]), .B(
        \pool/pool/pe_b/peij_1_0/add/fai_10/n3 ), .Z(
        \pool/pool/pe_b/peij_1_0/d_acc [10]) );
  INV_X2 \pool/pool/pe_b/peij_1_0/add/fai_10/U2  ( .A(
        \pool/pool/pe_b/peij_1_0/add/fai_10/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_0/add/c_out ) );
  AOI22_X2 \pool/pool/pe_b/peij_1_0/add/fai_10/U1  ( .A1(
        \pool/pool/pe_b/peij_1_0/add/notb [10]), .A2(
        \pool/pool/pe_b_o_data[1][43] ), .B1(
        \pool/pool/pe_b/peij_1_0/add/fai_10/n3 ), .B2(
        \pool/pool/pe_b/peij_1_0/add/cprop [10]), .ZN(
        \pool/pool/pe_b/peij_1_0/add/fai_10/n1 ) );
  INV_X1 \pool/pool/pe_b/peij_1_1/U22  ( .A(\pool/pool/pe_b/n6 ), .ZN(
        \pool/pool/pe_b/peij_1_1/n16 ) );
  INV_X1 \pool/pool/pe_b/peij_1_1/U14  ( .A(\pool/pool/pe_b/n6 ), .ZN(
        \pool/pool/pe_b/peij_1_1/n12 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_1/U13  ( .A1(
        \pool/pool/pe_b/peij_1_1/d_acc [0]), .A2(\pool/pool/pe_b/peij_1_1/n18 ), .ZN(\pool/pool/pe_b/peij_1_1/n11 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_1/U12  ( .A1(
        \pool/pool/pe_b/peij_1_1/d_acc [1]), .A2(\pool/pool/pe_b/peij_1_1/n18 ), .ZN(\pool/pool/pe_b/peij_1_1/n10 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_1/U11  ( .A1(
        \pool/pool/pe_b/peij_1_1/d_acc [2]), .A2(\pool/pool/pe_b/peij_1_1/n18 ), .ZN(\pool/pool/pe_b/peij_1_1/n9 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_1/U10  ( .A1(
        \pool/pool/pe_b/peij_1_1/d_acc [3]), .A2(\pool/pool/pe_b/peij_1_1/n18 ), .ZN(\pool/pool/pe_b/peij_1_1/n8 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_1/U9  ( .A1(
        \pool/pool/pe_b/peij_1_1/d_acc [4]), .A2(\pool/pool/pe_b/peij_1_1/n18 ), .ZN(\pool/pool/pe_b/peij_1_1/n7 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_1/U8  ( .A1(
        \pool/pool/pe_b/peij_1_1/d_acc [5]), .A2(\pool/pool/pe_b/peij_1_1/n18 ), .ZN(\pool/pool/pe_b/peij_1_1/n6 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_1/U7  ( .A1(
        \pool/pool/pe_b/peij_1_1/d_acc [6]), .A2(\pool/pool/pe_b/peij_1_1/n18 ), .ZN(\pool/pool/pe_b/peij_1_1/n5 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_1/U6  ( .A1(
        \pool/pool/pe_b/peij_1_1/d_acc [7]), .A2(\pool/pool/pe_b/peij_1_1/n18 ), .ZN(\pool/pool/pe_b/peij_1_1/n4 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_1/U5  ( .A1(
        \pool/pool/pe_b/peij_1_1/d_acc [8]), .A2(\pool/pool/pe_b/peij_1_1/n18 ), .ZN(\pool/pool/pe_b/peij_1_1/n3 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_1/U4  ( .A1(
        \pool/pool/pe_b/peij_1_1/d_acc [9]), .A2(\pool/pool/pe_b/peij_1_1/n18 ), .ZN(\pool/pool/pe_b/peij_1_1/n2 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_1/U3  ( .A1(
        \pool/pool/pe_b/peij_1_1/d_acc [10]), .A2(
        \pool/pool/pe_b/peij_1_1/n18 ), .ZN(\pool/pool/pe_b/peij_1_1/n1 ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_1/q_acc_reg[10]  ( .D(
        \pool/pool/pe_b/peij_1_1/n1 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_1/n16 ), .Q(\pool/pool/pe_b_o_data[1][32] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_1/q_acc_reg[9]  ( .D(
        \pool/pool/pe_b/peij_1_1/n2 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_1/n16 ), .Q(\pool/pool/pe_b_o_data[1][31] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_1/q_acc_reg[8]  ( .D(
        \pool/pool/pe_b/peij_1_1/n3 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_1/n16 ), .Q(\pool/pool/pe_b_o_data[1][30] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_1/q_acc_reg[7]  ( .D(
        \pool/pool/pe_b/peij_1_1/n4 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_1/n16 ), .Q(\pool/pool/pe_b_o_data[1][29] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_1/q_acc_reg[6]  ( .D(
        \pool/pool/pe_b/peij_1_1/n5 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_1/n16 ), .Q(\pool/pool/pe_b_o_data[1][28] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_1/q_acc_reg[5]  ( .D(
        \pool/pool/pe_b/peij_1_1/n6 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_1/n16 ), .Q(\pool/pool/pe_b_o_data[1][27] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_1/q_acc_reg[4]  ( .D(
        \pool/pool/pe_b/peij_1_1/n7 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_1/n16 ), .Q(\pool/pool/pe_b_o_data[1][26] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_1/q_acc_reg[3]  ( .D(
        \pool/pool/pe_b/peij_1_1/n8 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_1/n16 ), .Q(\pool/pool/pe_b_o_data[1][25] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_1/q_acc_reg[2]  ( .D(
        \pool/pool/pe_b/peij_1_1/n9 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_1/n16 ), .Q(\pool/pool/pe_b_o_data[1][24] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_1/q_acc_reg[1]  ( .D(
        \pool/pool/pe_b/peij_1_1/n10 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_1/n16 ), .Q(\pool/pool/pe_b_o_data[1][23] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_1/q_acc_reg[0]  ( .D(
        \pool/pool/pe_b/peij_1_1/n11 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_1/n16 ), .Q(\pool/pool/pe_b_o_data[1][22] ) );
  INV_X2 \pool/pool/pe_b/peij_1_1/U21  ( .A(\pool/sync_clr ), .ZN(
        \pool/pool/pe_b/peij_1_1/n18 ) );
  AND3_X2 \pool/pool/pe_b/peij_1_1/U20  ( .A1(\pool/pool/pe_b/int_pe_en[1][1] ), .A2(\pool/pool/pe_b/peij_1_1/n18 ), .A3(1'b1), .ZN(
        \pool/pool/pe_b/peij_1_1/n17 ) );
  AND2_X2 \pool/pool/pe_b/peij_1_1/U19  ( .A1(\pool/pool/pe_b_i_data[1][8] ), 
        .A2(\pool/pool/pe_b/peij_1_1/n17 ), .ZN(\pool/pool/pe_b/peij_1_1/N33 )
         );
  AND2_X2 \pool/pool/pe_b/peij_1_1/U18  ( .A1(\pool/pool/pe_b_i_data[1][9] ), 
        .A2(\pool/pool/pe_b/peij_1_1/n17 ), .ZN(\pool/pool/pe_b/peij_1_1/N34 )
         );
  AND2_X2 \pool/pool/pe_b/peij_1_1/U17  ( .A1(\pool/pool/pe_b_i_data[1][10] ), 
        .A2(\pool/pool/pe_b/peij_1_1/n17 ), .ZN(\pool/pool/pe_b/peij_1_1/N35 )
         );
  AND4_X4 \pool/pool/pe_b/peij_1_1/U16  ( .A1(1'b1), .A2(
        \pool/pool/pe_b_i_data[1][11] ), .A3(\pool/pool/pe_b/int_pe_en[1][1] ), 
        .A4(\pool/pool/pe_b/peij_1_1/n18 ), .ZN(\pool/pool/pe_b/peij_1_1/N36 )
         );
  DFFR_X1 \pool/pool/pe_b/peij_1_1/q_im_reg[0]  ( .D(
        \pool/pool/pe_b/peij_1_1/N33 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_1/n12 ), .Q(\pool/pool/pe_b/peij_1_1/sgnext [0]) );
  DFFR_X1 \pool/pool/pe_b/peij_1_1/q_im_reg[1]  ( .D(
        \pool/pool/pe_b/peij_1_1/N34 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_1/n12 ), .Q(\pool/pool/pe_b/peij_1_1/sgnext [1]) );
  DFFR_X1 \pool/pool/pe_b/peij_1_1/q_im_reg[2]  ( .D(
        \pool/pool/pe_b/peij_1_1/N35 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_1/n12 ), .Q(\pool/pool/pe_b/peij_1_1/sgnext [2]) );
  DFFR_X1 \pool/pool/pe_b/peij_1_1/q_im_reg[3]  ( .D(
        \pool/pool/pe_b/peij_1_1/N36 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_1/n12 ), .Q(\pool/pool/pe_b/peij_1_1/sgnext_10 ) );
  SDFFR_X1 \pool/pool/pe_b/peij_1_1/q_k_reg  ( .D(1'b0), .SI(
        \pool/pool/pe_b/peij_1_1/n18 ), .SE(1'b0), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_1/n12 ), .Q(\pool/pool/pe_b/peij_1_1/q_k ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/U11  ( .A(
        \pool/pool/pe_b/peij_1_1/sgnext [0]), .B(\pool/pool/pe_b/peij_1_1/q_k ), .Z(\pool/pool/pe_b/peij_1_1/add/notb [0]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/U10  ( .A(
        \pool/pool/pe_b/peij_1_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_1/q_k ), .Z(\pool/pool/pe_b/peij_1_1/add/notb [10]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/U9  ( .A(
        \pool/pool/pe_b/peij_1_1/sgnext [1]), .B(\pool/pool/pe_b/peij_1_1/q_k ), .Z(\pool/pool/pe_b/peij_1_1/add/notb [1]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/U8  ( .A(
        \pool/pool/pe_b/peij_1_1/sgnext [2]), .B(\pool/pool/pe_b/peij_1_1/q_k ), .Z(\pool/pool/pe_b/peij_1_1/add/notb [2]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/U7  ( .A(
        \pool/pool/pe_b/peij_1_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_1/q_k ), .Z(\pool/pool/pe_b/peij_1_1/add/notb [3]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/U6  ( .A(
        \pool/pool/pe_b/peij_1_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_1/q_k ), .Z(\pool/pool/pe_b/peij_1_1/add/notb [4]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/U5  ( .A(
        \pool/pool/pe_b/peij_1_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_1/q_k ), .Z(\pool/pool/pe_b/peij_1_1/add/notb [5]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/U4  ( .A(
        \pool/pool/pe_b/peij_1_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_1/q_k ), .Z(\pool/pool/pe_b/peij_1_1/add/notb [6]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/U3  ( .A(
        \pool/pool/pe_b/peij_1_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_1/q_k ), .Z(\pool/pool/pe_b/peij_1_1/add/notb [7]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/U2  ( .A(
        \pool/pool/pe_b/peij_1_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_1/q_k ), .Z(\pool/pool/pe_b/peij_1_1/add/notb [8]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/U1  ( .A(
        \pool/pool/pe_b/peij_1_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_1/q_k ), .Z(\pool/pool/pe_b/peij_1_1/add/notb [9]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_0/U4  ( .A(
        \pool/pool/pe_b_o_data[1][22] ), .B(
        \pool/pool/pe_b/peij_1_1/add/notb [0]), .Z(
        \pool/pool/pe_b/peij_1_1/add/fai_0/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_0/U3  ( .A(
        \pool/pool/pe_b/peij_1_1/q_k ), .B(
        \pool/pool/pe_b/peij_1_1/add/fai_0/n3 ), .Z(
        \pool/pool/pe_b/peij_1_1/d_acc [0]) );
  INV_X2 \pool/pool/pe_b/peij_1_1/add/fai_0/U2  ( .A(
        \pool/pool/pe_b/peij_1_1/add/fai_0/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_1/add/cprop [1]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_1/add/fai_0/U1  ( .A1(
        \pool/pool/pe_b/peij_1_1/add/notb [0]), .A2(
        \pool/pool/pe_b_o_data[1][22] ), .B1(
        \pool/pool/pe_b/peij_1_1/add/fai_0/n3 ), .B2(
        \pool/pool/pe_b/peij_1_1/q_k ), .ZN(
        \pool/pool/pe_b/peij_1_1/add/fai_0/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_1/U4  ( .A(
        \pool/pool/pe_b_o_data[1][23] ), .B(
        \pool/pool/pe_b/peij_1_1/add/notb [1]), .Z(
        \pool/pool/pe_b/peij_1_1/add/fai_1/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_1/U3  ( .A(
        \pool/pool/pe_b/peij_1_1/add/cprop [1]), .B(
        \pool/pool/pe_b/peij_1_1/add/fai_1/n3 ), .Z(
        \pool/pool/pe_b/peij_1_1/d_acc [1]) );
  INV_X2 \pool/pool/pe_b/peij_1_1/add/fai_1/U2  ( .A(
        \pool/pool/pe_b/peij_1_1/add/fai_1/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_1/add/cprop [2]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_1/add/fai_1/U1  ( .A1(
        \pool/pool/pe_b/peij_1_1/add/notb [1]), .A2(
        \pool/pool/pe_b_o_data[1][23] ), .B1(
        \pool/pool/pe_b/peij_1_1/add/fai_1/n3 ), .B2(
        \pool/pool/pe_b/peij_1_1/add/cprop [1]), .ZN(
        \pool/pool/pe_b/peij_1_1/add/fai_1/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_2/U4  ( .A(
        \pool/pool/pe_b_o_data[1][24] ), .B(
        \pool/pool/pe_b/peij_1_1/add/notb [2]), .Z(
        \pool/pool/pe_b/peij_1_1/add/fai_2/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_2/U3  ( .A(
        \pool/pool/pe_b/peij_1_1/add/cprop [2]), .B(
        \pool/pool/pe_b/peij_1_1/add/fai_2/n3 ), .Z(
        \pool/pool/pe_b/peij_1_1/d_acc [2]) );
  INV_X2 \pool/pool/pe_b/peij_1_1/add/fai_2/U2  ( .A(
        \pool/pool/pe_b/peij_1_1/add/fai_2/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_1/add/cprop [3]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_1/add/fai_2/U1  ( .A1(
        \pool/pool/pe_b/peij_1_1/add/notb [2]), .A2(
        \pool/pool/pe_b_o_data[1][24] ), .B1(
        \pool/pool/pe_b/peij_1_1/add/fai_2/n3 ), .B2(
        \pool/pool/pe_b/peij_1_1/add/cprop [2]), .ZN(
        \pool/pool/pe_b/peij_1_1/add/fai_2/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_3/U4  ( .A(
        \pool/pool/pe_b_o_data[1][25] ), .B(
        \pool/pool/pe_b/peij_1_1/add/notb [3]), .Z(
        \pool/pool/pe_b/peij_1_1/add/fai_3/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_3/U3  ( .A(
        \pool/pool/pe_b/peij_1_1/add/cprop [3]), .B(
        \pool/pool/pe_b/peij_1_1/add/fai_3/n3 ), .Z(
        \pool/pool/pe_b/peij_1_1/d_acc [3]) );
  INV_X2 \pool/pool/pe_b/peij_1_1/add/fai_3/U2  ( .A(
        \pool/pool/pe_b/peij_1_1/add/fai_3/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_1/add/cprop [4]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_1/add/fai_3/U1  ( .A1(
        \pool/pool/pe_b/peij_1_1/add/notb [3]), .A2(
        \pool/pool/pe_b_o_data[1][25] ), .B1(
        \pool/pool/pe_b/peij_1_1/add/fai_3/n3 ), .B2(
        \pool/pool/pe_b/peij_1_1/add/cprop [3]), .ZN(
        \pool/pool/pe_b/peij_1_1/add/fai_3/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_4/U4  ( .A(
        \pool/pool/pe_b_o_data[1][26] ), .B(
        \pool/pool/pe_b/peij_1_1/add/notb [4]), .Z(
        \pool/pool/pe_b/peij_1_1/add/fai_4/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_4/U3  ( .A(
        \pool/pool/pe_b/peij_1_1/add/cprop [4]), .B(
        \pool/pool/pe_b/peij_1_1/add/fai_4/n3 ), .Z(
        \pool/pool/pe_b/peij_1_1/d_acc [4]) );
  INV_X2 \pool/pool/pe_b/peij_1_1/add/fai_4/U2  ( .A(
        \pool/pool/pe_b/peij_1_1/add/fai_4/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_1/add/cprop [5]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_1/add/fai_4/U1  ( .A1(
        \pool/pool/pe_b/peij_1_1/add/notb [4]), .A2(
        \pool/pool/pe_b_o_data[1][26] ), .B1(
        \pool/pool/pe_b/peij_1_1/add/fai_4/n3 ), .B2(
        \pool/pool/pe_b/peij_1_1/add/cprop [4]), .ZN(
        \pool/pool/pe_b/peij_1_1/add/fai_4/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_5/U4  ( .A(
        \pool/pool/pe_b_o_data[1][27] ), .B(
        \pool/pool/pe_b/peij_1_1/add/notb [5]), .Z(
        \pool/pool/pe_b/peij_1_1/add/fai_5/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_5/U3  ( .A(
        \pool/pool/pe_b/peij_1_1/add/cprop [5]), .B(
        \pool/pool/pe_b/peij_1_1/add/fai_5/n3 ), .Z(
        \pool/pool/pe_b/peij_1_1/d_acc [5]) );
  INV_X2 \pool/pool/pe_b/peij_1_1/add/fai_5/U2  ( .A(
        \pool/pool/pe_b/peij_1_1/add/fai_5/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_1/add/cprop [6]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_1/add/fai_5/U1  ( .A1(
        \pool/pool/pe_b/peij_1_1/add/notb [5]), .A2(
        \pool/pool/pe_b_o_data[1][27] ), .B1(
        \pool/pool/pe_b/peij_1_1/add/fai_5/n3 ), .B2(
        \pool/pool/pe_b/peij_1_1/add/cprop [5]), .ZN(
        \pool/pool/pe_b/peij_1_1/add/fai_5/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_6/U4  ( .A(
        \pool/pool/pe_b_o_data[1][28] ), .B(
        \pool/pool/pe_b/peij_1_1/add/notb [6]), .Z(
        \pool/pool/pe_b/peij_1_1/add/fai_6/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_6/U3  ( .A(
        \pool/pool/pe_b/peij_1_1/add/cprop [6]), .B(
        \pool/pool/pe_b/peij_1_1/add/fai_6/n3 ), .Z(
        \pool/pool/pe_b/peij_1_1/d_acc [6]) );
  INV_X2 \pool/pool/pe_b/peij_1_1/add/fai_6/U2  ( .A(
        \pool/pool/pe_b/peij_1_1/add/fai_6/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_1/add/cprop [7]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_1/add/fai_6/U1  ( .A1(
        \pool/pool/pe_b/peij_1_1/add/notb [6]), .A2(
        \pool/pool/pe_b_o_data[1][28] ), .B1(
        \pool/pool/pe_b/peij_1_1/add/fai_6/n3 ), .B2(
        \pool/pool/pe_b/peij_1_1/add/cprop [6]), .ZN(
        \pool/pool/pe_b/peij_1_1/add/fai_6/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_7/U4  ( .A(
        \pool/pool/pe_b_o_data[1][29] ), .B(
        \pool/pool/pe_b/peij_1_1/add/notb [7]), .Z(
        \pool/pool/pe_b/peij_1_1/add/fai_7/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_7/U3  ( .A(
        \pool/pool/pe_b/peij_1_1/add/cprop [7]), .B(
        \pool/pool/pe_b/peij_1_1/add/fai_7/n3 ), .Z(
        \pool/pool/pe_b/peij_1_1/d_acc [7]) );
  INV_X2 \pool/pool/pe_b/peij_1_1/add/fai_7/U2  ( .A(
        \pool/pool/pe_b/peij_1_1/add/fai_7/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_1/add/cprop [8]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_1/add/fai_7/U1  ( .A1(
        \pool/pool/pe_b/peij_1_1/add/notb [7]), .A2(
        \pool/pool/pe_b_o_data[1][29] ), .B1(
        \pool/pool/pe_b/peij_1_1/add/fai_7/n3 ), .B2(
        \pool/pool/pe_b/peij_1_1/add/cprop [7]), .ZN(
        \pool/pool/pe_b/peij_1_1/add/fai_7/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_8/U4  ( .A(
        \pool/pool/pe_b_o_data[1][30] ), .B(
        \pool/pool/pe_b/peij_1_1/add/notb [8]), .Z(
        \pool/pool/pe_b/peij_1_1/add/fai_8/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_8/U3  ( .A(
        \pool/pool/pe_b/peij_1_1/add/cprop [8]), .B(
        \pool/pool/pe_b/peij_1_1/add/fai_8/n3 ), .Z(
        \pool/pool/pe_b/peij_1_1/d_acc [8]) );
  INV_X2 \pool/pool/pe_b/peij_1_1/add/fai_8/U2  ( .A(
        \pool/pool/pe_b/peij_1_1/add/fai_8/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_1/add/cprop [9]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_1/add/fai_8/U1  ( .A1(
        \pool/pool/pe_b/peij_1_1/add/notb [8]), .A2(
        \pool/pool/pe_b_o_data[1][30] ), .B1(
        \pool/pool/pe_b/peij_1_1/add/fai_8/n3 ), .B2(
        \pool/pool/pe_b/peij_1_1/add/cprop [8]), .ZN(
        \pool/pool/pe_b/peij_1_1/add/fai_8/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_9/U4  ( .A(
        \pool/pool/pe_b_o_data[1][31] ), .B(
        \pool/pool/pe_b/peij_1_1/add/notb [9]), .Z(
        \pool/pool/pe_b/peij_1_1/add/fai_9/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_9/U3  ( .A(
        \pool/pool/pe_b/peij_1_1/add/cprop [9]), .B(
        \pool/pool/pe_b/peij_1_1/add/fai_9/n3 ), .Z(
        \pool/pool/pe_b/peij_1_1/d_acc [9]) );
  INV_X2 \pool/pool/pe_b/peij_1_1/add/fai_9/U2  ( .A(
        \pool/pool/pe_b/peij_1_1/add/fai_9/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_1/add/cprop [10]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_1/add/fai_9/U1  ( .A1(
        \pool/pool/pe_b/peij_1_1/add/notb [9]), .A2(
        \pool/pool/pe_b_o_data[1][31] ), .B1(
        \pool/pool/pe_b/peij_1_1/add/fai_9/n3 ), .B2(
        \pool/pool/pe_b/peij_1_1/add/cprop [9]), .ZN(
        \pool/pool/pe_b/peij_1_1/add/fai_9/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_10/U4  ( .A(
        \pool/pool/pe_b_o_data[1][32] ), .B(
        \pool/pool/pe_b/peij_1_1/add/notb [10]), .Z(
        \pool/pool/pe_b/peij_1_1/add/fai_10/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_1/add/fai_10/U3  ( .A(
        \pool/pool/pe_b/peij_1_1/add/cprop [10]), .B(
        \pool/pool/pe_b/peij_1_1/add/fai_10/n3 ), .Z(
        \pool/pool/pe_b/peij_1_1/d_acc [10]) );
  INV_X2 \pool/pool/pe_b/peij_1_1/add/fai_10/U2  ( .A(
        \pool/pool/pe_b/peij_1_1/add/fai_10/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_1/add/c_out ) );
  AOI22_X2 \pool/pool/pe_b/peij_1_1/add/fai_10/U1  ( .A1(
        \pool/pool/pe_b/peij_1_1/add/notb [10]), .A2(
        \pool/pool/pe_b_o_data[1][32] ), .B1(
        \pool/pool/pe_b/peij_1_1/add/fai_10/n3 ), .B2(
        \pool/pool/pe_b/peij_1_1/add/cprop [10]), .ZN(
        \pool/pool/pe_b/peij_1_1/add/fai_10/n1 ) );
  INV_X1 \pool/pool/pe_b/peij_1_2/U22  ( .A(\pool/pool/pe_b/n6 ), .ZN(
        \pool/pool/pe_b/peij_1_2/n16 ) );
  INV_X1 \pool/pool/pe_b/peij_1_2/U14  ( .A(\pool/pool/pe_b/n6 ), .ZN(
        \pool/pool/pe_b/peij_1_2/n12 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_2/U13  ( .A1(
        \pool/pool/pe_b/peij_1_2/d_acc [0]), .A2(\pool/pool/pe_b/peij_1_2/n18 ), .ZN(\pool/pool/pe_b/peij_1_2/n11 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_2/U12  ( .A1(
        \pool/pool/pe_b/peij_1_2/d_acc [1]), .A2(\pool/pool/pe_b/peij_1_2/n18 ), .ZN(\pool/pool/pe_b/peij_1_2/n10 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_2/U11  ( .A1(
        \pool/pool/pe_b/peij_1_2/d_acc [2]), .A2(\pool/pool/pe_b/peij_1_2/n18 ), .ZN(\pool/pool/pe_b/peij_1_2/n9 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_2/U10  ( .A1(
        \pool/pool/pe_b/peij_1_2/d_acc [3]), .A2(\pool/pool/pe_b/peij_1_2/n18 ), .ZN(\pool/pool/pe_b/peij_1_2/n8 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_2/U9  ( .A1(
        \pool/pool/pe_b/peij_1_2/d_acc [4]), .A2(\pool/pool/pe_b/peij_1_2/n18 ), .ZN(\pool/pool/pe_b/peij_1_2/n7 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_2/U8  ( .A1(
        \pool/pool/pe_b/peij_1_2/d_acc [5]), .A2(\pool/pool/pe_b/peij_1_2/n18 ), .ZN(\pool/pool/pe_b/peij_1_2/n6 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_2/U7  ( .A1(
        \pool/pool/pe_b/peij_1_2/d_acc [6]), .A2(\pool/pool/pe_b/peij_1_2/n18 ), .ZN(\pool/pool/pe_b/peij_1_2/n5 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_2/U6  ( .A1(
        \pool/pool/pe_b/peij_1_2/d_acc [7]), .A2(\pool/pool/pe_b/peij_1_2/n18 ), .ZN(\pool/pool/pe_b/peij_1_2/n4 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_2/U5  ( .A1(
        \pool/pool/pe_b/peij_1_2/d_acc [8]), .A2(\pool/pool/pe_b/peij_1_2/n18 ), .ZN(\pool/pool/pe_b/peij_1_2/n3 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_2/U4  ( .A1(
        \pool/pool/pe_b/peij_1_2/d_acc [9]), .A2(\pool/pool/pe_b/peij_1_2/n18 ), .ZN(\pool/pool/pe_b/peij_1_2/n2 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_2/U3  ( .A1(
        \pool/pool/pe_b/peij_1_2/d_acc [10]), .A2(
        \pool/pool/pe_b/peij_1_2/n18 ), .ZN(\pool/pool/pe_b/peij_1_2/n1 ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_2/q_acc_reg[10]  ( .D(
        \pool/pool/pe_b/peij_1_2/n1 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_2/n16 ), .Q(\pool/pool/pe_b_o_data[1][21] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_2/q_acc_reg[9]  ( .D(
        \pool/pool/pe_b/peij_1_2/n2 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_2/n16 ), .Q(\pool/pool/pe_b_o_data[1][20] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_2/q_acc_reg[8]  ( .D(
        \pool/pool/pe_b/peij_1_2/n3 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_2/n16 ), .Q(\pool/pool/pe_b_o_data[1][19] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_2/q_acc_reg[7]  ( .D(
        \pool/pool/pe_b/peij_1_2/n4 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_2/n16 ), .Q(\pool/pool/pe_b_o_data[1][18] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_2/q_acc_reg[6]  ( .D(
        \pool/pool/pe_b/peij_1_2/n5 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_2/n16 ), .Q(\pool/pool/pe_b_o_data[1][17] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_2/q_acc_reg[5]  ( .D(
        \pool/pool/pe_b/peij_1_2/n6 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_2/n16 ), .Q(\pool/pool/pe_b_o_data[1][16] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_2/q_acc_reg[4]  ( .D(
        \pool/pool/pe_b/peij_1_2/n7 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_2/n16 ), .Q(\pool/pool/pe_b_o_data[1][15] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_2/q_acc_reg[3]  ( .D(
        \pool/pool/pe_b/peij_1_2/n8 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_2/n16 ), .Q(\pool/pool/pe_b_o_data[1][14] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_2/q_acc_reg[2]  ( .D(
        \pool/pool/pe_b/peij_1_2/n9 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_2/n16 ), .Q(\pool/pool/pe_b_o_data[1][13] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_2/q_acc_reg[1]  ( .D(
        \pool/pool/pe_b/peij_1_2/n10 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_2/n16 ), .Q(\pool/pool/pe_b_o_data[1][12] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_2/q_acc_reg[0]  ( .D(
        \pool/pool/pe_b/peij_1_2/n11 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_2/n16 ), .Q(\pool/pool/pe_b_o_data[1][11] ) );
  INV_X2 \pool/pool/pe_b/peij_1_2/U21  ( .A(\pool/sync_clr ), .ZN(
        \pool/pool/pe_b/peij_1_2/n18 ) );
  AND3_X2 \pool/pool/pe_b/peij_1_2/U20  ( .A1(\pool/pool/pe_b/int_pe_en[1][2] ), .A2(\pool/pool/pe_b/peij_1_2/n18 ), .A3(1'b1), .ZN(
        \pool/pool/pe_b/peij_1_2/n17 ) );
  AND2_X2 \pool/pool/pe_b/peij_1_2/U19  ( .A1(\pool/pool/pe_b_i_data[1][4] ), 
        .A2(\pool/pool/pe_b/peij_1_2/n17 ), .ZN(\pool/pool/pe_b/peij_1_2/N33 )
         );
  AND2_X2 \pool/pool/pe_b/peij_1_2/U18  ( .A1(\pool/pool/pe_b_i_data[1][5] ), 
        .A2(\pool/pool/pe_b/peij_1_2/n17 ), .ZN(\pool/pool/pe_b/peij_1_2/N34 )
         );
  AND2_X2 \pool/pool/pe_b/peij_1_2/U17  ( .A1(\pool/pool/pe_b_i_data[1][6] ), 
        .A2(\pool/pool/pe_b/peij_1_2/n17 ), .ZN(\pool/pool/pe_b/peij_1_2/N35 )
         );
  AND4_X4 \pool/pool/pe_b/peij_1_2/U16  ( .A1(1'b1), .A2(
        \pool/pool/pe_b_i_data[1][7] ), .A3(\pool/pool/pe_b/int_pe_en[1][2] ), 
        .A4(\pool/pool/pe_b/peij_1_2/n18 ), .ZN(\pool/pool/pe_b/peij_1_2/N36 )
         );
  DFFR_X1 \pool/pool/pe_b/peij_1_2/q_im_reg[0]  ( .D(
        \pool/pool/pe_b/peij_1_2/N33 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_2/n12 ), .Q(\pool/pool/pe_b/peij_1_2/sgnext [0]) );
  DFFR_X1 \pool/pool/pe_b/peij_1_2/q_im_reg[1]  ( .D(
        \pool/pool/pe_b/peij_1_2/N34 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_2/n12 ), .Q(\pool/pool/pe_b/peij_1_2/sgnext [1]) );
  DFFR_X1 \pool/pool/pe_b/peij_1_2/q_im_reg[2]  ( .D(
        \pool/pool/pe_b/peij_1_2/N35 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_2/n12 ), .Q(\pool/pool/pe_b/peij_1_2/sgnext [2]) );
  DFFR_X1 \pool/pool/pe_b/peij_1_2/q_im_reg[3]  ( .D(
        \pool/pool/pe_b/peij_1_2/N36 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_2/n12 ), .Q(\pool/pool/pe_b/peij_1_2/sgnext_10 ) );
  SDFFR_X1 \pool/pool/pe_b/peij_1_2/q_k_reg  ( .D(1'b0), .SI(
        \pool/pool/pe_b/peij_1_2/n18 ), .SE(1'b0), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_2/n12 ), .Q(\pool/pool/pe_b/peij_1_2/q_k ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/U11  ( .A(
        \pool/pool/pe_b/peij_1_2/sgnext [0]), .B(\pool/pool/pe_b/peij_1_2/q_k ), .Z(\pool/pool/pe_b/peij_1_2/add/notb [0]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/U10  ( .A(
        \pool/pool/pe_b/peij_1_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_2/q_k ), .Z(\pool/pool/pe_b/peij_1_2/add/notb [10]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/U9  ( .A(
        \pool/pool/pe_b/peij_1_2/sgnext [1]), .B(\pool/pool/pe_b/peij_1_2/q_k ), .Z(\pool/pool/pe_b/peij_1_2/add/notb [1]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/U8  ( .A(
        \pool/pool/pe_b/peij_1_2/sgnext [2]), .B(\pool/pool/pe_b/peij_1_2/q_k ), .Z(\pool/pool/pe_b/peij_1_2/add/notb [2]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/U7  ( .A(
        \pool/pool/pe_b/peij_1_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_2/q_k ), .Z(\pool/pool/pe_b/peij_1_2/add/notb [3]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/U6  ( .A(
        \pool/pool/pe_b/peij_1_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_2/q_k ), .Z(\pool/pool/pe_b/peij_1_2/add/notb [4]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/U5  ( .A(
        \pool/pool/pe_b/peij_1_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_2/q_k ), .Z(\pool/pool/pe_b/peij_1_2/add/notb [5]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/U4  ( .A(
        \pool/pool/pe_b/peij_1_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_2/q_k ), .Z(\pool/pool/pe_b/peij_1_2/add/notb [6]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/U3  ( .A(
        \pool/pool/pe_b/peij_1_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_2/q_k ), .Z(\pool/pool/pe_b/peij_1_2/add/notb [7]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/U2  ( .A(
        \pool/pool/pe_b/peij_1_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_2/q_k ), .Z(\pool/pool/pe_b/peij_1_2/add/notb [8]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/U1  ( .A(
        \pool/pool/pe_b/peij_1_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_2/q_k ), .Z(\pool/pool/pe_b/peij_1_2/add/notb [9]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_0/U4  ( .A(
        \pool/pool/pe_b_o_data[1][11] ), .B(
        \pool/pool/pe_b/peij_1_2/add/notb [0]), .Z(
        \pool/pool/pe_b/peij_1_2/add/fai_0/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_0/U3  ( .A(
        \pool/pool/pe_b/peij_1_2/q_k ), .B(
        \pool/pool/pe_b/peij_1_2/add/fai_0/n3 ), .Z(
        \pool/pool/pe_b/peij_1_2/d_acc [0]) );
  INV_X2 \pool/pool/pe_b/peij_1_2/add/fai_0/U2  ( .A(
        \pool/pool/pe_b/peij_1_2/add/fai_0/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_2/add/cprop [1]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_2/add/fai_0/U1  ( .A1(
        \pool/pool/pe_b/peij_1_2/add/notb [0]), .A2(
        \pool/pool/pe_b_o_data[1][11] ), .B1(
        \pool/pool/pe_b/peij_1_2/add/fai_0/n3 ), .B2(
        \pool/pool/pe_b/peij_1_2/q_k ), .ZN(
        \pool/pool/pe_b/peij_1_2/add/fai_0/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_1/U4  ( .A(
        \pool/pool/pe_b_o_data[1][12] ), .B(
        \pool/pool/pe_b/peij_1_2/add/notb [1]), .Z(
        \pool/pool/pe_b/peij_1_2/add/fai_1/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_1/U3  ( .A(
        \pool/pool/pe_b/peij_1_2/add/cprop [1]), .B(
        \pool/pool/pe_b/peij_1_2/add/fai_1/n3 ), .Z(
        \pool/pool/pe_b/peij_1_2/d_acc [1]) );
  INV_X2 \pool/pool/pe_b/peij_1_2/add/fai_1/U2  ( .A(
        \pool/pool/pe_b/peij_1_2/add/fai_1/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_2/add/cprop [2]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_2/add/fai_1/U1  ( .A1(
        \pool/pool/pe_b/peij_1_2/add/notb [1]), .A2(
        \pool/pool/pe_b_o_data[1][12] ), .B1(
        \pool/pool/pe_b/peij_1_2/add/fai_1/n3 ), .B2(
        \pool/pool/pe_b/peij_1_2/add/cprop [1]), .ZN(
        \pool/pool/pe_b/peij_1_2/add/fai_1/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_2/U4  ( .A(
        \pool/pool/pe_b_o_data[1][13] ), .B(
        \pool/pool/pe_b/peij_1_2/add/notb [2]), .Z(
        \pool/pool/pe_b/peij_1_2/add/fai_2/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_2/U3  ( .A(
        \pool/pool/pe_b/peij_1_2/add/cprop [2]), .B(
        \pool/pool/pe_b/peij_1_2/add/fai_2/n3 ), .Z(
        \pool/pool/pe_b/peij_1_2/d_acc [2]) );
  INV_X2 \pool/pool/pe_b/peij_1_2/add/fai_2/U2  ( .A(
        \pool/pool/pe_b/peij_1_2/add/fai_2/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_2/add/cprop [3]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_2/add/fai_2/U1  ( .A1(
        \pool/pool/pe_b/peij_1_2/add/notb [2]), .A2(
        \pool/pool/pe_b_o_data[1][13] ), .B1(
        \pool/pool/pe_b/peij_1_2/add/fai_2/n3 ), .B2(
        \pool/pool/pe_b/peij_1_2/add/cprop [2]), .ZN(
        \pool/pool/pe_b/peij_1_2/add/fai_2/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_3/U4  ( .A(
        \pool/pool/pe_b_o_data[1][14] ), .B(
        \pool/pool/pe_b/peij_1_2/add/notb [3]), .Z(
        \pool/pool/pe_b/peij_1_2/add/fai_3/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_3/U3  ( .A(
        \pool/pool/pe_b/peij_1_2/add/cprop [3]), .B(
        \pool/pool/pe_b/peij_1_2/add/fai_3/n3 ), .Z(
        \pool/pool/pe_b/peij_1_2/d_acc [3]) );
  INV_X2 \pool/pool/pe_b/peij_1_2/add/fai_3/U2  ( .A(
        \pool/pool/pe_b/peij_1_2/add/fai_3/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_2/add/cprop [4]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_2/add/fai_3/U1  ( .A1(
        \pool/pool/pe_b/peij_1_2/add/notb [3]), .A2(
        \pool/pool/pe_b_o_data[1][14] ), .B1(
        \pool/pool/pe_b/peij_1_2/add/fai_3/n3 ), .B2(
        \pool/pool/pe_b/peij_1_2/add/cprop [3]), .ZN(
        \pool/pool/pe_b/peij_1_2/add/fai_3/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_4/U4  ( .A(
        \pool/pool/pe_b_o_data[1][15] ), .B(
        \pool/pool/pe_b/peij_1_2/add/notb [4]), .Z(
        \pool/pool/pe_b/peij_1_2/add/fai_4/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_4/U3  ( .A(
        \pool/pool/pe_b/peij_1_2/add/cprop [4]), .B(
        \pool/pool/pe_b/peij_1_2/add/fai_4/n3 ), .Z(
        \pool/pool/pe_b/peij_1_2/d_acc [4]) );
  INV_X2 \pool/pool/pe_b/peij_1_2/add/fai_4/U2  ( .A(
        \pool/pool/pe_b/peij_1_2/add/fai_4/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_2/add/cprop [5]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_2/add/fai_4/U1  ( .A1(
        \pool/pool/pe_b/peij_1_2/add/notb [4]), .A2(
        \pool/pool/pe_b_o_data[1][15] ), .B1(
        \pool/pool/pe_b/peij_1_2/add/fai_4/n3 ), .B2(
        \pool/pool/pe_b/peij_1_2/add/cprop [4]), .ZN(
        \pool/pool/pe_b/peij_1_2/add/fai_4/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_5/U4  ( .A(
        \pool/pool/pe_b_o_data[1][16] ), .B(
        \pool/pool/pe_b/peij_1_2/add/notb [5]), .Z(
        \pool/pool/pe_b/peij_1_2/add/fai_5/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_5/U3  ( .A(
        \pool/pool/pe_b/peij_1_2/add/cprop [5]), .B(
        \pool/pool/pe_b/peij_1_2/add/fai_5/n3 ), .Z(
        \pool/pool/pe_b/peij_1_2/d_acc [5]) );
  INV_X2 \pool/pool/pe_b/peij_1_2/add/fai_5/U2  ( .A(
        \pool/pool/pe_b/peij_1_2/add/fai_5/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_2/add/cprop [6]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_2/add/fai_5/U1  ( .A1(
        \pool/pool/pe_b/peij_1_2/add/notb [5]), .A2(
        \pool/pool/pe_b_o_data[1][16] ), .B1(
        \pool/pool/pe_b/peij_1_2/add/fai_5/n3 ), .B2(
        \pool/pool/pe_b/peij_1_2/add/cprop [5]), .ZN(
        \pool/pool/pe_b/peij_1_2/add/fai_5/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_6/U4  ( .A(
        \pool/pool/pe_b_o_data[1][17] ), .B(
        \pool/pool/pe_b/peij_1_2/add/notb [6]), .Z(
        \pool/pool/pe_b/peij_1_2/add/fai_6/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_6/U3  ( .A(
        \pool/pool/pe_b/peij_1_2/add/cprop [6]), .B(
        \pool/pool/pe_b/peij_1_2/add/fai_6/n3 ), .Z(
        \pool/pool/pe_b/peij_1_2/d_acc [6]) );
  INV_X2 \pool/pool/pe_b/peij_1_2/add/fai_6/U2  ( .A(
        \pool/pool/pe_b/peij_1_2/add/fai_6/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_2/add/cprop [7]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_2/add/fai_6/U1  ( .A1(
        \pool/pool/pe_b/peij_1_2/add/notb [6]), .A2(
        \pool/pool/pe_b_o_data[1][17] ), .B1(
        \pool/pool/pe_b/peij_1_2/add/fai_6/n3 ), .B2(
        \pool/pool/pe_b/peij_1_2/add/cprop [6]), .ZN(
        \pool/pool/pe_b/peij_1_2/add/fai_6/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_7/U4  ( .A(
        \pool/pool/pe_b_o_data[1][18] ), .B(
        \pool/pool/pe_b/peij_1_2/add/notb [7]), .Z(
        \pool/pool/pe_b/peij_1_2/add/fai_7/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_7/U3  ( .A(
        \pool/pool/pe_b/peij_1_2/add/cprop [7]), .B(
        \pool/pool/pe_b/peij_1_2/add/fai_7/n3 ), .Z(
        \pool/pool/pe_b/peij_1_2/d_acc [7]) );
  INV_X2 \pool/pool/pe_b/peij_1_2/add/fai_7/U2  ( .A(
        \pool/pool/pe_b/peij_1_2/add/fai_7/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_2/add/cprop [8]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_2/add/fai_7/U1  ( .A1(
        \pool/pool/pe_b/peij_1_2/add/notb [7]), .A2(
        \pool/pool/pe_b_o_data[1][18] ), .B1(
        \pool/pool/pe_b/peij_1_2/add/fai_7/n3 ), .B2(
        \pool/pool/pe_b/peij_1_2/add/cprop [7]), .ZN(
        \pool/pool/pe_b/peij_1_2/add/fai_7/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_8/U4  ( .A(
        \pool/pool/pe_b_o_data[1][19] ), .B(
        \pool/pool/pe_b/peij_1_2/add/notb [8]), .Z(
        \pool/pool/pe_b/peij_1_2/add/fai_8/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_8/U3  ( .A(
        \pool/pool/pe_b/peij_1_2/add/cprop [8]), .B(
        \pool/pool/pe_b/peij_1_2/add/fai_8/n3 ), .Z(
        \pool/pool/pe_b/peij_1_2/d_acc [8]) );
  INV_X2 \pool/pool/pe_b/peij_1_2/add/fai_8/U2  ( .A(
        \pool/pool/pe_b/peij_1_2/add/fai_8/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_2/add/cprop [9]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_2/add/fai_8/U1  ( .A1(
        \pool/pool/pe_b/peij_1_2/add/notb [8]), .A2(
        \pool/pool/pe_b_o_data[1][19] ), .B1(
        \pool/pool/pe_b/peij_1_2/add/fai_8/n3 ), .B2(
        \pool/pool/pe_b/peij_1_2/add/cprop [8]), .ZN(
        \pool/pool/pe_b/peij_1_2/add/fai_8/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_9/U4  ( .A(
        \pool/pool/pe_b_o_data[1][20] ), .B(
        \pool/pool/pe_b/peij_1_2/add/notb [9]), .Z(
        \pool/pool/pe_b/peij_1_2/add/fai_9/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_9/U3  ( .A(
        \pool/pool/pe_b/peij_1_2/add/cprop [9]), .B(
        \pool/pool/pe_b/peij_1_2/add/fai_9/n3 ), .Z(
        \pool/pool/pe_b/peij_1_2/d_acc [9]) );
  INV_X2 \pool/pool/pe_b/peij_1_2/add/fai_9/U2  ( .A(
        \pool/pool/pe_b/peij_1_2/add/fai_9/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_2/add/cprop [10]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_2/add/fai_9/U1  ( .A1(
        \pool/pool/pe_b/peij_1_2/add/notb [9]), .A2(
        \pool/pool/pe_b_o_data[1][20] ), .B1(
        \pool/pool/pe_b/peij_1_2/add/fai_9/n3 ), .B2(
        \pool/pool/pe_b/peij_1_2/add/cprop [9]), .ZN(
        \pool/pool/pe_b/peij_1_2/add/fai_9/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_10/U4  ( .A(
        \pool/pool/pe_b_o_data[1][21] ), .B(
        \pool/pool/pe_b/peij_1_2/add/notb [10]), .Z(
        \pool/pool/pe_b/peij_1_2/add/fai_10/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_2/add/fai_10/U3  ( .A(
        \pool/pool/pe_b/peij_1_2/add/cprop [10]), .B(
        \pool/pool/pe_b/peij_1_2/add/fai_10/n3 ), .Z(
        \pool/pool/pe_b/peij_1_2/d_acc [10]) );
  INV_X2 \pool/pool/pe_b/peij_1_2/add/fai_10/U2  ( .A(
        \pool/pool/pe_b/peij_1_2/add/fai_10/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_2/add/c_out ) );
  AOI22_X2 \pool/pool/pe_b/peij_1_2/add/fai_10/U1  ( .A1(
        \pool/pool/pe_b/peij_1_2/add/notb [10]), .A2(
        \pool/pool/pe_b_o_data[1][21] ), .B1(
        \pool/pool/pe_b/peij_1_2/add/fai_10/n3 ), .B2(
        \pool/pool/pe_b/peij_1_2/add/cprop [10]), .ZN(
        \pool/pool/pe_b/peij_1_2/add/fai_10/n1 ) );
  INV_X1 \pool/pool/pe_b/peij_1_3/U22  ( .A(\pool/pool/pe_b/n6 ), .ZN(
        \pool/pool/pe_b/peij_1_3/n16 ) );
  INV_X1 \pool/pool/pe_b/peij_1_3/U14  ( .A(\pool/pool/pe_b/n6 ), .ZN(
        \pool/pool/pe_b/peij_1_3/n12 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_3/U13  ( .A1(
        \pool/pool/pe_b/peij_1_3/d_acc [0]), .A2(\pool/pool/pe_b/peij_1_3/n18 ), .ZN(\pool/pool/pe_b/peij_1_3/n11 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_3/U12  ( .A1(
        \pool/pool/pe_b/peij_1_3/d_acc [1]), .A2(\pool/pool/pe_b/peij_1_3/n18 ), .ZN(\pool/pool/pe_b/peij_1_3/n10 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_3/U11  ( .A1(
        \pool/pool/pe_b/peij_1_3/d_acc [2]), .A2(\pool/pool/pe_b/peij_1_3/n18 ), .ZN(\pool/pool/pe_b/peij_1_3/n9 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_3/U10  ( .A1(
        \pool/pool/pe_b/peij_1_3/d_acc [3]), .A2(\pool/pool/pe_b/peij_1_3/n18 ), .ZN(\pool/pool/pe_b/peij_1_3/n8 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_3/U9  ( .A1(
        \pool/pool/pe_b/peij_1_3/d_acc [4]), .A2(\pool/pool/pe_b/peij_1_3/n18 ), .ZN(\pool/pool/pe_b/peij_1_3/n7 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_3/U8  ( .A1(
        \pool/pool/pe_b/peij_1_3/d_acc [5]), .A2(\pool/pool/pe_b/peij_1_3/n18 ), .ZN(\pool/pool/pe_b/peij_1_3/n6 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_3/U7  ( .A1(
        \pool/pool/pe_b/peij_1_3/d_acc [6]), .A2(\pool/pool/pe_b/peij_1_3/n18 ), .ZN(\pool/pool/pe_b/peij_1_3/n5 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_3/U6  ( .A1(
        \pool/pool/pe_b/peij_1_3/d_acc [7]), .A2(\pool/pool/pe_b/peij_1_3/n18 ), .ZN(\pool/pool/pe_b/peij_1_3/n4 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_3/U5  ( .A1(
        \pool/pool/pe_b/peij_1_3/d_acc [8]), .A2(\pool/pool/pe_b/peij_1_3/n18 ), .ZN(\pool/pool/pe_b/peij_1_3/n3 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_3/U4  ( .A1(
        \pool/pool/pe_b/peij_1_3/d_acc [9]), .A2(\pool/pool/pe_b/peij_1_3/n18 ), .ZN(\pool/pool/pe_b/peij_1_3/n2 ) );
  AND2_X1 \pool/pool/pe_b/peij_1_3/U3  ( .A1(
        \pool/pool/pe_b/peij_1_3/d_acc [10]), .A2(
        \pool/pool/pe_b/peij_1_3/n18 ), .ZN(\pool/pool/pe_b/peij_1_3/n1 ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_3/q_acc_reg[10]  ( .D(
        \pool/pool/pe_b/peij_1_3/n1 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_3/n16 ), .Q(\pool/pool/pe_b_o_data[1][10] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_3/q_acc_reg[9]  ( .D(
        \pool/pool/pe_b/peij_1_3/n2 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_3/n16 ), .Q(\pool/pool/pe_b_o_data[1][9] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_3/q_acc_reg[8]  ( .D(
        \pool/pool/pe_b/peij_1_3/n3 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_3/n16 ), .Q(\pool/pool/pe_b_o_data[1][8] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_3/q_acc_reg[7]  ( .D(
        \pool/pool/pe_b/peij_1_3/n4 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_3/n16 ), .Q(\pool/pool/pe_b_o_data[1][7] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_3/q_acc_reg[6]  ( .D(
        \pool/pool/pe_b/peij_1_3/n5 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_3/n16 ), .Q(\pool/pool/pe_b_o_data[1][6] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_3/q_acc_reg[5]  ( .D(
        \pool/pool/pe_b/peij_1_3/n6 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_3/n16 ), .Q(\pool/pool/pe_b_o_data[1][5] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_3/q_acc_reg[4]  ( .D(
        \pool/pool/pe_b/peij_1_3/n7 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_3/n16 ), .Q(\pool/pool/pe_b_o_data[1][4] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_3/q_acc_reg[3]  ( .D(
        \pool/pool/pe_b/peij_1_3/n8 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_3/n16 ), .Q(\pool/pool/pe_b_o_data[1][3] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_3/q_acc_reg[2]  ( .D(
        \pool/pool/pe_b/peij_1_3/n9 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_3/n16 ), .Q(\pool/pool/pe_b_o_data[1][2] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_3/q_acc_reg[1]  ( .D(
        \pool/pool/pe_b/peij_1_3/n10 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_3/n16 ), .Q(\pool/pool/pe_b_o_data[1][1] ) );
  DFFR_X1 \pool/pool/pe_b/peij_1_3/q_acc_reg[0]  ( .D(
        \pool/pool/pe_b/peij_1_3/n11 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_3/n16 ), .Q(\pool/pool/pe_b_o_data[1][0] ) );
  INV_X2 \pool/pool/pe_b/peij_1_3/U21  ( .A(\pool/sync_clr ), .ZN(
        \pool/pool/pe_b/peij_1_3/n18 ) );
  AND3_X2 \pool/pool/pe_b/peij_1_3/U20  ( .A1(\pool/pool/pe_b/int_pe_en[1][3] ), .A2(\pool/pool/pe_b/peij_1_3/n18 ), .A3(1'b1), .ZN(
        \pool/pool/pe_b/peij_1_3/n17 ) );
  AND2_X2 \pool/pool/pe_b/peij_1_3/U19  ( .A1(\pool/pool/pe_b_i_data[1][0] ), 
        .A2(\pool/pool/pe_b/peij_1_3/n17 ), .ZN(\pool/pool/pe_b/peij_1_3/N33 )
         );
  AND2_X2 \pool/pool/pe_b/peij_1_3/U18  ( .A1(\pool/pool/pe_b_i_data[1][1] ), 
        .A2(\pool/pool/pe_b/peij_1_3/n17 ), .ZN(\pool/pool/pe_b/peij_1_3/N34 )
         );
  AND2_X2 \pool/pool/pe_b/peij_1_3/U17  ( .A1(\pool/pool/pe_b_i_data[1][2] ), 
        .A2(\pool/pool/pe_b/peij_1_3/n17 ), .ZN(\pool/pool/pe_b/peij_1_3/N35 )
         );
  AND4_X4 \pool/pool/pe_b/peij_1_3/U16  ( .A1(1'b1), .A2(
        \pool/pool/pe_b_i_data[1][3] ), .A3(\pool/pool/pe_b/int_pe_en[1][3] ), 
        .A4(\pool/pool/pe_b/peij_1_3/n18 ), .ZN(\pool/pool/pe_b/peij_1_3/N36 )
         );
  DFFR_X1 \pool/pool/pe_b/peij_1_3/q_im_reg[0]  ( .D(
        \pool/pool/pe_b/peij_1_3/N33 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_3/n12 ), .Q(\pool/pool/pe_b/peij_1_3/sgnext [0]) );
  DFFR_X1 \pool/pool/pe_b/peij_1_3/q_im_reg[1]  ( .D(
        \pool/pool/pe_b/peij_1_3/N34 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_3/n12 ), .Q(\pool/pool/pe_b/peij_1_3/sgnext [1]) );
  DFFR_X1 \pool/pool/pe_b/peij_1_3/q_im_reg[2]  ( .D(
        \pool/pool/pe_b/peij_1_3/N35 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_3/n12 ), .Q(\pool/pool/pe_b/peij_1_3/sgnext [2]) );
  DFFR_X1 \pool/pool/pe_b/peij_1_3/q_im_reg[3]  ( .D(
        \pool/pool/pe_b/peij_1_3/N36 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_3/n12 ), .Q(\pool/pool/pe_b/peij_1_3/sgnext_10 ) );
  SDFFR_X1 \pool/pool/pe_b/peij_1_3/q_k_reg  ( .D(1'b0), .SI(
        \pool/pool/pe_b/peij_1_3/n18 ), .SE(1'b0), .CK(clk), .RN(
        \pool/pool/pe_b/peij_1_3/n12 ), .Q(\pool/pool/pe_b/peij_1_3/q_k ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/U11  ( .A(
        \pool/pool/pe_b/peij_1_3/sgnext [0]), .B(\pool/pool/pe_b/peij_1_3/q_k ), .Z(\pool/pool/pe_b/peij_1_3/add/notb [0]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/U10  ( .A(
        \pool/pool/pe_b/peij_1_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_3/q_k ), .Z(\pool/pool/pe_b/peij_1_3/add/notb [10]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/U9  ( .A(
        \pool/pool/pe_b/peij_1_3/sgnext [1]), .B(\pool/pool/pe_b/peij_1_3/q_k ), .Z(\pool/pool/pe_b/peij_1_3/add/notb [1]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/U8  ( .A(
        \pool/pool/pe_b/peij_1_3/sgnext [2]), .B(\pool/pool/pe_b/peij_1_3/q_k ), .Z(\pool/pool/pe_b/peij_1_3/add/notb [2]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/U7  ( .A(
        \pool/pool/pe_b/peij_1_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_3/q_k ), .Z(\pool/pool/pe_b/peij_1_3/add/notb [3]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/U6  ( .A(
        \pool/pool/pe_b/peij_1_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_3/q_k ), .Z(\pool/pool/pe_b/peij_1_3/add/notb [4]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/U5  ( .A(
        \pool/pool/pe_b/peij_1_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_3/q_k ), .Z(\pool/pool/pe_b/peij_1_3/add/notb [5]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/U4  ( .A(
        \pool/pool/pe_b/peij_1_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_3/q_k ), .Z(\pool/pool/pe_b/peij_1_3/add/notb [6]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/U3  ( .A(
        \pool/pool/pe_b/peij_1_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_3/q_k ), .Z(\pool/pool/pe_b/peij_1_3/add/notb [7]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/U2  ( .A(
        \pool/pool/pe_b/peij_1_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_3/q_k ), .Z(\pool/pool/pe_b/peij_1_3/add/notb [8]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/U1  ( .A(
        \pool/pool/pe_b/peij_1_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_1_3/q_k ), .Z(\pool/pool/pe_b/peij_1_3/add/notb [9]) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_0/U4  ( .A(
        \pool/pool/pe_b_o_data[1][0] ), .B(
        \pool/pool/pe_b/peij_1_3/add/notb [0]), .Z(
        \pool/pool/pe_b/peij_1_3/add/fai_0/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_0/U3  ( .A(
        \pool/pool/pe_b/peij_1_3/q_k ), .B(
        \pool/pool/pe_b/peij_1_3/add/fai_0/n3 ), .Z(
        \pool/pool/pe_b/peij_1_3/d_acc [0]) );
  INV_X2 \pool/pool/pe_b/peij_1_3/add/fai_0/U2  ( .A(
        \pool/pool/pe_b/peij_1_3/add/fai_0/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_3/add/cprop [1]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_3/add/fai_0/U1  ( .A1(
        \pool/pool/pe_b/peij_1_3/add/notb [0]), .A2(
        \pool/pool/pe_b_o_data[1][0] ), .B1(
        \pool/pool/pe_b/peij_1_3/add/fai_0/n3 ), .B2(
        \pool/pool/pe_b/peij_1_3/q_k ), .ZN(
        \pool/pool/pe_b/peij_1_3/add/fai_0/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_1/U4  ( .A(
        \pool/pool/pe_b_o_data[1][1] ), .B(
        \pool/pool/pe_b/peij_1_3/add/notb [1]), .Z(
        \pool/pool/pe_b/peij_1_3/add/fai_1/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_1/U3  ( .A(
        \pool/pool/pe_b/peij_1_3/add/cprop [1]), .B(
        \pool/pool/pe_b/peij_1_3/add/fai_1/n3 ), .Z(
        \pool/pool/pe_b/peij_1_3/d_acc [1]) );
  INV_X2 \pool/pool/pe_b/peij_1_3/add/fai_1/U2  ( .A(
        \pool/pool/pe_b/peij_1_3/add/fai_1/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_3/add/cprop [2]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_3/add/fai_1/U1  ( .A1(
        \pool/pool/pe_b/peij_1_3/add/notb [1]), .A2(
        \pool/pool/pe_b_o_data[1][1] ), .B1(
        \pool/pool/pe_b/peij_1_3/add/fai_1/n3 ), .B2(
        \pool/pool/pe_b/peij_1_3/add/cprop [1]), .ZN(
        \pool/pool/pe_b/peij_1_3/add/fai_1/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_2/U4  ( .A(
        \pool/pool/pe_b_o_data[1][2] ), .B(
        \pool/pool/pe_b/peij_1_3/add/notb [2]), .Z(
        \pool/pool/pe_b/peij_1_3/add/fai_2/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_2/U3  ( .A(
        \pool/pool/pe_b/peij_1_3/add/cprop [2]), .B(
        \pool/pool/pe_b/peij_1_3/add/fai_2/n3 ), .Z(
        \pool/pool/pe_b/peij_1_3/d_acc [2]) );
  INV_X2 \pool/pool/pe_b/peij_1_3/add/fai_2/U2  ( .A(
        \pool/pool/pe_b/peij_1_3/add/fai_2/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_3/add/cprop [3]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_3/add/fai_2/U1  ( .A1(
        \pool/pool/pe_b/peij_1_3/add/notb [2]), .A2(
        \pool/pool/pe_b_o_data[1][2] ), .B1(
        \pool/pool/pe_b/peij_1_3/add/fai_2/n3 ), .B2(
        \pool/pool/pe_b/peij_1_3/add/cprop [2]), .ZN(
        \pool/pool/pe_b/peij_1_3/add/fai_2/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_3/U4  ( .A(
        \pool/pool/pe_b_o_data[1][3] ), .B(
        \pool/pool/pe_b/peij_1_3/add/notb [3]), .Z(
        \pool/pool/pe_b/peij_1_3/add/fai_3/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_3/U3  ( .A(
        \pool/pool/pe_b/peij_1_3/add/cprop [3]), .B(
        \pool/pool/pe_b/peij_1_3/add/fai_3/n3 ), .Z(
        \pool/pool/pe_b/peij_1_3/d_acc [3]) );
  INV_X2 \pool/pool/pe_b/peij_1_3/add/fai_3/U2  ( .A(
        \pool/pool/pe_b/peij_1_3/add/fai_3/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_3/add/cprop [4]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_3/add/fai_3/U1  ( .A1(
        \pool/pool/pe_b/peij_1_3/add/notb [3]), .A2(
        \pool/pool/pe_b_o_data[1][3] ), .B1(
        \pool/pool/pe_b/peij_1_3/add/fai_3/n3 ), .B2(
        \pool/pool/pe_b/peij_1_3/add/cprop [3]), .ZN(
        \pool/pool/pe_b/peij_1_3/add/fai_3/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_4/U4  ( .A(
        \pool/pool/pe_b_o_data[1][4] ), .B(
        \pool/pool/pe_b/peij_1_3/add/notb [4]), .Z(
        \pool/pool/pe_b/peij_1_3/add/fai_4/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_4/U3  ( .A(
        \pool/pool/pe_b/peij_1_3/add/cprop [4]), .B(
        \pool/pool/pe_b/peij_1_3/add/fai_4/n3 ), .Z(
        \pool/pool/pe_b/peij_1_3/d_acc [4]) );
  INV_X2 \pool/pool/pe_b/peij_1_3/add/fai_4/U2  ( .A(
        \pool/pool/pe_b/peij_1_3/add/fai_4/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_3/add/cprop [5]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_3/add/fai_4/U1  ( .A1(
        \pool/pool/pe_b/peij_1_3/add/notb [4]), .A2(
        \pool/pool/pe_b_o_data[1][4] ), .B1(
        \pool/pool/pe_b/peij_1_3/add/fai_4/n3 ), .B2(
        \pool/pool/pe_b/peij_1_3/add/cprop [4]), .ZN(
        \pool/pool/pe_b/peij_1_3/add/fai_4/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_5/U4  ( .A(
        \pool/pool/pe_b_o_data[1][5] ), .B(
        \pool/pool/pe_b/peij_1_3/add/notb [5]), .Z(
        \pool/pool/pe_b/peij_1_3/add/fai_5/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_5/U3  ( .A(
        \pool/pool/pe_b/peij_1_3/add/cprop [5]), .B(
        \pool/pool/pe_b/peij_1_3/add/fai_5/n3 ), .Z(
        \pool/pool/pe_b/peij_1_3/d_acc [5]) );
  INV_X2 \pool/pool/pe_b/peij_1_3/add/fai_5/U2  ( .A(
        \pool/pool/pe_b/peij_1_3/add/fai_5/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_3/add/cprop [6]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_3/add/fai_5/U1  ( .A1(
        \pool/pool/pe_b/peij_1_3/add/notb [5]), .A2(
        \pool/pool/pe_b_o_data[1][5] ), .B1(
        \pool/pool/pe_b/peij_1_3/add/fai_5/n3 ), .B2(
        \pool/pool/pe_b/peij_1_3/add/cprop [5]), .ZN(
        \pool/pool/pe_b/peij_1_3/add/fai_5/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_6/U4  ( .A(
        \pool/pool/pe_b_o_data[1][6] ), .B(
        \pool/pool/pe_b/peij_1_3/add/notb [6]), .Z(
        \pool/pool/pe_b/peij_1_3/add/fai_6/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_6/U3  ( .A(
        \pool/pool/pe_b/peij_1_3/add/cprop [6]), .B(
        \pool/pool/pe_b/peij_1_3/add/fai_6/n3 ), .Z(
        \pool/pool/pe_b/peij_1_3/d_acc [6]) );
  INV_X2 \pool/pool/pe_b/peij_1_3/add/fai_6/U2  ( .A(
        \pool/pool/pe_b/peij_1_3/add/fai_6/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_3/add/cprop [7]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_3/add/fai_6/U1  ( .A1(
        \pool/pool/pe_b/peij_1_3/add/notb [6]), .A2(
        \pool/pool/pe_b_o_data[1][6] ), .B1(
        \pool/pool/pe_b/peij_1_3/add/fai_6/n3 ), .B2(
        \pool/pool/pe_b/peij_1_3/add/cprop [6]), .ZN(
        \pool/pool/pe_b/peij_1_3/add/fai_6/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_7/U4  ( .A(
        \pool/pool/pe_b_o_data[1][7] ), .B(
        \pool/pool/pe_b/peij_1_3/add/notb [7]), .Z(
        \pool/pool/pe_b/peij_1_3/add/fai_7/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_7/U3  ( .A(
        \pool/pool/pe_b/peij_1_3/add/cprop [7]), .B(
        \pool/pool/pe_b/peij_1_3/add/fai_7/n3 ), .Z(
        \pool/pool/pe_b/peij_1_3/d_acc [7]) );
  INV_X2 \pool/pool/pe_b/peij_1_3/add/fai_7/U2  ( .A(
        \pool/pool/pe_b/peij_1_3/add/fai_7/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_3/add/cprop [8]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_3/add/fai_7/U1  ( .A1(
        \pool/pool/pe_b/peij_1_3/add/notb [7]), .A2(
        \pool/pool/pe_b_o_data[1][7] ), .B1(
        \pool/pool/pe_b/peij_1_3/add/fai_7/n3 ), .B2(
        \pool/pool/pe_b/peij_1_3/add/cprop [7]), .ZN(
        \pool/pool/pe_b/peij_1_3/add/fai_7/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_8/U4  ( .A(
        \pool/pool/pe_b_o_data[1][8] ), .B(
        \pool/pool/pe_b/peij_1_3/add/notb [8]), .Z(
        \pool/pool/pe_b/peij_1_3/add/fai_8/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_8/U3  ( .A(
        \pool/pool/pe_b/peij_1_3/add/cprop [8]), .B(
        \pool/pool/pe_b/peij_1_3/add/fai_8/n3 ), .Z(
        \pool/pool/pe_b/peij_1_3/d_acc [8]) );
  INV_X2 \pool/pool/pe_b/peij_1_3/add/fai_8/U2  ( .A(
        \pool/pool/pe_b/peij_1_3/add/fai_8/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_3/add/cprop [9]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_3/add/fai_8/U1  ( .A1(
        \pool/pool/pe_b/peij_1_3/add/notb [8]), .A2(
        \pool/pool/pe_b_o_data[1][8] ), .B1(
        \pool/pool/pe_b/peij_1_3/add/fai_8/n3 ), .B2(
        \pool/pool/pe_b/peij_1_3/add/cprop [8]), .ZN(
        \pool/pool/pe_b/peij_1_3/add/fai_8/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_9/U4  ( .A(
        \pool/pool/pe_b_o_data[1][9] ), .B(
        \pool/pool/pe_b/peij_1_3/add/notb [9]), .Z(
        \pool/pool/pe_b/peij_1_3/add/fai_9/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_9/U3  ( .A(
        \pool/pool/pe_b/peij_1_3/add/cprop [9]), .B(
        \pool/pool/pe_b/peij_1_3/add/fai_9/n3 ), .Z(
        \pool/pool/pe_b/peij_1_3/d_acc [9]) );
  INV_X2 \pool/pool/pe_b/peij_1_3/add/fai_9/U2  ( .A(
        \pool/pool/pe_b/peij_1_3/add/fai_9/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_3/add/cprop [10]) );
  AOI22_X2 \pool/pool/pe_b/peij_1_3/add/fai_9/U1  ( .A1(
        \pool/pool/pe_b/peij_1_3/add/notb [9]), .A2(
        \pool/pool/pe_b_o_data[1][9] ), .B1(
        \pool/pool/pe_b/peij_1_3/add/fai_9/n3 ), .B2(
        \pool/pool/pe_b/peij_1_3/add/cprop [9]), .ZN(
        \pool/pool/pe_b/peij_1_3/add/fai_9/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_10/U4  ( .A(
        \pool/pool/pe_b_o_data[1][10] ), .B(
        \pool/pool/pe_b/peij_1_3/add/notb [10]), .Z(
        \pool/pool/pe_b/peij_1_3/add/fai_10/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_1_3/add/fai_10/U3  ( .A(
        \pool/pool/pe_b/peij_1_3/add/cprop [10]), .B(
        \pool/pool/pe_b/peij_1_3/add/fai_10/n3 ), .Z(
        \pool/pool/pe_b/peij_1_3/d_acc [10]) );
  INV_X2 \pool/pool/pe_b/peij_1_3/add/fai_10/U2  ( .A(
        \pool/pool/pe_b/peij_1_3/add/fai_10/n1 ), .ZN(
        \pool/pool/pe_b/peij_1_3/add/c_out ) );
  AOI22_X2 \pool/pool/pe_b/peij_1_3/add/fai_10/U1  ( .A1(
        \pool/pool/pe_b/peij_1_3/add/notb [10]), .A2(
        \pool/pool/pe_b_o_data[1][10] ), .B1(
        \pool/pool/pe_b/peij_1_3/add/fai_10/n3 ), .B2(
        \pool/pool/pe_b/peij_1_3/add/cprop [10]), .ZN(
        \pool/pool/pe_b/peij_1_3/add/fai_10/n1 ) );
  INV_X1 \pool/pool/pe_b/peij_2_0/U22  ( .A(\pool/pool/pe_b/n6 ), .ZN(
        \pool/pool/pe_b/peij_2_0/n16 ) );
  INV_X1 \pool/pool/pe_b/peij_2_0/U14  ( .A(\pool/pool/pe_b/n6 ), .ZN(
        \pool/pool/pe_b/peij_2_0/n12 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_0/U13  ( .A1(
        \pool/pool/pe_b/peij_2_0/d_acc [0]), .A2(\pool/pool/pe_b/peij_2_0/n18 ), .ZN(\pool/pool/pe_b/peij_2_0/n11 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_0/U12  ( .A1(
        \pool/pool/pe_b/peij_2_0/d_acc [1]), .A2(\pool/pool/pe_b/peij_2_0/n18 ), .ZN(\pool/pool/pe_b/peij_2_0/n10 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_0/U11  ( .A1(
        \pool/pool/pe_b/peij_2_0/d_acc [2]), .A2(\pool/pool/pe_b/peij_2_0/n18 ), .ZN(\pool/pool/pe_b/peij_2_0/n9 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_0/U10  ( .A1(
        \pool/pool/pe_b/peij_2_0/d_acc [3]), .A2(\pool/pool/pe_b/peij_2_0/n18 ), .ZN(\pool/pool/pe_b/peij_2_0/n8 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_0/U9  ( .A1(
        \pool/pool/pe_b/peij_2_0/d_acc [4]), .A2(\pool/pool/pe_b/peij_2_0/n18 ), .ZN(\pool/pool/pe_b/peij_2_0/n7 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_0/U8  ( .A1(
        \pool/pool/pe_b/peij_2_0/d_acc [5]), .A2(\pool/pool/pe_b/peij_2_0/n18 ), .ZN(\pool/pool/pe_b/peij_2_0/n6 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_0/U7  ( .A1(
        \pool/pool/pe_b/peij_2_0/d_acc [6]), .A2(\pool/pool/pe_b/peij_2_0/n18 ), .ZN(\pool/pool/pe_b/peij_2_0/n5 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_0/U6  ( .A1(
        \pool/pool/pe_b/peij_2_0/d_acc [7]), .A2(\pool/pool/pe_b/peij_2_0/n18 ), .ZN(\pool/pool/pe_b/peij_2_0/n4 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_0/U5  ( .A1(
        \pool/pool/pe_b/peij_2_0/d_acc [8]), .A2(\pool/pool/pe_b/peij_2_0/n18 ), .ZN(\pool/pool/pe_b/peij_2_0/n3 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_0/U4  ( .A1(
        \pool/pool/pe_b/peij_2_0/d_acc [9]), .A2(\pool/pool/pe_b/peij_2_0/n18 ), .ZN(\pool/pool/pe_b/peij_2_0/n2 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_0/U3  ( .A1(
        \pool/pool/pe_b/peij_2_0/d_acc [10]), .A2(
        \pool/pool/pe_b/peij_2_0/n18 ), .ZN(\pool/pool/pe_b/peij_2_0/n1 ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_0/q_acc_reg[10]  ( .D(
        \pool/pool/pe_b/peij_2_0/n1 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_0/n16 ), .Q(\pool/pool/pe_b_o_data[2][43] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_0/q_acc_reg[9]  ( .D(
        \pool/pool/pe_b/peij_2_0/n2 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_0/n16 ), .Q(\pool/pool/pe_b_o_data[2][42] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_0/q_acc_reg[8]  ( .D(
        \pool/pool/pe_b/peij_2_0/n3 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_0/n16 ), .Q(\pool/pool/pe_b_o_data[2][41] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_0/q_acc_reg[7]  ( .D(
        \pool/pool/pe_b/peij_2_0/n4 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_0/n16 ), .Q(\pool/pool/pe_b_o_data[2][40] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_0/q_acc_reg[6]  ( .D(
        \pool/pool/pe_b/peij_2_0/n5 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_0/n16 ), .Q(\pool/pool/pe_b_o_data[2][39] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_0/q_acc_reg[5]  ( .D(
        \pool/pool/pe_b/peij_2_0/n6 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_0/n16 ), .Q(\pool/pool/pe_b_o_data[2][38] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_0/q_acc_reg[4]  ( .D(
        \pool/pool/pe_b/peij_2_0/n7 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_0/n16 ), .Q(\pool/pool/pe_b_o_data[2][37] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_0/q_acc_reg[3]  ( .D(
        \pool/pool/pe_b/peij_2_0/n8 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_0/n16 ), .Q(\pool/pool/pe_b_o_data[2][36] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_0/q_acc_reg[2]  ( .D(
        \pool/pool/pe_b/peij_2_0/n9 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_0/n16 ), .Q(\pool/pool/pe_b_o_data[2][35] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_0/q_acc_reg[1]  ( .D(
        \pool/pool/pe_b/peij_2_0/n10 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_0/n16 ), .Q(\pool/pool/pe_b_o_data[2][34] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_0/q_acc_reg[0]  ( .D(
        \pool/pool/pe_b/peij_2_0/n11 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_0/n16 ), .Q(\pool/pool/pe_b_o_data[2][33] ) );
  INV_X2 \pool/pool/pe_b/peij_2_0/U21  ( .A(\pool/sync_clr ), .ZN(
        \pool/pool/pe_b/peij_2_0/n18 ) );
  AND3_X2 \pool/pool/pe_b/peij_2_0/U20  ( .A1(\pool/pool/pe_b/int_pe_en[2][0] ), .A2(\pool/pool/pe_b/peij_2_0/n18 ), .A3(1'b1), .ZN(
        \pool/pool/pe_b/peij_2_0/n17 ) );
  AND2_X2 \pool/pool/pe_b/peij_2_0/U19  ( .A1(\pool/pool/pe_b_i_data[2][12] ), 
        .A2(\pool/pool/pe_b/peij_2_0/n17 ), .ZN(\pool/pool/pe_b/peij_2_0/N33 )
         );
  AND2_X2 \pool/pool/pe_b/peij_2_0/U18  ( .A1(\pool/pool/pe_b_i_data[2][13] ), 
        .A2(\pool/pool/pe_b/peij_2_0/n17 ), .ZN(\pool/pool/pe_b/peij_2_0/N34 )
         );
  AND2_X2 \pool/pool/pe_b/peij_2_0/U17  ( .A1(\pool/pool/pe_b_i_data[2][14] ), 
        .A2(\pool/pool/pe_b/peij_2_0/n17 ), .ZN(\pool/pool/pe_b/peij_2_0/N35 )
         );
  AND4_X4 \pool/pool/pe_b/peij_2_0/U16  ( .A1(1'b1), .A2(
        \pool/pool/pe_b_i_data[2][15] ), .A3(\pool/pool/pe_b/int_pe_en[2][0] ), 
        .A4(\pool/pool/pe_b/peij_2_0/n18 ), .ZN(\pool/pool/pe_b/peij_2_0/N36 )
         );
  DFFR_X1 \pool/pool/pe_b/peij_2_0/q_im_reg[0]  ( .D(
        \pool/pool/pe_b/peij_2_0/N33 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_0/n12 ), .Q(\pool/pool/pe_b/peij_2_0/sgnext [0]) );
  DFFR_X1 \pool/pool/pe_b/peij_2_0/q_im_reg[1]  ( .D(
        \pool/pool/pe_b/peij_2_0/N34 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_0/n12 ), .Q(\pool/pool/pe_b/peij_2_0/sgnext [1]) );
  DFFR_X1 \pool/pool/pe_b/peij_2_0/q_im_reg[2]  ( .D(
        \pool/pool/pe_b/peij_2_0/N35 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_0/n12 ), .Q(\pool/pool/pe_b/peij_2_0/sgnext [2]) );
  DFFR_X1 \pool/pool/pe_b/peij_2_0/q_im_reg[3]  ( .D(
        \pool/pool/pe_b/peij_2_0/N36 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_0/n12 ), .Q(\pool/pool/pe_b/peij_2_0/sgnext_10 ) );
  SDFFR_X1 \pool/pool/pe_b/peij_2_0/q_k_reg  ( .D(1'b0), .SI(
        \pool/pool/pe_b/peij_2_0/n18 ), .SE(1'b0), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_0/n12 ), .Q(\pool/pool/pe_b/peij_2_0/q_k ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/U11  ( .A(
        \pool/pool/pe_b/peij_2_0/sgnext [0]), .B(\pool/pool/pe_b/peij_2_0/q_k ), .Z(\pool/pool/pe_b/peij_2_0/add/notb [0]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/U10  ( .A(
        \pool/pool/pe_b/peij_2_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_0/q_k ), .Z(\pool/pool/pe_b/peij_2_0/add/notb [10]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/U9  ( .A(
        \pool/pool/pe_b/peij_2_0/sgnext [1]), .B(\pool/pool/pe_b/peij_2_0/q_k ), .Z(\pool/pool/pe_b/peij_2_0/add/notb [1]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/U8  ( .A(
        \pool/pool/pe_b/peij_2_0/sgnext [2]), .B(\pool/pool/pe_b/peij_2_0/q_k ), .Z(\pool/pool/pe_b/peij_2_0/add/notb [2]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/U7  ( .A(
        \pool/pool/pe_b/peij_2_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_0/q_k ), .Z(\pool/pool/pe_b/peij_2_0/add/notb [3]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/U6  ( .A(
        \pool/pool/pe_b/peij_2_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_0/q_k ), .Z(\pool/pool/pe_b/peij_2_0/add/notb [4]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/U5  ( .A(
        \pool/pool/pe_b/peij_2_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_0/q_k ), .Z(\pool/pool/pe_b/peij_2_0/add/notb [5]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/U4  ( .A(
        \pool/pool/pe_b/peij_2_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_0/q_k ), .Z(\pool/pool/pe_b/peij_2_0/add/notb [6]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/U3  ( .A(
        \pool/pool/pe_b/peij_2_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_0/q_k ), .Z(\pool/pool/pe_b/peij_2_0/add/notb [7]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/U2  ( .A(
        \pool/pool/pe_b/peij_2_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_0/q_k ), .Z(\pool/pool/pe_b/peij_2_0/add/notb [8]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/U1  ( .A(
        \pool/pool/pe_b/peij_2_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_0/q_k ), .Z(\pool/pool/pe_b/peij_2_0/add/notb [9]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_0/U4  ( .A(
        \pool/pool/pe_b_o_data[2][33] ), .B(
        \pool/pool/pe_b/peij_2_0/add/notb [0]), .Z(
        \pool/pool/pe_b/peij_2_0/add/fai_0/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_0/U3  ( .A(
        \pool/pool/pe_b/peij_2_0/q_k ), .B(
        \pool/pool/pe_b/peij_2_0/add/fai_0/n3 ), .Z(
        \pool/pool/pe_b/peij_2_0/d_acc [0]) );
  INV_X2 \pool/pool/pe_b/peij_2_0/add/fai_0/U2  ( .A(
        \pool/pool/pe_b/peij_2_0/add/fai_0/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_0/add/cprop [1]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_0/add/fai_0/U1  ( .A1(
        \pool/pool/pe_b/peij_2_0/add/notb [0]), .A2(
        \pool/pool/pe_b_o_data[2][33] ), .B1(
        \pool/pool/pe_b/peij_2_0/add/fai_0/n3 ), .B2(
        \pool/pool/pe_b/peij_2_0/q_k ), .ZN(
        \pool/pool/pe_b/peij_2_0/add/fai_0/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_1/U4  ( .A(
        \pool/pool/pe_b_o_data[2][34] ), .B(
        \pool/pool/pe_b/peij_2_0/add/notb [1]), .Z(
        \pool/pool/pe_b/peij_2_0/add/fai_1/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_1/U3  ( .A(
        \pool/pool/pe_b/peij_2_0/add/cprop [1]), .B(
        \pool/pool/pe_b/peij_2_0/add/fai_1/n3 ), .Z(
        \pool/pool/pe_b/peij_2_0/d_acc [1]) );
  INV_X2 \pool/pool/pe_b/peij_2_0/add/fai_1/U2  ( .A(
        \pool/pool/pe_b/peij_2_0/add/fai_1/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_0/add/cprop [2]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_0/add/fai_1/U1  ( .A1(
        \pool/pool/pe_b/peij_2_0/add/notb [1]), .A2(
        \pool/pool/pe_b_o_data[2][34] ), .B1(
        \pool/pool/pe_b/peij_2_0/add/fai_1/n3 ), .B2(
        \pool/pool/pe_b/peij_2_0/add/cprop [1]), .ZN(
        \pool/pool/pe_b/peij_2_0/add/fai_1/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_2/U4  ( .A(
        \pool/pool/pe_b_o_data[2][35] ), .B(
        \pool/pool/pe_b/peij_2_0/add/notb [2]), .Z(
        \pool/pool/pe_b/peij_2_0/add/fai_2/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_2/U3  ( .A(
        \pool/pool/pe_b/peij_2_0/add/cprop [2]), .B(
        \pool/pool/pe_b/peij_2_0/add/fai_2/n3 ), .Z(
        \pool/pool/pe_b/peij_2_0/d_acc [2]) );
  INV_X2 \pool/pool/pe_b/peij_2_0/add/fai_2/U2  ( .A(
        \pool/pool/pe_b/peij_2_0/add/fai_2/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_0/add/cprop [3]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_0/add/fai_2/U1  ( .A1(
        \pool/pool/pe_b/peij_2_0/add/notb [2]), .A2(
        \pool/pool/pe_b_o_data[2][35] ), .B1(
        \pool/pool/pe_b/peij_2_0/add/fai_2/n3 ), .B2(
        \pool/pool/pe_b/peij_2_0/add/cprop [2]), .ZN(
        \pool/pool/pe_b/peij_2_0/add/fai_2/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_3/U4  ( .A(
        \pool/pool/pe_b_o_data[2][36] ), .B(
        \pool/pool/pe_b/peij_2_0/add/notb [3]), .Z(
        \pool/pool/pe_b/peij_2_0/add/fai_3/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_3/U3  ( .A(
        \pool/pool/pe_b/peij_2_0/add/cprop [3]), .B(
        \pool/pool/pe_b/peij_2_0/add/fai_3/n3 ), .Z(
        \pool/pool/pe_b/peij_2_0/d_acc [3]) );
  INV_X2 \pool/pool/pe_b/peij_2_0/add/fai_3/U2  ( .A(
        \pool/pool/pe_b/peij_2_0/add/fai_3/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_0/add/cprop [4]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_0/add/fai_3/U1  ( .A1(
        \pool/pool/pe_b/peij_2_0/add/notb [3]), .A2(
        \pool/pool/pe_b_o_data[2][36] ), .B1(
        \pool/pool/pe_b/peij_2_0/add/fai_3/n3 ), .B2(
        \pool/pool/pe_b/peij_2_0/add/cprop [3]), .ZN(
        \pool/pool/pe_b/peij_2_0/add/fai_3/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_4/U4  ( .A(
        \pool/pool/pe_b_o_data[2][37] ), .B(
        \pool/pool/pe_b/peij_2_0/add/notb [4]), .Z(
        \pool/pool/pe_b/peij_2_0/add/fai_4/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_4/U3  ( .A(
        \pool/pool/pe_b/peij_2_0/add/cprop [4]), .B(
        \pool/pool/pe_b/peij_2_0/add/fai_4/n3 ), .Z(
        \pool/pool/pe_b/peij_2_0/d_acc [4]) );
  INV_X2 \pool/pool/pe_b/peij_2_0/add/fai_4/U2  ( .A(
        \pool/pool/pe_b/peij_2_0/add/fai_4/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_0/add/cprop [5]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_0/add/fai_4/U1  ( .A1(
        \pool/pool/pe_b/peij_2_0/add/notb [4]), .A2(
        \pool/pool/pe_b_o_data[2][37] ), .B1(
        \pool/pool/pe_b/peij_2_0/add/fai_4/n3 ), .B2(
        \pool/pool/pe_b/peij_2_0/add/cprop [4]), .ZN(
        \pool/pool/pe_b/peij_2_0/add/fai_4/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_5/U4  ( .A(
        \pool/pool/pe_b_o_data[2][38] ), .B(
        \pool/pool/pe_b/peij_2_0/add/notb [5]), .Z(
        \pool/pool/pe_b/peij_2_0/add/fai_5/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_5/U3  ( .A(
        \pool/pool/pe_b/peij_2_0/add/cprop [5]), .B(
        \pool/pool/pe_b/peij_2_0/add/fai_5/n3 ), .Z(
        \pool/pool/pe_b/peij_2_0/d_acc [5]) );
  INV_X2 \pool/pool/pe_b/peij_2_0/add/fai_5/U2  ( .A(
        \pool/pool/pe_b/peij_2_0/add/fai_5/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_0/add/cprop [6]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_0/add/fai_5/U1  ( .A1(
        \pool/pool/pe_b/peij_2_0/add/notb [5]), .A2(
        \pool/pool/pe_b_o_data[2][38] ), .B1(
        \pool/pool/pe_b/peij_2_0/add/fai_5/n3 ), .B2(
        \pool/pool/pe_b/peij_2_0/add/cprop [5]), .ZN(
        \pool/pool/pe_b/peij_2_0/add/fai_5/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_6/U4  ( .A(
        \pool/pool/pe_b_o_data[2][39] ), .B(
        \pool/pool/pe_b/peij_2_0/add/notb [6]), .Z(
        \pool/pool/pe_b/peij_2_0/add/fai_6/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_6/U3  ( .A(
        \pool/pool/pe_b/peij_2_0/add/cprop [6]), .B(
        \pool/pool/pe_b/peij_2_0/add/fai_6/n3 ), .Z(
        \pool/pool/pe_b/peij_2_0/d_acc [6]) );
  INV_X2 \pool/pool/pe_b/peij_2_0/add/fai_6/U2  ( .A(
        \pool/pool/pe_b/peij_2_0/add/fai_6/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_0/add/cprop [7]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_0/add/fai_6/U1  ( .A1(
        \pool/pool/pe_b/peij_2_0/add/notb [6]), .A2(
        \pool/pool/pe_b_o_data[2][39] ), .B1(
        \pool/pool/pe_b/peij_2_0/add/fai_6/n3 ), .B2(
        \pool/pool/pe_b/peij_2_0/add/cprop [6]), .ZN(
        \pool/pool/pe_b/peij_2_0/add/fai_6/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_7/U4  ( .A(
        \pool/pool/pe_b_o_data[2][40] ), .B(
        \pool/pool/pe_b/peij_2_0/add/notb [7]), .Z(
        \pool/pool/pe_b/peij_2_0/add/fai_7/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_7/U3  ( .A(
        \pool/pool/pe_b/peij_2_0/add/cprop [7]), .B(
        \pool/pool/pe_b/peij_2_0/add/fai_7/n3 ), .Z(
        \pool/pool/pe_b/peij_2_0/d_acc [7]) );
  INV_X2 \pool/pool/pe_b/peij_2_0/add/fai_7/U2  ( .A(
        \pool/pool/pe_b/peij_2_0/add/fai_7/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_0/add/cprop [8]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_0/add/fai_7/U1  ( .A1(
        \pool/pool/pe_b/peij_2_0/add/notb [7]), .A2(
        \pool/pool/pe_b_o_data[2][40] ), .B1(
        \pool/pool/pe_b/peij_2_0/add/fai_7/n3 ), .B2(
        \pool/pool/pe_b/peij_2_0/add/cprop [7]), .ZN(
        \pool/pool/pe_b/peij_2_0/add/fai_7/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_8/U4  ( .A(
        \pool/pool/pe_b_o_data[2][41] ), .B(
        \pool/pool/pe_b/peij_2_0/add/notb [8]), .Z(
        \pool/pool/pe_b/peij_2_0/add/fai_8/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_8/U3  ( .A(
        \pool/pool/pe_b/peij_2_0/add/cprop [8]), .B(
        \pool/pool/pe_b/peij_2_0/add/fai_8/n3 ), .Z(
        \pool/pool/pe_b/peij_2_0/d_acc [8]) );
  INV_X2 \pool/pool/pe_b/peij_2_0/add/fai_8/U2  ( .A(
        \pool/pool/pe_b/peij_2_0/add/fai_8/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_0/add/cprop [9]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_0/add/fai_8/U1  ( .A1(
        \pool/pool/pe_b/peij_2_0/add/notb [8]), .A2(
        \pool/pool/pe_b_o_data[2][41] ), .B1(
        \pool/pool/pe_b/peij_2_0/add/fai_8/n3 ), .B2(
        \pool/pool/pe_b/peij_2_0/add/cprop [8]), .ZN(
        \pool/pool/pe_b/peij_2_0/add/fai_8/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_9/U4  ( .A(
        \pool/pool/pe_b_o_data[2][42] ), .B(
        \pool/pool/pe_b/peij_2_0/add/notb [9]), .Z(
        \pool/pool/pe_b/peij_2_0/add/fai_9/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_9/U3  ( .A(
        \pool/pool/pe_b/peij_2_0/add/cprop [9]), .B(
        \pool/pool/pe_b/peij_2_0/add/fai_9/n3 ), .Z(
        \pool/pool/pe_b/peij_2_0/d_acc [9]) );
  INV_X2 \pool/pool/pe_b/peij_2_0/add/fai_9/U2  ( .A(
        \pool/pool/pe_b/peij_2_0/add/fai_9/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_0/add/cprop [10]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_0/add/fai_9/U1  ( .A1(
        \pool/pool/pe_b/peij_2_0/add/notb [9]), .A2(
        \pool/pool/pe_b_o_data[2][42] ), .B1(
        \pool/pool/pe_b/peij_2_0/add/fai_9/n3 ), .B2(
        \pool/pool/pe_b/peij_2_0/add/cprop [9]), .ZN(
        \pool/pool/pe_b/peij_2_0/add/fai_9/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_10/U4  ( .A(
        \pool/pool/pe_b_o_data[2][43] ), .B(
        \pool/pool/pe_b/peij_2_0/add/notb [10]), .Z(
        \pool/pool/pe_b/peij_2_0/add/fai_10/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_0/add/fai_10/U3  ( .A(
        \pool/pool/pe_b/peij_2_0/add/cprop [10]), .B(
        \pool/pool/pe_b/peij_2_0/add/fai_10/n3 ), .Z(
        \pool/pool/pe_b/peij_2_0/d_acc [10]) );
  INV_X2 \pool/pool/pe_b/peij_2_0/add/fai_10/U2  ( .A(
        \pool/pool/pe_b/peij_2_0/add/fai_10/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_0/add/c_out ) );
  AOI22_X2 \pool/pool/pe_b/peij_2_0/add/fai_10/U1  ( .A1(
        \pool/pool/pe_b/peij_2_0/add/notb [10]), .A2(
        \pool/pool/pe_b_o_data[2][43] ), .B1(
        \pool/pool/pe_b/peij_2_0/add/fai_10/n3 ), .B2(
        \pool/pool/pe_b/peij_2_0/add/cprop [10]), .ZN(
        \pool/pool/pe_b/peij_2_0/add/fai_10/n1 ) );
  INV_X1 \pool/pool/pe_b/peij_2_1/U22  ( .A(\pool/pool/pe_b/n6 ), .ZN(
        \pool/pool/pe_b/peij_2_1/n16 ) );
  INV_X1 \pool/pool/pe_b/peij_2_1/U14  ( .A(\pool/pool/pe_b/n6 ), .ZN(
        \pool/pool/pe_b/peij_2_1/n12 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_1/U13  ( .A1(
        \pool/pool/pe_b/peij_2_1/d_acc [0]), .A2(\pool/pool/pe_b/peij_2_1/n18 ), .ZN(\pool/pool/pe_b/peij_2_1/n11 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_1/U12  ( .A1(
        \pool/pool/pe_b/peij_2_1/d_acc [1]), .A2(\pool/pool/pe_b/peij_2_1/n18 ), .ZN(\pool/pool/pe_b/peij_2_1/n10 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_1/U11  ( .A1(
        \pool/pool/pe_b/peij_2_1/d_acc [2]), .A2(\pool/pool/pe_b/peij_2_1/n18 ), .ZN(\pool/pool/pe_b/peij_2_1/n9 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_1/U10  ( .A1(
        \pool/pool/pe_b/peij_2_1/d_acc [3]), .A2(\pool/pool/pe_b/peij_2_1/n18 ), .ZN(\pool/pool/pe_b/peij_2_1/n8 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_1/U9  ( .A1(
        \pool/pool/pe_b/peij_2_1/d_acc [4]), .A2(\pool/pool/pe_b/peij_2_1/n18 ), .ZN(\pool/pool/pe_b/peij_2_1/n7 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_1/U8  ( .A1(
        \pool/pool/pe_b/peij_2_1/d_acc [5]), .A2(\pool/pool/pe_b/peij_2_1/n18 ), .ZN(\pool/pool/pe_b/peij_2_1/n6 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_1/U7  ( .A1(
        \pool/pool/pe_b/peij_2_1/d_acc [6]), .A2(\pool/pool/pe_b/peij_2_1/n18 ), .ZN(\pool/pool/pe_b/peij_2_1/n5 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_1/U6  ( .A1(
        \pool/pool/pe_b/peij_2_1/d_acc [7]), .A2(\pool/pool/pe_b/peij_2_1/n18 ), .ZN(\pool/pool/pe_b/peij_2_1/n4 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_1/U5  ( .A1(
        \pool/pool/pe_b/peij_2_1/d_acc [8]), .A2(\pool/pool/pe_b/peij_2_1/n18 ), .ZN(\pool/pool/pe_b/peij_2_1/n3 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_1/U4  ( .A1(
        \pool/pool/pe_b/peij_2_1/d_acc [9]), .A2(\pool/pool/pe_b/peij_2_1/n18 ), .ZN(\pool/pool/pe_b/peij_2_1/n2 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_1/U3  ( .A1(
        \pool/pool/pe_b/peij_2_1/d_acc [10]), .A2(
        \pool/pool/pe_b/peij_2_1/n18 ), .ZN(\pool/pool/pe_b/peij_2_1/n1 ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_1/q_acc_reg[10]  ( .D(
        \pool/pool/pe_b/peij_2_1/n1 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_1/n16 ), .Q(\pool/pool/pe_b_o_data[2][32] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_1/q_acc_reg[9]  ( .D(
        \pool/pool/pe_b/peij_2_1/n2 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_1/n16 ), .Q(\pool/pool/pe_b_o_data[2][31] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_1/q_acc_reg[8]  ( .D(
        \pool/pool/pe_b/peij_2_1/n3 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_1/n16 ), .Q(\pool/pool/pe_b_o_data[2][30] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_1/q_acc_reg[7]  ( .D(
        \pool/pool/pe_b/peij_2_1/n4 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_1/n16 ), .Q(\pool/pool/pe_b_o_data[2][29] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_1/q_acc_reg[6]  ( .D(
        \pool/pool/pe_b/peij_2_1/n5 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_1/n16 ), .Q(\pool/pool/pe_b_o_data[2][28] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_1/q_acc_reg[5]  ( .D(
        \pool/pool/pe_b/peij_2_1/n6 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_1/n16 ), .Q(\pool/pool/pe_b_o_data[2][27] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_1/q_acc_reg[4]  ( .D(
        \pool/pool/pe_b/peij_2_1/n7 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_1/n16 ), .Q(\pool/pool/pe_b_o_data[2][26] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_1/q_acc_reg[3]  ( .D(
        \pool/pool/pe_b/peij_2_1/n8 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_1/n16 ), .Q(\pool/pool/pe_b_o_data[2][25] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_1/q_acc_reg[2]  ( .D(
        \pool/pool/pe_b/peij_2_1/n9 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_1/n16 ), .Q(\pool/pool/pe_b_o_data[2][24] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_1/q_acc_reg[1]  ( .D(
        \pool/pool/pe_b/peij_2_1/n10 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_1/n16 ), .Q(\pool/pool/pe_b_o_data[2][23] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_1/q_acc_reg[0]  ( .D(
        \pool/pool/pe_b/peij_2_1/n11 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_1/n16 ), .Q(\pool/pool/pe_b_o_data[2][22] ) );
  INV_X2 \pool/pool/pe_b/peij_2_1/U21  ( .A(\pool/sync_clr ), .ZN(
        \pool/pool/pe_b/peij_2_1/n18 ) );
  AND3_X2 \pool/pool/pe_b/peij_2_1/U20  ( .A1(\pool/pool/pe_b/int_pe_en[2][1] ), .A2(\pool/pool/pe_b/peij_2_1/n18 ), .A3(1'b1), .ZN(
        \pool/pool/pe_b/peij_2_1/n17 ) );
  AND2_X2 \pool/pool/pe_b/peij_2_1/U19  ( .A1(\pool/pool/pe_b_i_data[2][8] ), 
        .A2(\pool/pool/pe_b/peij_2_1/n17 ), .ZN(\pool/pool/pe_b/peij_2_1/N33 )
         );
  AND2_X2 \pool/pool/pe_b/peij_2_1/U18  ( .A1(\pool/pool/pe_b_i_data[2][9] ), 
        .A2(\pool/pool/pe_b/peij_2_1/n17 ), .ZN(\pool/pool/pe_b/peij_2_1/N34 )
         );
  AND2_X2 \pool/pool/pe_b/peij_2_1/U17  ( .A1(\pool/pool/pe_b_i_data[2][10] ), 
        .A2(\pool/pool/pe_b/peij_2_1/n17 ), .ZN(\pool/pool/pe_b/peij_2_1/N35 )
         );
  AND4_X4 \pool/pool/pe_b/peij_2_1/U16  ( .A1(1'b1), .A2(
        \pool/pool/pe_b_i_data[2][11] ), .A3(\pool/pool/pe_b/int_pe_en[2][1] ), 
        .A4(\pool/pool/pe_b/peij_2_1/n18 ), .ZN(\pool/pool/pe_b/peij_2_1/N36 )
         );
  DFFR_X1 \pool/pool/pe_b/peij_2_1/q_im_reg[0]  ( .D(
        \pool/pool/pe_b/peij_2_1/N33 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_1/n12 ), .Q(\pool/pool/pe_b/peij_2_1/sgnext [0]) );
  DFFR_X1 \pool/pool/pe_b/peij_2_1/q_im_reg[1]  ( .D(
        \pool/pool/pe_b/peij_2_1/N34 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_1/n12 ), .Q(\pool/pool/pe_b/peij_2_1/sgnext [1]) );
  DFFR_X1 \pool/pool/pe_b/peij_2_1/q_im_reg[2]  ( .D(
        \pool/pool/pe_b/peij_2_1/N35 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_1/n12 ), .Q(\pool/pool/pe_b/peij_2_1/sgnext [2]) );
  DFFR_X1 \pool/pool/pe_b/peij_2_1/q_im_reg[3]  ( .D(
        \pool/pool/pe_b/peij_2_1/N36 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_1/n12 ), .Q(\pool/pool/pe_b/peij_2_1/sgnext_10 ) );
  SDFFR_X1 \pool/pool/pe_b/peij_2_1/q_k_reg  ( .D(1'b0), .SI(
        \pool/pool/pe_b/peij_2_1/n18 ), .SE(1'b0), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_1/n12 ), .Q(\pool/pool/pe_b/peij_2_1/q_k ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/U11  ( .A(
        \pool/pool/pe_b/peij_2_1/sgnext [0]), .B(\pool/pool/pe_b/peij_2_1/q_k ), .Z(\pool/pool/pe_b/peij_2_1/add/notb [0]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/U10  ( .A(
        \pool/pool/pe_b/peij_2_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_1/q_k ), .Z(\pool/pool/pe_b/peij_2_1/add/notb [10]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/U9  ( .A(
        \pool/pool/pe_b/peij_2_1/sgnext [1]), .B(\pool/pool/pe_b/peij_2_1/q_k ), .Z(\pool/pool/pe_b/peij_2_1/add/notb [1]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/U8  ( .A(
        \pool/pool/pe_b/peij_2_1/sgnext [2]), .B(\pool/pool/pe_b/peij_2_1/q_k ), .Z(\pool/pool/pe_b/peij_2_1/add/notb [2]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/U7  ( .A(
        \pool/pool/pe_b/peij_2_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_1/q_k ), .Z(\pool/pool/pe_b/peij_2_1/add/notb [3]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/U6  ( .A(
        \pool/pool/pe_b/peij_2_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_1/q_k ), .Z(\pool/pool/pe_b/peij_2_1/add/notb [4]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/U5  ( .A(
        \pool/pool/pe_b/peij_2_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_1/q_k ), .Z(\pool/pool/pe_b/peij_2_1/add/notb [5]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/U4  ( .A(
        \pool/pool/pe_b/peij_2_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_1/q_k ), .Z(\pool/pool/pe_b/peij_2_1/add/notb [6]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/U3  ( .A(
        \pool/pool/pe_b/peij_2_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_1/q_k ), .Z(\pool/pool/pe_b/peij_2_1/add/notb [7]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/U2  ( .A(
        \pool/pool/pe_b/peij_2_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_1/q_k ), .Z(\pool/pool/pe_b/peij_2_1/add/notb [8]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/U1  ( .A(
        \pool/pool/pe_b/peij_2_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_1/q_k ), .Z(\pool/pool/pe_b/peij_2_1/add/notb [9]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_0/U4  ( .A(
        \pool/pool/pe_b_o_data[2][22] ), .B(
        \pool/pool/pe_b/peij_2_1/add/notb [0]), .Z(
        \pool/pool/pe_b/peij_2_1/add/fai_0/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_0/U3  ( .A(
        \pool/pool/pe_b/peij_2_1/q_k ), .B(
        \pool/pool/pe_b/peij_2_1/add/fai_0/n3 ), .Z(
        \pool/pool/pe_b/peij_2_1/d_acc [0]) );
  INV_X2 \pool/pool/pe_b/peij_2_1/add/fai_0/U2  ( .A(
        \pool/pool/pe_b/peij_2_1/add/fai_0/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_1/add/cprop [1]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_1/add/fai_0/U1  ( .A1(
        \pool/pool/pe_b/peij_2_1/add/notb [0]), .A2(
        \pool/pool/pe_b_o_data[2][22] ), .B1(
        \pool/pool/pe_b/peij_2_1/add/fai_0/n3 ), .B2(
        \pool/pool/pe_b/peij_2_1/q_k ), .ZN(
        \pool/pool/pe_b/peij_2_1/add/fai_0/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_1/U4  ( .A(
        \pool/pool/pe_b_o_data[2][23] ), .B(
        \pool/pool/pe_b/peij_2_1/add/notb [1]), .Z(
        \pool/pool/pe_b/peij_2_1/add/fai_1/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_1/U3  ( .A(
        \pool/pool/pe_b/peij_2_1/add/cprop [1]), .B(
        \pool/pool/pe_b/peij_2_1/add/fai_1/n3 ), .Z(
        \pool/pool/pe_b/peij_2_1/d_acc [1]) );
  INV_X2 \pool/pool/pe_b/peij_2_1/add/fai_1/U2  ( .A(
        \pool/pool/pe_b/peij_2_1/add/fai_1/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_1/add/cprop [2]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_1/add/fai_1/U1  ( .A1(
        \pool/pool/pe_b/peij_2_1/add/notb [1]), .A2(
        \pool/pool/pe_b_o_data[2][23] ), .B1(
        \pool/pool/pe_b/peij_2_1/add/fai_1/n3 ), .B2(
        \pool/pool/pe_b/peij_2_1/add/cprop [1]), .ZN(
        \pool/pool/pe_b/peij_2_1/add/fai_1/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_2/U4  ( .A(
        \pool/pool/pe_b_o_data[2][24] ), .B(
        \pool/pool/pe_b/peij_2_1/add/notb [2]), .Z(
        \pool/pool/pe_b/peij_2_1/add/fai_2/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_2/U3  ( .A(
        \pool/pool/pe_b/peij_2_1/add/cprop [2]), .B(
        \pool/pool/pe_b/peij_2_1/add/fai_2/n3 ), .Z(
        \pool/pool/pe_b/peij_2_1/d_acc [2]) );
  INV_X2 \pool/pool/pe_b/peij_2_1/add/fai_2/U2  ( .A(
        \pool/pool/pe_b/peij_2_1/add/fai_2/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_1/add/cprop [3]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_1/add/fai_2/U1  ( .A1(
        \pool/pool/pe_b/peij_2_1/add/notb [2]), .A2(
        \pool/pool/pe_b_o_data[2][24] ), .B1(
        \pool/pool/pe_b/peij_2_1/add/fai_2/n3 ), .B2(
        \pool/pool/pe_b/peij_2_1/add/cprop [2]), .ZN(
        \pool/pool/pe_b/peij_2_1/add/fai_2/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_3/U4  ( .A(
        \pool/pool/pe_b_o_data[2][25] ), .B(
        \pool/pool/pe_b/peij_2_1/add/notb [3]), .Z(
        \pool/pool/pe_b/peij_2_1/add/fai_3/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_3/U3  ( .A(
        \pool/pool/pe_b/peij_2_1/add/cprop [3]), .B(
        \pool/pool/pe_b/peij_2_1/add/fai_3/n3 ), .Z(
        \pool/pool/pe_b/peij_2_1/d_acc [3]) );
  INV_X2 \pool/pool/pe_b/peij_2_1/add/fai_3/U2  ( .A(
        \pool/pool/pe_b/peij_2_1/add/fai_3/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_1/add/cprop [4]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_1/add/fai_3/U1  ( .A1(
        \pool/pool/pe_b/peij_2_1/add/notb [3]), .A2(
        \pool/pool/pe_b_o_data[2][25] ), .B1(
        \pool/pool/pe_b/peij_2_1/add/fai_3/n3 ), .B2(
        \pool/pool/pe_b/peij_2_1/add/cprop [3]), .ZN(
        \pool/pool/pe_b/peij_2_1/add/fai_3/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_4/U4  ( .A(
        \pool/pool/pe_b_o_data[2][26] ), .B(
        \pool/pool/pe_b/peij_2_1/add/notb [4]), .Z(
        \pool/pool/pe_b/peij_2_1/add/fai_4/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_4/U3  ( .A(
        \pool/pool/pe_b/peij_2_1/add/cprop [4]), .B(
        \pool/pool/pe_b/peij_2_1/add/fai_4/n3 ), .Z(
        \pool/pool/pe_b/peij_2_1/d_acc [4]) );
  INV_X2 \pool/pool/pe_b/peij_2_1/add/fai_4/U2  ( .A(
        \pool/pool/pe_b/peij_2_1/add/fai_4/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_1/add/cprop [5]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_1/add/fai_4/U1  ( .A1(
        \pool/pool/pe_b/peij_2_1/add/notb [4]), .A2(
        \pool/pool/pe_b_o_data[2][26] ), .B1(
        \pool/pool/pe_b/peij_2_1/add/fai_4/n3 ), .B2(
        \pool/pool/pe_b/peij_2_1/add/cprop [4]), .ZN(
        \pool/pool/pe_b/peij_2_1/add/fai_4/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_5/U4  ( .A(
        \pool/pool/pe_b_o_data[2][27] ), .B(
        \pool/pool/pe_b/peij_2_1/add/notb [5]), .Z(
        \pool/pool/pe_b/peij_2_1/add/fai_5/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_5/U3  ( .A(
        \pool/pool/pe_b/peij_2_1/add/cprop [5]), .B(
        \pool/pool/pe_b/peij_2_1/add/fai_5/n3 ), .Z(
        \pool/pool/pe_b/peij_2_1/d_acc [5]) );
  INV_X2 \pool/pool/pe_b/peij_2_1/add/fai_5/U2  ( .A(
        \pool/pool/pe_b/peij_2_1/add/fai_5/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_1/add/cprop [6]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_1/add/fai_5/U1  ( .A1(
        \pool/pool/pe_b/peij_2_1/add/notb [5]), .A2(
        \pool/pool/pe_b_o_data[2][27] ), .B1(
        \pool/pool/pe_b/peij_2_1/add/fai_5/n3 ), .B2(
        \pool/pool/pe_b/peij_2_1/add/cprop [5]), .ZN(
        \pool/pool/pe_b/peij_2_1/add/fai_5/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_6/U4  ( .A(
        \pool/pool/pe_b_o_data[2][28] ), .B(
        \pool/pool/pe_b/peij_2_1/add/notb [6]), .Z(
        \pool/pool/pe_b/peij_2_1/add/fai_6/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_6/U3  ( .A(
        \pool/pool/pe_b/peij_2_1/add/cprop [6]), .B(
        \pool/pool/pe_b/peij_2_1/add/fai_6/n3 ), .Z(
        \pool/pool/pe_b/peij_2_1/d_acc [6]) );
  INV_X2 \pool/pool/pe_b/peij_2_1/add/fai_6/U2  ( .A(
        \pool/pool/pe_b/peij_2_1/add/fai_6/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_1/add/cprop [7]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_1/add/fai_6/U1  ( .A1(
        \pool/pool/pe_b/peij_2_1/add/notb [6]), .A2(
        \pool/pool/pe_b_o_data[2][28] ), .B1(
        \pool/pool/pe_b/peij_2_1/add/fai_6/n3 ), .B2(
        \pool/pool/pe_b/peij_2_1/add/cprop [6]), .ZN(
        \pool/pool/pe_b/peij_2_1/add/fai_6/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_7/U4  ( .A(
        \pool/pool/pe_b_o_data[2][29] ), .B(
        \pool/pool/pe_b/peij_2_1/add/notb [7]), .Z(
        \pool/pool/pe_b/peij_2_1/add/fai_7/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_7/U3  ( .A(
        \pool/pool/pe_b/peij_2_1/add/cprop [7]), .B(
        \pool/pool/pe_b/peij_2_1/add/fai_7/n3 ), .Z(
        \pool/pool/pe_b/peij_2_1/d_acc [7]) );
  INV_X2 \pool/pool/pe_b/peij_2_1/add/fai_7/U2  ( .A(
        \pool/pool/pe_b/peij_2_1/add/fai_7/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_1/add/cprop [8]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_1/add/fai_7/U1  ( .A1(
        \pool/pool/pe_b/peij_2_1/add/notb [7]), .A2(
        \pool/pool/pe_b_o_data[2][29] ), .B1(
        \pool/pool/pe_b/peij_2_1/add/fai_7/n3 ), .B2(
        \pool/pool/pe_b/peij_2_1/add/cprop [7]), .ZN(
        \pool/pool/pe_b/peij_2_1/add/fai_7/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_8/U4  ( .A(
        \pool/pool/pe_b_o_data[2][30] ), .B(
        \pool/pool/pe_b/peij_2_1/add/notb [8]), .Z(
        \pool/pool/pe_b/peij_2_1/add/fai_8/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_8/U3  ( .A(
        \pool/pool/pe_b/peij_2_1/add/cprop [8]), .B(
        \pool/pool/pe_b/peij_2_1/add/fai_8/n3 ), .Z(
        \pool/pool/pe_b/peij_2_1/d_acc [8]) );
  INV_X2 \pool/pool/pe_b/peij_2_1/add/fai_8/U2  ( .A(
        \pool/pool/pe_b/peij_2_1/add/fai_8/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_1/add/cprop [9]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_1/add/fai_8/U1  ( .A1(
        \pool/pool/pe_b/peij_2_1/add/notb [8]), .A2(
        \pool/pool/pe_b_o_data[2][30] ), .B1(
        \pool/pool/pe_b/peij_2_1/add/fai_8/n3 ), .B2(
        \pool/pool/pe_b/peij_2_1/add/cprop [8]), .ZN(
        \pool/pool/pe_b/peij_2_1/add/fai_8/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_9/U4  ( .A(
        \pool/pool/pe_b_o_data[2][31] ), .B(
        \pool/pool/pe_b/peij_2_1/add/notb [9]), .Z(
        \pool/pool/pe_b/peij_2_1/add/fai_9/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_9/U3  ( .A(
        \pool/pool/pe_b/peij_2_1/add/cprop [9]), .B(
        \pool/pool/pe_b/peij_2_1/add/fai_9/n3 ), .Z(
        \pool/pool/pe_b/peij_2_1/d_acc [9]) );
  INV_X2 \pool/pool/pe_b/peij_2_1/add/fai_9/U2  ( .A(
        \pool/pool/pe_b/peij_2_1/add/fai_9/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_1/add/cprop [10]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_1/add/fai_9/U1  ( .A1(
        \pool/pool/pe_b/peij_2_1/add/notb [9]), .A2(
        \pool/pool/pe_b_o_data[2][31] ), .B1(
        \pool/pool/pe_b/peij_2_1/add/fai_9/n3 ), .B2(
        \pool/pool/pe_b/peij_2_1/add/cprop [9]), .ZN(
        \pool/pool/pe_b/peij_2_1/add/fai_9/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_10/U4  ( .A(
        \pool/pool/pe_b_o_data[2][32] ), .B(
        \pool/pool/pe_b/peij_2_1/add/notb [10]), .Z(
        \pool/pool/pe_b/peij_2_1/add/fai_10/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_1/add/fai_10/U3  ( .A(
        \pool/pool/pe_b/peij_2_1/add/cprop [10]), .B(
        \pool/pool/pe_b/peij_2_1/add/fai_10/n3 ), .Z(
        \pool/pool/pe_b/peij_2_1/d_acc [10]) );
  INV_X2 \pool/pool/pe_b/peij_2_1/add/fai_10/U2  ( .A(
        \pool/pool/pe_b/peij_2_1/add/fai_10/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_1/add/c_out ) );
  AOI22_X2 \pool/pool/pe_b/peij_2_1/add/fai_10/U1  ( .A1(
        \pool/pool/pe_b/peij_2_1/add/notb [10]), .A2(
        \pool/pool/pe_b_o_data[2][32] ), .B1(
        \pool/pool/pe_b/peij_2_1/add/fai_10/n3 ), .B2(
        \pool/pool/pe_b/peij_2_1/add/cprop [10]), .ZN(
        \pool/pool/pe_b/peij_2_1/add/fai_10/n1 ) );
  INV_X1 \pool/pool/pe_b/peij_2_2/U22  ( .A(\pool/pool/pe_b/n7 ), .ZN(
        \pool/pool/pe_b/peij_2_2/n16 ) );
  INV_X1 \pool/pool/pe_b/peij_2_2/U14  ( .A(\pool/pool/pe_b/n7 ), .ZN(
        \pool/pool/pe_b/peij_2_2/n12 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_2/U13  ( .A1(
        \pool/pool/pe_b/peij_2_2/d_acc [0]), .A2(\pool/pool/pe_b/peij_2_2/n18 ), .ZN(\pool/pool/pe_b/peij_2_2/n11 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_2/U12  ( .A1(
        \pool/pool/pe_b/peij_2_2/d_acc [1]), .A2(\pool/pool/pe_b/peij_2_2/n18 ), .ZN(\pool/pool/pe_b/peij_2_2/n10 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_2/U11  ( .A1(
        \pool/pool/pe_b/peij_2_2/d_acc [2]), .A2(\pool/pool/pe_b/peij_2_2/n18 ), .ZN(\pool/pool/pe_b/peij_2_2/n9 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_2/U10  ( .A1(
        \pool/pool/pe_b/peij_2_2/d_acc [3]), .A2(\pool/pool/pe_b/peij_2_2/n18 ), .ZN(\pool/pool/pe_b/peij_2_2/n8 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_2/U9  ( .A1(
        \pool/pool/pe_b/peij_2_2/d_acc [4]), .A2(\pool/pool/pe_b/peij_2_2/n18 ), .ZN(\pool/pool/pe_b/peij_2_2/n7 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_2/U8  ( .A1(
        \pool/pool/pe_b/peij_2_2/d_acc [5]), .A2(\pool/pool/pe_b/peij_2_2/n18 ), .ZN(\pool/pool/pe_b/peij_2_2/n6 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_2/U7  ( .A1(
        \pool/pool/pe_b/peij_2_2/d_acc [6]), .A2(\pool/pool/pe_b/peij_2_2/n18 ), .ZN(\pool/pool/pe_b/peij_2_2/n5 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_2/U6  ( .A1(
        \pool/pool/pe_b/peij_2_2/d_acc [7]), .A2(\pool/pool/pe_b/peij_2_2/n18 ), .ZN(\pool/pool/pe_b/peij_2_2/n4 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_2/U5  ( .A1(
        \pool/pool/pe_b/peij_2_2/d_acc [8]), .A2(\pool/pool/pe_b/peij_2_2/n18 ), .ZN(\pool/pool/pe_b/peij_2_2/n3 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_2/U4  ( .A1(
        \pool/pool/pe_b/peij_2_2/d_acc [9]), .A2(\pool/pool/pe_b/peij_2_2/n18 ), .ZN(\pool/pool/pe_b/peij_2_2/n2 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_2/U3  ( .A1(
        \pool/pool/pe_b/peij_2_2/d_acc [10]), .A2(
        \pool/pool/pe_b/peij_2_2/n18 ), .ZN(\pool/pool/pe_b/peij_2_2/n1 ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_2/q_acc_reg[10]  ( .D(
        \pool/pool/pe_b/peij_2_2/n1 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_2/n16 ), .Q(\pool/pool/pe_b_o_data[2][21] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_2/q_acc_reg[9]  ( .D(
        \pool/pool/pe_b/peij_2_2/n2 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_2/n16 ), .Q(\pool/pool/pe_b_o_data[2][20] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_2/q_acc_reg[8]  ( .D(
        \pool/pool/pe_b/peij_2_2/n3 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_2/n16 ), .Q(\pool/pool/pe_b_o_data[2][19] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_2/q_acc_reg[7]  ( .D(
        \pool/pool/pe_b/peij_2_2/n4 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_2/n16 ), .Q(\pool/pool/pe_b_o_data[2][18] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_2/q_acc_reg[6]  ( .D(
        \pool/pool/pe_b/peij_2_2/n5 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_2/n16 ), .Q(\pool/pool/pe_b_o_data[2][17] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_2/q_acc_reg[5]  ( .D(
        \pool/pool/pe_b/peij_2_2/n6 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_2/n16 ), .Q(\pool/pool/pe_b_o_data[2][16] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_2/q_acc_reg[4]  ( .D(
        \pool/pool/pe_b/peij_2_2/n7 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_2/n16 ), .Q(\pool/pool/pe_b_o_data[2][15] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_2/q_acc_reg[3]  ( .D(
        \pool/pool/pe_b/peij_2_2/n8 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_2/n16 ), .Q(\pool/pool/pe_b_o_data[2][14] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_2/q_acc_reg[2]  ( .D(
        \pool/pool/pe_b/peij_2_2/n9 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_2/n16 ), .Q(\pool/pool/pe_b_o_data[2][13] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_2/q_acc_reg[1]  ( .D(
        \pool/pool/pe_b/peij_2_2/n10 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_2/n16 ), .Q(\pool/pool/pe_b_o_data[2][12] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_2/q_acc_reg[0]  ( .D(
        \pool/pool/pe_b/peij_2_2/n11 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_2/n16 ), .Q(\pool/pool/pe_b_o_data[2][11] ) );
  INV_X2 \pool/pool/pe_b/peij_2_2/U21  ( .A(\pool/sync_clr ), .ZN(
        \pool/pool/pe_b/peij_2_2/n18 ) );
  AND3_X2 \pool/pool/pe_b/peij_2_2/U20  ( .A1(\pool/pool/pe_b/int_pe_en[2][2] ), .A2(\pool/pool/pe_b/peij_2_2/n18 ), .A3(1'b1), .ZN(
        \pool/pool/pe_b/peij_2_2/n17 ) );
  AND2_X2 \pool/pool/pe_b/peij_2_2/U19  ( .A1(\pool/pool/pe_b_i_data[2][4] ), 
        .A2(\pool/pool/pe_b/peij_2_2/n17 ), .ZN(\pool/pool/pe_b/peij_2_2/N33 )
         );
  AND2_X2 \pool/pool/pe_b/peij_2_2/U18  ( .A1(\pool/pool/pe_b_i_data[2][5] ), 
        .A2(\pool/pool/pe_b/peij_2_2/n17 ), .ZN(\pool/pool/pe_b/peij_2_2/N34 )
         );
  AND2_X2 \pool/pool/pe_b/peij_2_2/U17  ( .A1(\pool/pool/pe_b_i_data[2][6] ), 
        .A2(\pool/pool/pe_b/peij_2_2/n17 ), .ZN(\pool/pool/pe_b/peij_2_2/N35 )
         );
  AND4_X4 \pool/pool/pe_b/peij_2_2/U16  ( .A1(1'b1), .A2(
        \pool/pool/pe_b_i_data[2][7] ), .A3(\pool/pool/pe_b/int_pe_en[2][2] ), 
        .A4(\pool/pool/pe_b/peij_2_2/n18 ), .ZN(\pool/pool/pe_b/peij_2_2/N36 )
         );
  DFFR_X1 \pool/pool/pe_b/peij_2_2/q_im_reg[0]  ( .D(
        \pool/pool/pe_b/peij_2_2/N33 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_2/n12 ), .Q(\pool/pool/pe_b/peij_2_2/sgnext [0]) );
  DFFR_X1 \pool/pool/pe_b/peij_2_2/q_im_reg[1]  ( .D(
        \pool/pool/pe_b/peij_2_2/N34 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_2/n12 ), .Q(\pool/pool/pe_b/peij_2_2/sgnext [1]) );
  DFFR_X1 \pool/pool/pe_b/peij_2_2/q_im_reg[2]  ( .D(
        \pool/pool/pe_b/peij_2_2/N35 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_2/n12 ), .Q(\pool/pool/pe_b/peij_2_2/sgnext [2]) );
  DFFR_X1 \pool/pool/pe_b/peij_2_2/q_im_reg[3]  ( .D(
        \pool/pool/pe_b/peij_2_2/N36 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_2/n12 ), .Q(\pool/pool/pe_b/peij_2_2/sgnext_10 ) );
  SDFFR_X1 \pool/pool/pe_b/peij_2_2/q_k_reg  ( .D(1'b0), .SI(
        \pool/pool/pe_b/peij_2_2/n18 ), .SE(1'b0), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_2/n12 ), .Q(\pool/pool/pe_b/peij_2_2/q_k ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/U11  ( .A(
        \pool/pool/pe_b/peij_2_2/sgnext [0]), .B(\pool/pool/pe_b/peij_2_2/q_k ), .Z(\pool/pool/pe_b/peij_2_2/add/notb [0]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/U10  ( .A(
        \pool/pool/pe_b/peij_2_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_2/q_k ), .Z(\pool/pool/pe_b/peij_2_2/add/notb [10]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/U9  ( .A(
        \pool/pool/pe_b/peij_2_2/sgnext [1]), .B(\pool/pool/pe_b/peij_2_2/q_k ), .Z(\pool/pool/pe_b/peij_2_2/add/notb [1]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/U8  ( .A(
        \pool/pool/pe_b/peij_2_2/sgnext [2]), .B(\pool/pool/pe_b/peij_2_2/q_k ), .Z(\pool/pool/pe_b/peij_2_2/add/notb [2]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/U7  ( .A(
        \pool/pool/pe_b/peij_2_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_2/q_k ), .Z(\pool/pool/pe_b/peij_2_2/add/notb [3]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/U6  ( .A(
        \pool/pool/pe_b/peij_2_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_2/q_k ), .Z(\pool/pool/pe_b/peij_2_2/add/notb [4]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/U5  ( .A(
        \pool/pool/pe_b/peij_2_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_2/q_k ), .Z(\pool/pool/pe_b/peij_2_2/add/notb [5]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/U4  ( .A(
        \pool/pool/pe_b/peij_2_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_2/q_k ), .Z(\pool/pool/pe_b/peij_2_2/add/notb [6]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/U3  ( .A(
        \pool/pool/pe_b/peij_2_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_2/q_k ), .Z(\pool/pool/pe_b/peij_2_2/add/notb [7]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/U2  ( .A(
        \pool/pool/pe_b/peij_2_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_2/q_k ), .Z(\pool/pool/pe_b/peij_2_2/add/notb [8]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/U1  ( .A(
        \pool/pool/pe_b/peij_2_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_2/q_k ), .Z(\pool/pool/pe_b/peij_2_2/add/notb [9]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_0/U4  ( .A(
        \pool/pool/pe_b_o_data[2][11] ), .B(
        \pool/pool/pe_b/peij_2_2/add/notb [0]), .Z(
        \pool/pool/pe_b/peij_2_2/add/fai_0/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_0/U3  ( .A(
        \pool/pool/pe_b/peij_2_2/q_k ), .B(
        \pool/pool/pe_b/peij_2_2/add/fai_0/n3 ), .Z(
        \pool/pool/pe_b/peij_2_2/d_acc [0]) );
  INV_X2 \pool/pool/pe_b/peij_2_2/add/fai_0/U2  ( .A(
        \pool/pool/pe_b/peij_2_2/add/fai_0/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_2/add/cprop [1]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_2/add/fai_0/U1  ( .A1(
        \pool/pool/pe_b/peij_2_2/add/notb [0]), .A2(
        \pool/pool/pe_b_o_data[2][11] ), .B1(
        \pool/pool/pe_b/peij_2_2/add/fai_0/n3 ), .B2(
        \pool/pool/pe_b/peij_2_2/q_k ), .ZN(
        \pool/pool/pe_b/peij_2_2/add/fai_0/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_1/U4  ( .A(
        \pool/pool/pe_b_o_data[2][12] ), .B(
        \pool/pool/pe_b/peij_2_2/add/notb [1]), .Z(
        \pool/pool/pe_b/peij_2_2/add/fai_1/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_1/U3  ( .A(
        \pool/pool/pe_b/peij_2_2/add/cprop [1]), .B(
        \pool/pool/pe_b/peij_2_2/add/fai_1/n3 ), .Z(
        \pool/pool/pe_b/peij_2_2/d_acc [1]) );
  INV_X2 \pool/pool/pe_b/peij_2_2/add/fai_1/U2  ( .A(
        \pool/pool/pe_b/peij_2_2/add/fai_1/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_2/add/cprop [2]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_2/add/fai_1/U1  ( .A1(
        \pool/pool/pe_b/peij_2_2/add/notb [1]), .A2(
        \pool/pool/pe_b_o_data[2][12] ), .B1(
        \pool/pool/pe_b/peij_2_2/add/fai_1/n3 ), .B2(
        \pool/pool/pe_b/peij_2_2/add/cprop [1]), .ZN(
        \pool/pool/pe_b/peij_2_2/add/fai_1/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_2/U4  ( .A(
        \pool/pool/pe_b_o_data[2][13] ), .B(
        \pool/pool/pe_b/peij_2_2/add/notb [2]), .Z(
        \pool/pool/pe_b/peij_2_2/add/fai_2/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_2/U3  ( .A(
        \pool/pool/pe_b/peij_2_2/add/cprop [2]), .B(
        \pool/pool/pe_b/peij_2_2/add/fai_2/n3 ), .Z(
        \pool/pool/pe_b/peij_2_2/d_acc [2]) );
  INV_X2 \pool/pool/pe_b/peij_2_2/add/fai_2/U2  ( .A(
        \pool/pool/pe_b/peij_2_2/add/fai_2/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_2/add/cprop [3]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_2/add/fai_2/U1  ( .A1(
        \pool/pool/pe_b/peij_2_2/add/notb [2]), .A2(
        \pool/pool/pe_b_o_data[2][13] ), .B1(
        \pool/pool/pe_b/peij_2_2/add/fai_2/n3 ), .B2(
        \pool/pool/pe_b/peij_2_2/add/cprop [2]), .ZN(
        \pool/pool/pe_b/peij_2_2/add/fai_2/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_3/U4  ( .A(
        \pool/pool/pe_b_o_data[2][14] ), .B(
        \pool/pool/pe_b/peij_2_2/add/notb [3]), .Z(
        \pool/pool/pe_b/peij_2_2/add/fai_3/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_3/U3  ( .A(
        \pool/pool/pe_b/peij_2_2/add/cprop [3]), .B(
        \pool/pool/pe_b/peij_2_2/add/fai_3/n3 ), .Z(
        \pool/pool/pe_b/peij_2_2/d_acc [3]) );
  INV_X2 \pool/pool/pe_b/peij_2_2/add/fai_3/U2  ( .A(
        \pool/pool/pe_b/peij_2_2/add/fai_3/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_2/add/cprop [4]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_2/add/fai_3/U1  ( .A1(
        \pool/pool/pe_b/peij_2_2/add/notb [3]), .A2(
        \pool/pool/pe_b_o_data[2][14] ), .B1(
        \pool/pool/pe_b/peij_2_2/add/fai_3/n3 ), .B2(
        \pool/pool/pe_b/peij_2_2/add/cprop [3]), .ZN(
        \pool/pool/pe_b/peij_2_2/add/fai_3/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_4/U4  ( .A(
        \pool/pool/pe_b_o_data[2][15] ), .B(
        \pool/pool/pe_b/peij_2_2/add/notb [4]), .Z(
        \pool/pool/pe_b/peij_2_2/add/fai_4/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_4/U3  ( .A(
        \pool/pool/pe_b/peij_2_2/add/cprop [4]), .B(
        \pool/pool/pe_b/peij_2_2/add/fai_4/n3 ), .Z(
        \pool/pool/pe_b/peij_2_2/d_acc [4]) );
  INV_X2 \pool/pool/pe_b/peij_2_2/add/fai_4/U2  ( .A(
        \pool/pool/pe_b/peij_2_2/add/fai_4/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_2/add/cprop [5]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_2/add/fai_4/U1  ( .A1(
        \pool/pool/pe_b/peij_2_2/add/notb [4]), .A2(
        \pool/pool/pe_b_o_data[2][15] ), .B1(
        \pool/pool/pe_b/peij_2_2/add/fai_4/n3 ), .B2(
        \pool/pool/pe_b/peij_2_2/add/cprop [4]), .ZN(
        \pool/pool/pe_b/peij_2_2/add/fai_4/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_5/U4  ( .A(
        \pool/pool/pe_b_o_data[2][16] ), .B(
        \pool/pool/pe_b/peij_2_2/add/notb [5]), .Z(
        \pool/pool/pe_b/peij_2_2/add/fai_5/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_5/U3  ( .A(
        \pool/pool/pe_b/peij_2_2/add/cprop [5]), .B(
        \pool/pool/pe_b/peij_2_2/add/fai_5/n3 ), .Z(
        \pool/pool/pe_b/peij_2_2/d_acc [5]) );
  INV_X2 \pool/pool/pe_b/peij_2_2/add/fai_5/U2  ( .A(
        \pool/pool/pe_b/peij_2_2/add/fai_5/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_2/add/cprop [6]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_2/add/fai_5/U1  ( .A1(
        \pool/pool/pe_b/peij_2_2/add/notb [5]), .A2(
        \pool/pool/pe_b_o_data[2][16] ), .B1(
        \pool/pool/pe_b/peij_2_2/add/fai_5/n3 ), .B2(
        \pool/pool/pe_b/peij_2_2/add/cprop [5]), .ZN(
        \pool/pool/pe_b/peij_2_2/add/fai_5/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_6/U4  ( .A(
        \pool/pool/pe_b_o_data[2][17] ), .B(
        \pool/pool/pe_b/peij_2_2/add/notb [6]), .Z(
        \pool/pool/pe_b/peij_2_2/add/fai_6/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_6/U3  ( .A(
        \pool/pool/pe_b/peij_2_2/add/cprop [6]), .B(
        \pool/pool/pe_b/peij_2_2/add/fai_6/n3 ), .Z(
        \pool/pool/pe_b/peij_2_2/d_acc [6]) );
  INV_X2 \pool/pool/pe_b/peij_2_2/add/fai_6/U2  ( .A(
        \pool/pool/pe_b/peij_2_2/add/fai_6/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_2/add/cprop [7]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_2/add/fai_6/U1  ( .A1(
        \pool/pool/pe_b/peij_2_2/add/notb [6]), .A2(
        \pool/pool/pe_b_o_data[2][17] ), .B1(
        \pool/pool/pe_b/peij_2_2/add/fai_6/n3 ), .B2(
        \pool/pool/pe_b/peij_2_2/add/cprop [6]), .ZN(
        \pool/pool/pe_b/peij_2_2/add/fai_6/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_7/U4  ( .A(
        \pool/pool/pe_b_o_data[2][18] ), .B(
        \pool/pool/pe_b/peij_2_2/add/notb [7]), .Z(
        \pool/pool/pe_b/peij_2_2/add/fai_7/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_7/U3  ( .A(
        \pool/pool/pe_b/peij_2_2/add/cprop [7]), .B(
        \pool/pool/pe_b/peij_2_2/add/fai_7/n3 ), .Z(
        \pool/pool/pe_b/peij_2_2/d_acc [7]) );
  INV_X2 \pool/pool/pe_b/peij_2_2/add/fai_7/U2  ( .A(
        \pool/pool/pe_b/peij_2_2/add/fai_7/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_2/add/cprop [8]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_2/add/fai_7/U1  ( .A1(
        \pool/pool/pe_b/peij_2_2/add/notb [7]), .A2(
        \pool/pool/pe_b_o_data[2][18] ), .B1(
        \pool/pool/pe_b/peij_2_2/add/fai_7/n3 ), .B2(
        \pool/pool/pe_b/peij_2_2/add/cprop [7]), .ZN(
        \pool/pool/pe_b/peij_2_2/add/fai_7/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_8/U4  ( .A(
        \pool/pool/pe_b_o_data[2][19] ), .B(
        \pool/pool/pe_b/peij_2_2/add/notb [8]), .Z(
        \pool/pool/pe_b/peij_2_2/add/fai_8/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_8/U3  ( .A(
        \pool/pool/pe_b/peij_2_2/add/cprop [8]), .B(
        \pool/pool/pe_b/peij_2_2/add/fai_8/n3 ), .Z(
        \pool/pool/pe_b/peij_2_2/d_acc [8]) );
  INV_X2 \pool/pool/pe_b/peij_2_2/add/fai_8/U2  ( .A(
        \pool/pool/pe_b/peij_2_2/add/fai_8/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_2/add/cprop [9]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_2/add/fai_8/U1  ( .A1(
        \pool/pool/pe_b/peij_2_2/add/notb [8]), .A2(
        \pool/pool/pe_b_o_data[2][19] ), .B1(
        \pool/pool/pe_b/peij_2_2/add/fai_8/n3 ), .B2(
        \pool/pool/pe_b/peij_2_2/add/cprop [8]), .ZN(
        \pool/pool/pe_b/peij_2_2/add/fai_8/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_9/U4  ( .A(
        \pool/pool/pe_b_o_data[2][20] ), .B(
        \pool/pool/pe_b/peij_2_2/add/notb [9]), .Z(
        \pool/pool/pe_b/peij_2_2/add/fai_9/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_9/U3  ( .A(
        \pool/pool/pe_b/peij_2_2/add/cprop [9]), .B(
        \pool/pool/pe_b/peij_2_2/add/fai_9/n3 ), .Z(
        \pool/pool/pe_b/peij_2_2/d_acc [9]) );
  INV_X2 \pool/pool/pe_b/peij_2_2/add/fai_9/U2  ( .A(
        \pool/pool/pe_b/peij_2_2/add/fai_9/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_2/add/cprop [10]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_2/add/fai_9/U1  ( .A1(
        \pool/pool/pe_b/peij_2_2/add/notb [9]), .A2(
        \pool/pool/pe_b_o_data[2][20] ), .B1(
        \pool/pool/pe_b/peij_2_2/add/fai_9/n3 ), .B2(
        \pool/pool/pe_b/peij_2_2/add/cprop [9]), .ZN(
        \pool/pool/pe_b/peij_2_2/add/fai_9/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_10/U4  ( .A(
        \pool/pool/pe_b_o_data[2][21] ), .B(
        \pool/pool/pe_b/peij_2_2/add/notb [10]), .Z(
        \pool/pool/pe_b/peij_2_2/add/fai_10/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_2/add/fai_10/U3  ( .A(
        \pool/pool/pe_b/peij_2_2/add/cprop [10]), .B(
        \pool/pool/pe_b/peij_2_2/add/fai_10/n3 ), .Z(
        \pool/pool/pe_b/peij_2_2/d_acc [10]) );
  INV_X2 \pool/pool/pe_b/peij_2_2/add/fai_10/U2  ( .A(
        \pool/pool/pe_b/peij_2_2/add/fai_10/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_2/add/c_out ) );
  AOI22_X2 \pool/pool/pe_b/peij_2_2/add/fai_10/U1  ( .A1(
        \pool/pool/pe_b/peij_2_2/add/notb [10]), .A2(
        \pool/pool/pe_b_o_data[2][21] ), .B1(
        \pool/pool/pe_b/peij_2_2/add/fai_10/n3 ), .B2(
        \pool/pool/pe_b/peij_2_2/add/cprop [10]), .ZN(
        \pool/pool/pe_b/peij_2_2/add/fai_10/n1 ) );
  INV_X1 \pool/pool/pe_b/peij_2_3/U22  ( .A(\pool/pool/pe_b/n7 ), .ZN(
        \pool/pool/pe_b/peij_2_3/n16 ) );
  INV_X1 \pool/pool/pe_b/peij_2_3/U14  ( .A(\pool/pool/pe_b/n7 ), .ZN(
        \pool/pool/pe_b/peij_2_3/n12 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_3/U13  ( .A1(
        \pool/pool/pe_b/peij_2_3/d_acc [0]), .A2(\pool/pool/pe_b/peij_2_3/n18 ), .ZN(\pool/pool/pe_b/peij_2_3/n11 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_3/U12  ( .A1(
        \pool/pool/pe_b/peij_2_3/d_acc [1]), .A2(\pool/pool/pe_b/peij_2_3/n18 ), .ZN(\pool/pool/pe_b/peij_2_3/n10 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_3/U11  ( .A1(
        \pool/pool/pe_b/peij_2_3/d_acc [2]), .A2(\pool/pool/pe_b/peij_2_3/n18 ), .ZN(\pool/pool/pe_b/peij_2_3/n9 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_3/U10  ( .A1(
        \pool/pool/pe_b/peij_2_3/d_acc [3]), .A2(\pool/pool/pe_b/peij_2_3/n18 ), .ZN(\pool/pool/pe_b/peij_2_3/n8 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_3/U9  ( .A1(
        \pool/pool/pe_b/peij_2_3/d_acc [4]), .A2(\pool/pool/pe_b/peij_2_3/n18 ), .ZN(\pool/pool/pe_b/peij_2_3/n7 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_3/U8  ( .A1(
        \pool/pool/pe_b/peij_2_3/d_acc [5]), .A2(\pool/pool/pe_b/peij_2_3/n18 ), .ZN(\pool/pool/pe_b/peij_2_3/n6 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_3/U7  ( .A1(
        \pool/pool/pe_b/peij_2_3/d_acc [6]), .A2(\pool/pool/pe_b/peij_2_3/n18 ), .ZN(\pool/pool/pe_b/peij_2_3/n5 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_3/U6  ( .A1(
        \pool/pool/pe_b/peij_2_3/d_acc [7]), .A2(\pool/pool/pe_b/peij_2_3/n18 ), .ZN(\pool/pool/pe_b/peij_2_3/n4 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_3/U5  ( .A1(
        \pool/pool/pe_b/peij_2_3/d_acc [8]), .A2(\pool/pool/pe_b/peij_2_3/n18 ), .ZN(\pool/pool/pe_b/peij_2_3/n3 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_3/U4  ( .A1(
        \pool/pool/pe_b/peij_2_3/d_acc [9]), .A2(\pool/pool/pe_b/peij_2_3/n18 ), .ZN(\pool/pool/pe_b/peij_2_3/n2 ) );
  AND2_X1 \pool/pool/pe_b/peij_2_3/U3  ( .A1(
        \pool/pool/pe_b/peij_2_3/d_acc [10]), .A2(
        \pool/pool/pe_b/peij_2_3/n18 ), .ZN(\pool/pool/pe_b/peij_2_3/n1 ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_3/q_acc_reg[10]  ( .D(
        \pool/pool/pe_b/peij_2_3/n1 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_3/n16 ), .Q(\pool/pool/pe_b_o_data[2][10] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_3/q_acc_reg[9]  ( .D(
        \pool/pool/pe_b/peij_2_3/n2 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_3/n16 ), .Q(\pool/pool/pe_b_o_data[2][9] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_3/q_acc_reg[8]  ( .D(
        \pool/pool/pe_b/peij_2_3/n3 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_3/n16 ), .Q(\pool/pool/pe_b_o_data[2][8] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_3/q_acc_reg[7]  ( .D(
        \pool/pool/pe_b/peij_2_3/n4 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_3/n16 ), .Q(\pool/pool/pe_b_o_data[2][7] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_3/q_acc_reg[6]  ( .D(
        \pool/pool/pe_b/peij_2_3/n5 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_3/n16 ), .Q(\pool/pool/pe_b_o_data[2][6] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_3/q_acc_reg[5]  ( .D(
        \pool/pool/pe_b/peij_2_3/n6 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_3/n16 ), .Q(\pool/pool/pe_b_o_data[2][5] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_3/q_acc_reg[4]  ( .D(
        \pool/pool/pe_b/peij_2_3/n7 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_3/n16 ), .Q(\pool/pool/pe_b_o_data[2][4] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_3/q_acc_reg[3]  ( .D(
        \pool/pool/pe_b/peij_2_3/n8 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_3/n16 ), .Q(\pool/pool/pe_b_o_data[2][3] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_3/q_acc_reg[2]  ( .D(
        \pool/pool/pe_b/peij_2_3/n9 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_3/n16 ), .Q(\pool/pool/pe_b_o_data[2][2] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_3/q_acc_reg[1]  ( .D(
        \pool/pool/pe_b/peij_2_3/n10 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_3/n16 ), .Q(\pool/pool/pe_b_o_data[2][1] ) );
  DFFR_X1 \pool/pool/pe_b/peij_2_3/q_acc_reg[0]  ( .D(
        \pool/pool/pe_b/peij_2_3/n11 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_3/n16 ), .Q(\pool/pool/pe_b_o_data[2][0] ) );
  INV_X2 \pool/pool/pe_b/peij_2_3/U21  ( .A(\pool/sync_clr ), .ZN(
        \pool/pool/pe_b/peij_2_3/n18 ) );
  AND3_X2 \pool/pool/pe_b/peij_2_3/U20  ( .A1(\pool/pool/pe_b/int_pe_en[2][3] ), .A2(\pool/pool/pe_b/peij_2_3/n18 ), .A3(1'b1), .ZN(
        \pool/pool/pe_b/peij_2_3/n17 ) );
  AND2_X2 \pool/pool/pe_b/peij_2_3/U19  ( .A1(\pool/pool/pe_b_i_data[2][0] ), 
        .A2(\pool/pool/pe_b/peij_2_3/n17 ), .ZN(\pool/pool/pe_b/peij_2_3/N33 )
         );
  AND2_X2 \pool/pool/pe_b/peij_2_3/U18  ( .A1(\pool/pool/pe_b_i_data[2][1] ), 
        .A2(\pool/pool/pe_b/peij_2_3/n17 ), .ZN(\pool/pool/pe_b/peij_2_3/N34 )
         );
  AND2_X2 \pool/pool/pe_b/peij_2_3/U17  ( .A1(\pool/pool/pe_b_i_data[2][2] ), 
        .A2(\pool/pool/pe_b/peij_2_3/n17 ), .ZN(\pool/pool/pe_b/peij_2_3/N35 )
         );
  AND4_X4 \pool/pool/pe_b/peij_2_3/U16  ( .A1(1'b1), .A2(
        \pool/pool/pe_b_i_data[2][3] ), .A3(\pool/pool/pe_b/int_pe_en[2][3] ), 
        .A4(\pool/pool/pe_b/peij_2_3/n18 ), .ZN(\pool/pool/pe_b/peij_2_3/N36 )
         );
  DFFR_X1 \pool/pool/pe_b/peij_2_3/q_im_reg[0]  ( .D(
        \pool/pool/pe_b/peij_2_3/N33 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_3/n12 ), .Q(\pool/pool/pe_b/peij_2_3/sgnext [0]) );
  DFFR_X1 \pool/pool/pe_b/peij_2_3/q_im_reg[1]  ( .D(
        \pool/pool/pe_b/peij_2_3/N34 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_3/n12 ), .Q(\pool/pool/pe_b/peij_2_3/sgnext [1]) );
  DFFR_X1 \pool/pool/pe_b/peij_2_3/q_im_reg[2]  ( .D(
        \pool/pool/pe_b/peij_2_3/N35 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_3/n12 ), .Q(\pool/pool/pe_b/peij_2_3/sgnext [2]) );
  DFFR_X1 \pool/pool/pe_b/peij_2_3/q_im_reg[3]  ( .D(
        \pool/pool/pe_b/peij_2_3/N36 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_3/n12 ), .Q(\pool/pool/pe_b/peij_2_3/sgnext_10 ) );
  SDFFR_X1 \pool/pool/pe_b/peij_2_3/q_k_reg  ( .D(1'b0), .SI(
        \pool/pool/pe_b/peij_2_3/n18 ), .SE(1'b0), .CK(clk), .RN(
        \pool/pool/pe_b/peij_2_3/n12 ), .Q(\pool/pool/pe_b/peij_2_3/q_k ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/U11  ( .A(
        \pool/pool/pe_b/peij_2_3/sgnext [0]), .B(\pool/pool/pe_b/peij_2_3/q_k ), .Z(\pool/pool/pe_b/peij_2_3/add/notb [0]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/U10  ( .A(
        \pool/pool/pe_b/peij_2_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_3/q_k ), .Z(\pool/pool/pe_b/peij_2_3/add/notb [10]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/U9  ( .A(
        \pool/pool/pe_b/peij_2_3/sgnext [1]), .B(\pool/pool/pe_b/peij_2_3/q_k ), .Z(\pool/pool/pe_b/peij_2_3/add/notb [1]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/U8  ( .A(
        \pool/pool/pe_b/peij_2_3/sgnext [2]), .B(\pool/pool/pe_b/peij_2_3/q_k ), .Z(\pool/pool/pe_b/peij_2_3/add/notb [2]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/U7  ( .A(
        \pool/pool/pe_b/peij_2_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_3/q_k ), .Z(\pool/pool/pe_b/peij_2_3/add/notb [3]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/U6  ( .A(
        \pool/pool/pe_b/peij_2_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_3/q_k ), .Z(\pool/pool/pe_b/peij_2_3/add/notb [4]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/U5  ( .A(
        \pool/pool/pe_b/peij_2_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_3/q_k ), .Z(\pool/pool/pe_b/peij_2_3/add/notb [5]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/U4  ( .A(
        \pool/pool/pe_b/peij_2_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_3/q_k ), .Z(\pool/pool/pe_b/peij_2_3/add/notb [6]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/U3  ( .A(
        \pool/pool/pe_b/peij_2_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_3/q_k ), .Z(\pool/pool/pe_b/peij_2_3/add/notb [7]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/U2  ( .A(
        \pool/pool/pe_b/peij_2_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_3/q_k ), .Z(\pool/pool/pe_b/peij_2_3/add/notb [8]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/U1  ( .A(
        \pool/pool/pe_b/peij_2_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_2_3/q_k ), .Z(\pool/pool/pe_b/peij_2_3/add/notb [9]) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_0/U4  ( .A(
        \pool/pool/pe_b_o_data[2][0] ), .B(
        \pool/pool/pe_b/peij_2_3/add/notb [0]), .Z(
        \pool/pool/pe_b/peij_2_3/add/fai_0/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_0/U3  ( .A(
        \pool/pool/pe_b/peij_2_3/q_k ), .B(
        \pool/pool/pe_b/peij_2_3/add/fai_0/n3 ), .Z(
        \pool/pool/pe_b/peij_2_3/d_acc [0]) );
  INV_X2 \pool/pool/pe_b/peij_2_3/add/fai_0/U2  ( .A(
        \pool/pool/pe_b/peij_2_3/add/fai_0/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_3/add/cprop [1]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_3/add/fai_0/U1  ( .A1(
        \pool/pool/pe_b/peij_2_3/add/notb [0]), .A2(
        \pool/pool/pe_b_o_data[2][0] ), .B1(
        \pool/pool/pe_b/peij_2_3/add/fai_0/n3 ), .B2(
        \pool/pool/pe_b/peij_2_3/q_k ), .ZN(
        \pool/pool/pe_b/peij_2_3/add/fai_0/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_1/U4  ( .A(
        \pool/pool/pe_b_o_data[2][1] ), .B(
        \pool/pool/pe_b/peij_2_3/add/notb [1]), .Z(
        \pool/pool/pe_b/peij_2_3/add/fai_1/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_1/U3  ( .A(
        \pool/pool/pe_b/peij_2_3/add/cprop [1]), .B(
        \pool/pool/pe_b/peij_2_3/add/fai_1/n3 ), .Z(
        \pool/pool/pe_b/peij_2_3/d_acc [1]) );
  INV_X2 \pool/pool/pe_b/peij_2_3/add/fai_1/U2  ( .A(
        \pool/pool/pe_b/peij_2_3/add/fai_1/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_3/add/cprop [2]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_3/add/fai_1/U1  ( .A1(
        \pool/pool/pe_b/peij_2_3/add/notb [1]), .A2(
        \pool/pool/pe_b_o_data[2][1] ), .B1(
        \pool/pool/pe_b/peij_2_3/add/fai_1/n3 ), .B2(
        \pool/pool/pe_b/peij_2_3/add/cprop [1]), .ZN(
        \pool/pool/pe_b/peij_2_3/add/fai_1/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_2/U4  ( .A(
        \pool/pool/pe_b_o_data[2][2] ), .B(
        \pool/pool/pe_b/peij_2_3/add/notb [2]), .Z(
        \pool/pool/pe_b/peij_2_3/add/fai_2/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_2/U3  ( .A(
        \pool/pool/pe_b/peij_2_3/add/cprop [2]), .B(
        \pool/pool/pe_b/peij_2_3/add/fai_2/n3 ), .Z(
        \pool/pool/pe_b/peij_2_3/d_acc [2]) );
  INV_X2 \pool/pool/pe_b/peij_2_3/add/fai_2/U2  ( .A(
        \pool/pool/pe_b/peij_2_3/add/fai_2/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_3/add/cprop [3]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_3/add/fai_2/U1  ( .A1(
        \pool/pool/pe_b/peij_2_3/add/notb [2]), .A2(
        \pool/pool/pe_b_o_data[2][2] ), .B1(
        \pool/pool/pe_b/peij_2_3/add/fai_2/n3 ), .B2(
        \pool/pool/pe_b/peij_2_3/add/cprop [2]), .ZN(
        \pool/pool/pe_b/peij_2_3/add/fai_2/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_3/U4  ( .A(
        \pool/pool/pe_b_o_data[2][3] ), .B(
        \pool/pool/pe_b/peij_2_3/add/notb [3]), .Z(
        \pool/pool/pe_b/peij_2_3/add/fai_3/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_3/U3  ( .A(
        \pool/pool/pe_b/peij_2_3/add/cprop [3]), .B(
        \pool/pool/pe_b/peij_2_3/add/fai_3/n3 ), .Z(
        \pool/pool/pe_b/peij_2_3/d_acc [3]) );
  INV_X2 \pool/pool/pe_b/peij_2_3/add/fai_3/U2  ( .A(
        \pool/pool/pe_b/peij_2_3/add/fai_3/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_3/add/cprop [4]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_3/add/fai_3/U1  ( .A1(
        \pool/pool/pe_b/peij_2_3/add/notb [3]), .A2(
        \pool/pool/pe_b_o_data[2][3] ), .B1(
        \pool/pool/pe_b/peij_2_3/add/fai_3/n3 ), .B2(
        \pool/pool/pe_b/peij_2_3/add/cprop [3]), .ZN(
        \pool/pool/pe_b/peij_2_3/add/fai_3/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_4/U4  ( .A(
        \pool/pool/pe_b_o_data[2][4] ), .B(
        \pool/pool/pe_b/peij_2_3/add/notb [4]), .Z(
        \pool/pool/pe_b/peij_2_3/add/fai_4/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_4/U3  ( .A(
        \pool/pool/pe_b/peij_2_3/add/cprop [4]), .B(
        \pool/pool/pe_b/peij_2_3/add/fai_4/n3 ), .Z(
        \pool/pool/pe_b/peij_2_3/d_acc [4]) );
  INV_X2 \pool/pool/pe_b/peij_2_3/add/fai_4/U2  ( .A(
        \pool/pool/pe_b/peij_2_3/add/fai_4/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_3/add/cprop [5]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_3/add/fai_4/U1  ( .A1(
        \pool/pool/pe_b/peij_2_3/add/notb [4]), .A2(
        \pool/pool/pe_b_o_data[2][4] ), .B1(
        \pool/pool/pe_b/peij_2_3/add/fai_4/n3 ), .B2(
        \pool/pool/pe_b/peij_2_3/add/cprop [4]), .ZN(
        \pool/pool/pe_b/peij_2_3/add/fai_4/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_5/U4  ( .A(
        \pool/pool/pe_b_o_data[2][5] ), .B(
        \pool/pool/pe_b/peij_2_3/add/notb [5]), .Z(
        \pool/pool/pe_b/peij_2_3/add/fai_5/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_5/U3  ( .A(
        \pool/pool/pe_b/peij_2_3/add/cprop [5]), .B(
        \pool/pool/pe_b/peij_2_3/add/fai_5/n3 ), .Z(
        \pool/pool/pe_b/peij_2_3/d_acc [5]) );
  INV_X2 \pool/pool/pe_b/peij_2_3/add/fai_5/U2  ( .A(
        \pool/pool/pe_b/peij_2_3/add/fai_5/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_3/add/cprop [6]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_3/add/fai_5/U1  ( .A1(
        \pool/pool/pe_b/peij_2_3/add/notb [5]), .A2(
        \pool/pool/pe_b_o_data[2][5] ), .B1(
        \pool/pool/pe_b/peij_2_3/add/fai_5/n3 ), .B2(
        \pool/pool/pe_b/peij_2_3/add/cprop [5]), .ZN(
        \pool/pool/pe_b/peij_2_3/add/fai_5/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_6/U4  ( .A(
        \pool/pool/pe_b_o_data[2][6] ), .B(
        \pool/pool/pe_b/peij_2_3/add/notb [6]), .Z(
        \pool/pool/pe_b/peij_2_3/add/fai_6/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_6/U3  ( .A(
        \pool/pool/pe_b/peij_2_3/add/cprop [6]), .B(
        \pool/pool/pe_b/peij_2_3/add/fai_6/n3 ), .Z(
        \pool/pool/pe_b/peij_2_3/d_acc [6]) );
  INV_X2 \pool/pool/pe_b/peij_2_3/add/fai_6/U2  ( .A(
        \pool/pool/pe_b/peij_2_3/add/fai_6/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_3/add/cprop [7]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_3/add/fai_6/U1  ( .A1(
        \pool/pool/pe_b/peij_2_3/add/notb [6]), .A2(
        \pool/pool/pe_b_o_data[2][6] ), .B1(
        \pool/pool/pe_b/peij_2_3/add/fai_6/n3 ), .B2(
        \pool/pool/pe_b/peij_2_3/add/cprop [6]), .ZN(
        \pool/pool/pe_b/peij_2_3/add/fai_6/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_7/U4  ( .A(
        \pool/pool/pe_b_o_data[2][7] ), .B(
        \pool/pool/pe_b/peij_2_3/add/notb [7]), .Z(
        \pool/pool/pe_b/peij_2_3/add/fai_7/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_7/U3  ( .A(
        \pool/pool/pe_b/peij_2_3/add/cprop [7]), .B(
        \pool/pool/pe_b/peij_2_3/add/fai_7/n3 ), .Z(
        \pool/pool/pe_b/peij_2_3/d_acc [7]) );
  INV_X2 \pool/pool/pe_b/peij_2_3/add/fai_7/U2  ( .A(
        \pool/pool/pe_b/peij_2_3/add/fai_7/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_3/add/cprop [8]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_3/add/fai_7/U1  ( .A1(
        \pool/pool/pe_b/peij_2_3/add/notb [7]), .A2(
        \pool/pool/pe_b_o_data[2][7] ), .B1(
        \pool/pool/pe_b/peij_2_3/add/fai_7/n3 ), .B2(
        \pool/pool/pe_b/peij_2_3/add/cprop [7]), .ZN(
        \pool/pool/pe_b/peij_2_3/add/fai_7/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_8/U4  ( .A(
        \pool/pool/pe_b_o_data[2][8] ), .B(
        \pool/pool/pe_b/peij_2_3/add/notb [8]), .Z(
        \pool/pool/pe_b/peij_2_3/add/fai_8/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_8/U3  ( .A(
        \pool/pool/pe_b/peij_2_3/add/cprop [8]), .B(
        \pool/pool/pe_b/peij_2_3/add/fai_8/n3 ), .Z(
        \pool/pool/pe_b/peij_2_3/d_acc [8]) );
  INV_X2 \pool/pool/pe_b/peij_2_3/add/fai_8/U2  ( .A(
        \pool/pool/pe_b/peij_2_3/add/fai_8/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_3/add/cprop [9]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_3/add/fai_8/U1  ( .A1(
        \pool/pool/pe_b/peij_2_3/add/notb [8]), .A2(
        \pool/pool/pe_b_o_data[2][8] ), .B1(
        \pool/pool/pe_b/peij_2_3/add/fai_8/n3 ), .B2(
        \pool/pool/pe_b/peij_2_3/add/cprop [8]), .ZN(
        \pool/pool/pe_b/peij_2_3/add/fai_8/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_9/U4  ( .A(
        \pool/pool/pe_b_o_data[2][9] ), .B(
        \pool/pool/pe_b/peij_2_3/add/notb [9]), .Z(
        \pool/pool/pe_b/peij_2_3/add/fai_9/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_9/U3  ( .A(
        \pool/pool/pe_b/peij_2_3/add/cprop [9]), .B(
        \pool/pool/pe_b/peij_2_3/add/fai_9/n3 ), .Z(
        \pool/pool/pe_b/peij_2_3/d_acc [9]) );
  INV_X2 \pool/pool/pe_b/peij_2_3/add/fai_9/U2  ( .A(
        \pool/pool/pe_b/peij_2_3/add/fai_9/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_3/add/cprop [10]) );
  AOI22_X2 \pool/pool/pe_b/peij_2_3/add/fai_9/U1  ( .A1(
        \pool/pool/pe_b/peij_2_3/add/notb [9]), .A2(
        \pool/pool/pe_b_o_data[2][9] ), .B1(
        \pool/pool/pe_b/peij_2_3/add/fai_9/n3 ), .B2(
        \pool/pool/pe_b/peij_2_3/add/cprop [9]), .ZN(
        \pool/pool/pe_b/peij_2_3/add/fai_9/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_10/U4  ( .A(
        \pool/pool/pe_b_o_data[2][10] ), .B(
        \pool/pool/pe_b/peij_2_3/add/notb [10]), .Z(
        \pool/pool/pe_b/peij_2_3/add/fai_10/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_2_3/add/fai_10/U3  ( .A(
        \pool/pool/pe_b/peij_2_3/add/cprop [10]), .B(
        \pool/pool/pe_b/peij_2_3/add/fai_10/n3 ), .Z(
        \pool/pool/pe_b/peij_2_3/d_acc [10]) );
  INV_X2 \pool/pool/pe_b/peij_2_3/add/fai_10/U2  ( .A(
        \pool/pool/pe_b/peij_2_3/add/fai_10/n1 ), .ZN(
        \pool/pool/pe_b/peij_2_3/add/c_out ) );
  AOI22_X2 \pool/pool/pe_b/peij_2_3/add/fai_10/U1  ( .A1(
        \pool/pool/pe_b/peij_2_3/add/notb [10]), .A2(
        \pool/pool/pe_b_o_data[2][10] ), .B1(
        \pool/pool/pe_b/peij_2_3/add/fai_10/n3 ), .B2(
        \pool/pool/pe_b/peij_2_3/add/cprop [10]), .ZN(
        \pool/pool/pe_b/peij_2_3/add/fai_10/n1 ) );
  INV_X1 \pool/pool/pe_b/peij_3_0/U22  ( .A(\pool/pool/pe_b/n7 ), .ZN(
        \pool/pool/pe_b/peij_3_0/n16 ) );
  INV_X1 \pool/pool/pe_b/peij_3_0/U14  ( .A(\pool/pool/pe_b/n7 ), .ZN(
        \pool/pool/pe_b/peij_3_0/n12 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_0/U13  ( .A1(
        \pool/pool/pe_b/peij_3_0/d_acc [0]), .A2(\pool/pool/pe_b/peij_3_0/n18 ), .ZN(\pool/pool/pe_b/peij_3_0/n11 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_0/U12  ( .A1(
        \pool/pool/pe_b/peij_3_0/d_acc [1]), .A2(\pool/pool/pe_b/peij_3_0/n18 ), .ZN(\pool/pool/pe_b/peij_3_0/n10 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_0/U11  ( .A1(
        \pool/pool/pe_b/peij_3_0/d_acc [2]), .A2(\pool/pool/pe_b/peij_3_0/n18 ), .ZN(\pool/pool/pe_b/peij_3_0/n9 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_0/U10  ( .A1(
        \pool/pool/pe_b/peij_3_0/d_acc [3]), .A2(\pool/pool/pe_b/peij_3_0/n18 ), .ZN(\pool/pool/pe_b/peij_3_0/n8 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_0/U9  ( .A1(
        \pool/pool/pe_b/peij_3_0/d_acc [4]), .A2(\pool/pool/pe_b/peij_3_0/n18 ), .ZN(\pool/pool/pe_b/peij_3_0/n7 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_0/U8  ( .A1(
        \pool/pool/pe_b/peij_3_0/d_acc [5]), .A2(\pool/pool/pe_b/peij_3_0/n18 ), .ZN(\pool/pool/pe_b/peij_3_0/n6 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_0/U7  ( .A1(
        \pool/pool/pe_b/peij_3_0/d_acc [6]), .A2(\pool/pool/pe_b/peij_3_0/n18 ), .ZN(\pool/pool/pe_b/peij_3_0/n5 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_0/U6  ( .A1(
        \pool/pool/pe_b/peij_3_0/d_acc [7]), .A2(\pool/pool/pe_b/peij_3_0/n18 ), .ZN(\pool/pool/pe_b/peij_3_0/n4 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_0/U5  ( .A1(
        \pool/pool/pe_b/peij_3_0/d_acc [8]), .A2(\pool/pool/pe_b/peij_3_0/n18 ), .ZN(\pool/pool/pe_b/peij_3_0/n3 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_0/U4  ( .A1(
        \pool/pool/pe_b/peij_3_0/d_acc [9]), .A2(\pool/pool/pe_b/peij_3_0/n18 ), .ZN(\pool/pool/pe_b/peij_3_0/n2 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_0/U3  ( .A1(
        \pool/pool/pe_b/peij_3_0/d_acc [10]), .A2(
        \pool/pool/pe_b/peij_3_0/n18 ), .ZN(\pool/pool/pe_b/peij_3_0/n1 ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_0/q_acc_reg[10]  ( .D(
        \pool/pool/pe_b/peij_3_0/n1 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_0/n16 ), .Q(\pool/pool/pe_b_o_data[3][43] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_0/q_acc_reg[9]  ( .D(
        \pool/pool/pe_b/peij_3_0/n2 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_0/n16 ), .Q(\pool/pool/pe_b_o_data[3][42] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_0/q_acc_reg[8]  ( .D(
        \pool/pool/pe_b/peij_3_0/n3 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_0/n16 ), .Q(\pool/pool/pe_b_o_data[3][41] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_0/q_acc_reg[7]  ( .D(
        \pool/pool/pe_b/peij_3_0/n4 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_0/n16 ), .Q(\pool/pool/pe_b_o_data[3][40] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_0/q_acc_reg[6]  ( .D(
        \pool/pool/pe_b/peij_3_0/n5 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_0/n16 ), .Q(\pool/pool/pe_b_o_data[3][39] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_0/q_acc_reg[5]  ( .D(
        \pool/pool/pe_b/peij_3_0/n6 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_0/n16 ), .Q(\pool/pool/pe_b_o_data[3][38] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_0/q_acc_reg[4]  ( .D(
        \pool/pool/pe_b/peij_3_0/n7 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_0/n16 ), .Q(\pool/pool/pe_b_o_data[3][37] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_0/q_acc_reg[3]  ( .D(
        \pool/pool/pe_b/peij_3_0/n8 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_0/n16 ), .Q(\pool/pool/pe_b_o_data[3][36] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_0/q_acc_reg[2]  ( .D(
        \pool/pool/pe_b/peij_3_0/n9 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_0/n16 ), .Q(\pool/pool/pe_b_o_data[3][35] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_0/q_acc_reg[1]  ( .D(
        \pool/pool/pe_b/peij_3_0/n10 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_0/n16 ), .Q(\pool/pool/pe_b_o_data[3][34] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_0/q_acc_reg[0]  ( .D(
        \pool/pool/pe_b/peij_3_0/n11 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_0/n16 ), .Q(\pool/pool/pe_b_o_data[3][33] ) );
  INV_X2 \pool/pool/pe_b/peij_3_0/U21  ( .A(\pool/sync_clr ), .ZN(
        \pool/pool/pe_b/peij_3_0/n18 ) );
  AND3_X2 \pool/pool/pe_b/peij_3_0/U20  ( .A1(\pool/pool/pe_b/int_pe_en[3][0] ), .A2(\pool/pool/pe_b/peij_3_0/n18 ), .A3(1'b1), .ZN(
        \pool/pool/pe_b/peij_3_0/n17 ) );
  AND2_X2 \pool/pool/pe_b/peij_3_0/U19  ( .A1(\pool/pool/pe_b_i_data[3][12] ), 
        .A2(\pool/pool/pe_b/peij_3_0/n17 ), .ZN(\pool/pool/pe_b/peij_3_0/N33 )
         );
  AND2_X2 \pool/pool/pe_b/peij_3_0/U18  ( .A1(\pool/pool/pe_b_i_data[3][13] ), 
        .A2(\pool/pool/pe_b/peij_3_0/n17 ), .ZN(\pool/pool/pe_b/peij_3_0/N34 )
         );
  AND2_X2 \pool/pool/pe_b/peij_3_0/U17  ( .A1(\pool/pool/pe_b_i_data[3][14] ), 
        .A2(\pool/pool/pe_b/peij_3_0/n17 ), .ZN(\pool/pool/pe_b/peij_3_0/N35 )
         );
  AND4_X4 \pool/pool/pe_b/peij_3_0/U16  ( .A1(1'b1), .A2(
        \pool/pool/pe_b_i_data[3][15] ), .A3(\pool/pool/pe_b/int_pe_en[3][0] ), 
        .A4(\pool/pool/pe_b/peij_3_0/n18 ), .ZN(\pool/pool/pe_b/peij_3_0/N36 )
         );
  DFFR_X1 \pool/pool/pe_b/peij_3_0/q_im_reg[0]  ( .D(
        \pool/pool/pe_b/peij_3_0/N33 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_0/n12 ), .Q(\pool/pool/pe_b/peij_3_0/sgnext [0]) );
  DFFR_X1 \pool/pool/pe_b/peij_3_0/q_im_reg[1]  ( .D(
        \pool/pool/pe_b/peij_3_0/N34 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_0/n12 ), .Q(\pool/pool/pe_b/peij_3_0/sgnext [1]) );
  DFFR_X1 \pool/pool/pe_b/peij_3_0/q_im_reg[2]  ( .D(
        \pool/pool/pe_b/peij_3_0/N35 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_0/n12 ), .Q(\pool/pool/pe_b/peij_3_0/sgnext [2]) );
  DFFR_X1 \pool/pool/pe_b/peij_3_0/q_im_reg[3]  ( .D(
        \pool/pool/pe_b/peij_3_0/N36 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_0/n12 ), .Q(\pool/pool/pe_b/peij_3_0/sgnext_10 ) );
  SDFFR_X1 \pool/pool/pe_b/peij_3_0/q_k_reg  ( .D(1'b0), .SI(
        \pool/pool/pe_b/peij_3_0/n18 ), .SE(1'b0), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_0/n12 ), .Q(\pool/pool/pe_b/peij_3_0/q_k ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/U11  ( .A(
        \pool/pool/pe_b/peij_3_0/sgnext [0]), .B(\pool/pool/pe_b/peij_3_0/q_k ), .Z(\pool/pool/pe_b/peij_3_0/add/notb [0]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/U10  ( .A(
        \pool/pool/pe_b/peij_3_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_0/q_k ), .Z(\pool/pool/pe_b/peij_3_0/add/notb [10]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/U9  ( .A(
        \pool/pool/pe_b/peij_3_0/sgnext [1]), .B(\pool/pool/pe_b/peij_3_0/q_k ), .Z(\pool/pool/pe_b/peij_3_0/add/notb [1]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/U8  ( .A(
        \pool/pool/pe_b/peij_3_0/sgnext [2]), .B(\pool/pool/pe_b/peij_3_0/q_k ), .Z(\pool/pool/pe_b/peij_3_0/add/notb [2]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/U7  ( .A(
        \pool/pool/pe_b/peij_3_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_0/q_k ), .Z(\pool/pool/pe_b/peij_3_0/add/notb [3]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/U6  ( .A(
        \pool/pool/pe_b/peij_3_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_0/q_k ), .Z(\pool/pool/pe_b/peij_3_0/add/notb [4]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/U5  ( .A(
        \pool/pool/pe_b/peij_3_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_0/q_k ), .Z(\pool/pool/pe_b/peij_3_0/add/notb [5]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/U4  ( .A(
        \pool/pool/pe_b/peij_3_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_0/q_k ), .Z(\pool/pool/pe_b/peij_3_0/add/notb [6]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/U3  ( .A(
        \pool/pool/pe_b/peij_3_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_0/q_k ), .Z(\pool/pool/pe_b/peij_3_0/add/notb [7]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/U2  ( .A(
        \pool/pool/pe_b/peij_3_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_0/q_k ), .Z(\pool/pool/pe_b/peij_3_0/add/notb [8]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/U1  ( .A(
        \pool/pool/pe_b/peij_3_0/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_0/q_k ), .Z(\pool/pool/pe_b/peij_3_0/add/notb [9]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_0/U4  ( .A(
        \pool/pool/pe_b_o_data[3][33] ), .B(
        \pool/pool/pe_b/peij_3_0/add/notb [0]), .Z(
        \pool/pool/pe_b/peij_3_0/add/fai_0/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_0/U3  ( .A(
        \pool/pool/pe_b/peij_3_0/q_k ), .B(
        \pool/pool/pe_b/peij_3_0/add/fai_0/n3 ), .Z(
        \pool/pool/pe_b/peij_3_0/d_acc [0]) );
  INV_X2 \pool/pool/pe_b/peij_3_0/add/fai_0/U2  ( .A(
        \pool/pool/pe_b/peij_3_0/add/fai_0/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_0/add/cprop [1]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_0/add/fai_0/U1  ( .A1(
        \pool/pool/pe_b/peij_3_0/add/notb [0]), .A2(
        \pool/pool/pe_b_o_data[3][33] ), .B1(
        \pool/pool/pe_b/peij_3_0/add/fai_0/n3 ), .B2(
        \pool/pool/pe_b/peij_3_0/q_k ), .ZN(
        \pool/pool/pe_b/peij_3_0/add/fai_0/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_1/U4  ( .A(
        \pool/pool/pe_b_o_data[3][34] ), .B(
        \pool/pool/pe_b/peij_3_0/add/notb [1]), .Z(
        \pool/pool/pe_b/peij_3_0/add/fai_1/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_1/U3  ( .A(
        \pool/pool/pe_b/peij_3_0/add/cprop [1]), .B(
        \pool/pool/pe_b/peij_3_0/add/fai_1/n3 ), .Z(
        \pool/pool/pe_b/peij_3_0/d_acc [1]) );
  INV_X2 \pool/pool/pe_b/peij_3_0/add/fai_1/U2  ( .A(
        \pool/pool/pe_b/peij_3_0/add/fai_1/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_0/add/cprop [2]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_0/add/fai_1/U1  ( .A1(
        \pool/pool/pe_b/peij_3_0/add/notb [1]), .A2(
        \pool/pool/pe_b_o_data[3][34] ), .B1(
        \pool/pool/pe_b/peij_3_0/add/fai_1/n3 ), .B2(
        \pool/pool/pe_b/peij_3_0/add/cprop [1]), .ZN(
        \pool/pool/pe_b/peij_3_0/add/fai_1/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_2/U4  ( .A(
        \pool/pool/pe_b_o_data[3][35] ), .B(
        \pool/pool/pe_b/peij_3_0/add/notb [2]), .Z(
        \pool/pool/pe_b/peij_3_0/add/fai_2/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_2/U3  ( .A(
        \pool/pool/pe_b/peij_3_0/add/cprop [2]), .B(
        \pool/pool/pe_b/peij_3_0/add/fai_2/n3 ), .Z(
        \pool/pool/pe_b/peij_3_0/d_acc [2]) );
  INV_X2 \pool/pool/pe_b/peij_3_0/add/fai_2/U2  ( .A(
        \pool/pool/pe_b/peij_3_0/add/fai_2/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_0/add/cprop [3]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_0/add/fai_2/U1  ( .A1(
        \pool/pool/pe_b/peij_3_0/add/notb [2]), .A2(
        \pool/pool/pe_b_o_data[3][35] ), .B1(
        \pool/pool/pe_b/peij_3_0/add/fai_2/n3 ), .B2(
        \pool/pool/pe_b/peij_3_0/add/cprop [2]), .ZN(
        \pool/pool/pe_b/peij_3_0/add/fai_2/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_3/U4  ( .A(
        \pool/pool/pe_b_o_data[3][36] ), .B(
        \pool/pool/pe_b/peij_3_0/add/notb [3]), .Z(
        \pool/pool/pe_b/peij_3_0/add/fai_3/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_3/U3  ( .A(
        \pool/pool/pe_b/peij_3_0/add/cprop [3]), .B(
        \pool/pool/pe_b/peij_3_0/add/fai_3/n3 ), .Z(
        \pool/pool/pe_b/peij_3_0/d_acc [3]) );
  INV_X2 \pool/pool/pe_b/peij_3_0/add/fai_3/U2  ( .A(
        \pool/pool/pe_b/peij_3_0/add/fai_3/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_0/add/cprop [4]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_0/add/fai_3/U1  ( .A1(
        \pool/pool/pe_b/peij_3_0/add/notb [3]), .A2(
        \pool/pool/pe_b_o_data[3][36] ), .B1(
        \pool/pool/pe_b/peij_3_0/add/fai_3/n3 ), .B2(
        \pool/pool/pe_b/peij_3_0/add/cprop [3]), .ZN(
        \pool/pool/pe_b/peij_3_0/add/fai_3/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_4/U4  ( .A(
        \pool/pool/pe_b_o_data[3][37] ), .B(
        \pool/pool/pe_b/peij_3_0/add/notb [4]), .Z(
        \pool/pool/pe_b/peij_3_0/add/fai_4/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_4/U3  ( .A(
        \pool/pool/pe_b/peij_3_0/add/cprop [4]), .B(
        \pool/pool/pe_b/peij_3_0/add/fai_4/n3 ), .Z(
        \pool/pool/pe_b/peij_3_0/d_acc [4]) );
  INV_X2 \pool/pool/pe_b/peij_3_0/add/fai_4/U2  ( .A(
        \pool/pool/pe_b/peij_3_0/add/fai_4/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_0/add/cprop [5]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_0/add/fai_4/U1  ( .A1(
        \pool/pool/pe_b/peij_3_0/add/notb [4]), .A2(
        \pool/pool/pe_b_o_data[3][37] ), .B1(
        \pool/pool/pe_b/peij_3_0/add/fai_4/n3 ), .B2(
        \pool/pool/pe_b/peij_3_0/add/cprop [4]), .ZN(
        \pool/pool/pe_b/peij_3_0/add/fai_4/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_5/U4  ( .A(
        \pool/pool/pe_b_o_data[3][38] ), .B(
        \pool/pool/pe_b/peij_3_0/add/notb [5]), .Z(
        \pool/pool/pe_b/peij_3_0/add/fai_5/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_5/U3  ( .A(
        \pool/pool/pe_b/peij_3_0/add/cprop [5]), .B(
        \pool/pool/pe_b/peij_3_0/add/fai_5/n3 ), .Z(
        \pool/pool/pe_b/peij_3_0/d_acc [5]) );
  INV_X2 \pool/pool/pe_b/peij_3_0/add/fai_5/U2  ( .A(
        \pool/pool/pe_b/peij_3_0/add/fai_5/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_0/add/cprop [6]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_0/add/fai_5/U1  ( .A1(
        \pool/pool/pe_b/peij_3_0/add/notb [5]), .A2(
        \pool/pool/pe_b_o_data[3][38] ), .B1(
        \pool/pool/pe_b/peij_3_0/add/fai_5/n3 ), .B2(
        \pool/pool/pe_b/peij_3_0/add/cprop [5]), .ZN(
        \pool/pool/pe_b/peij_3_0/add/fai_5/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_6/U4  ( .A(
        \pool/pool/pe_b_o_data[3][39] ), .B(
        \pool/pool/pe_b/peij_3_0/add/notb [6]), .Z(
        \pool/pool/pe_b/peij_3_0/add/fai_6/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_6/U3  ( .A(
        \pool/pool/pe_b/peij_3_0/add/cprop [6]), .B(
        \pool/pool/pe_b/peij_3_0/add/fai_6/n3 ), .Z(
        \pool/pool/pe_b/peij_3_0/d_acc [6]) );
  INV_X2 \pool/pool/pe_b/peij_3_0/add/fai_6/U2  ( .A(
        \pool/pool/pe_b/peij_3_0/add/fai_6/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_0/add/cprop [7]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_0/add/fai_6/U1  ( .A1(
        \pool/pool/pe_b/peij_3_0/add/notb [6]), .A2(
        \pool/pool/pe_b_o_data[3][39] ), .B1(
        \pool/pool/pe_b/peij_3_0/add/fai_6/n3 ), .B2(
        \pool/pool/pe_b/peij_3_0/add/cprop [6]), .ZN(
        \pool/pool/pe_b/peij_3_0/add/fai_6/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_7/U4  ( .A(
        \pool/pool/pe_b_o_data[3][40] ), .B(
        \pool/pool/pe_b/peij_3_0/add/notb [7]), .Z(
        \pool/pool/pe_b/peij_3_0/add/fai_7/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_7/U3  ( .A(
        \pool/pool/pe_b/peij_3_0/add/cprop [7]), .B(
        \pool/pool/pe_b/peij_3_0/add/fai_7/n3 ), .Z(
        \pool/pool/pe_b/peij_3_0/d_acc [7]) );
  INV_X2 \pool/pool/pe_b/peij_3_0/add/fai_7/U2  ( .A(
        \pool/pool/pe_b/peij_3_0/add/fai_7/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_0/add/cprop [8]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_0/add/fai_7/U1  ( .A1(
        \pool/pool/pe_b/peij_3_0/add/notb [7]), .A2(
        \pool/pool/pe_b_o_data[3][40] ), .B1(
        \pool/pool/pe_b/peij_3_0/add/fai_7/n3 ), .B2(
        \pool/pool/pe_b/peij_3_0/add/cprop [7]), .ZN(
        \pool/pool/pe_b/peij_3_0/add/fai_7/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_8/U4  ( .A(
        \pool/pool/pe_b_o_data[3][41] ), .B(
        \pool/pool/pe_b/peij_3_0/add/notb [8]), .Z(
        \pool/pool/pe_b/peij_3_0/add/fai_8/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_8/U3  ( .A(
        \pool/pool/pe_b/peij_3_0/add/cprop [8]), .B(
        \pool/pool/pe_b/peij_3_0/add/fai_8/n3 ), .Z(
        \pool/pool/pe_b/peij_3_0/d_acc [8]) );
  INV_X2 \pool/pool/pe_b/peij_3_0/add/fai_8/U2  ( .A(
        \pool/pool/pe_b/peij_3_0/add/fai_8/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_0/add/cprop [9]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_0/add/fai_8/U1  ( .A1(
        \pool/pool/pe_b/peij_3_0/add/notb [8]), .A2(
        \pool/pool/pe_b_o_data[3][41] ), .B1(
        \pool/pool/pe_b/peij_3_0/add/fai_8/n3 ), .B2(
        \pool/pool/pe_b/peij_3_0/add/cprop [8]), .ZN(
        \pool/pool/pe_b/peij_3_0/add/fai_8/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_9/U4  ( .A(
        \pool/pool/pe_b_o_data[3][42] ), .B(
        \pool/pool/pe_b/peij_3_0/add/notb [9]), .Z(
        \pool/pool/pe_b/peij_3_0/add/fai_9/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_9/U3  ( .A(
        \pool/pool/pe_b/peij_3_0/add/cprop [9]), .B(
        \pool/pool/pe_b/peij_3_0/add/fai_9/n3 ), .Z(
        \pool/pool/pe_b/peij_3_0/d_acc [9]) );
  INV_X2 \pool/pool/pe_b/peij_3_0/add/fai_9/U2  ( .A(
        \pool/pool/pe_b/peij_3_0/add/fai_9/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_0/add/cprop [10]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_0/add/fai_9/U1  ( .A1(
        \pool/pool/pe_b/peij_3_0/add/notb [9]), .A2(
        \pool/pool/pe_b_o_data[3][42] ), .B1(
        \pool/pool/pe_b/peij_3_0/add/fai_9/n3 ), .B2(
        \pool/pool/pe_b/peij_3_0/add/cprop [9]), .ZN(
        \pool/pool/pe_b/peij_3_0/add/fai_9/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_10/U4  ( .A(
        \pool/pool/pe_b_o_data[3][43] ), .B(
        \pool/pool/pe_b/peij_3_0/add/notb [10]), .Z(
        \pool/pool/pe_b/peij_3_0/add/fai_10/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_0/add/fai_10/U3  ( .A(
        \pool/pool/pe_b/peij_3_0/add/cprop [10]), .B(
        \pool/pool/pe_b/peij_3_0/add/fai_10/n3 ), .Z(
        \pool/pool/pe_b/peij_3_0/d_acc [10]) );
  INV_X2 \pool/pool/pe_b/peij_3_0/add/fai_10/U2  ( .A(
        \pool/pool/pe_b/peij_3_0/add/fai_10/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_0/add/c_out ) );
  AOI22_X2 \pool/pool/pe_b/peij_3_0/add/fai_10/U1  ( .A1(
        \pool/pool/pe_b/peij_3_0/add/notb [10]), .A2(
        \pool/pool/pe_b_o_data[3][43] ), .B1(
        \pool/pool/pe_b/peij_3_0/add/fai_10/n3 ), .B2(
        \pool/pool/pe_b/peij_3_0/add/cprop [10]), .ZN(
        \pool/pool/pe_b/peij_3_0/add/fai_10/n1 ) );
  INV_X1 \pool/pool/pe_b/peij_3_1/U22  ( .A(\pool/pool/pe_b/n7 ), .ZN(
        \pool/pool/pe_b/peij_3_1/n16 ) );
  INV_X1 \pool/pool/pe_b/peij_3_1/U14  ( .A(\pool/pool/pe_b/n7 ), .ZN(
        \pool/pool/pe_b/peij_3_1/n12 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_1/U13  ( .A1(
        \pool/pool/pe_b/peij_3_1/d_acc [0]), .A2(\pool/pool/pe_b/peij_3_1/n18 ), .ZN(\pool/pool/pe_b/peij_3_1/n11 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_1/U12  ( .A1(
        \pool/pool/pe_b/peij_3_1/d_acc [1]), .A2(\pool/pool/pe_b/peij_3_1/n18 ), .ZN(\pool/pool/pe_b/peij_3_1/n10 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_1/U11  ( .A1(
        \pool/pool/pe_b/peij_3_1/d_acc [2]), .A2(\pool/pool/pe_b/peij_3_1/n18 ), .ZN(\pool/pool/pe_b/peij_3_1/n9 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_1/U10  ( .A1(
        \pool/pool/pe_b/peij_3_1/d_acc [3]), .A2(\pool/pool/pe_b/peij_3_1/n18 ), .ZN(\pool/pool/pe_b/peij_3_1/n8 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_1/U9  ( .A1(
        \pool/pool/pe_b/peij_3_1/d_acc [4]), .A2(\pool/pool/pe_b/peij_3_1/n18 ), .ZN(\pool/pool/pe_b/peij_3_1/n7 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_1/U8  ( .A1(
        \pool/pool/pe_b/peij_3_1/d_acc [5]), .A2(\pool/pool/pe_b/peij_3_1/n18 ), .ZN(\pool/pool/pe_b/peij_3_1/n6 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_1/U7  ( .A1(
        \pool/pool/pe_b/peij_3_1/d_acc [6]), .A2(\pool/pool/pe_b/peij_3_1/n18 ), .ZN(\pool/pool/pe_b/peij_3_1/n5 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_1/U6  ( .A1(
        \pool/pool/pe_b/peij_3_1/d_acc [7]), .A2(\pool/pool/pe_b/peij_3_1/n18 ), .ZN(\pool/pool/pe_b/peij_3_1/n4 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_1/U5  ( .A1(
        \pool/pool/pe_b/peij_3_1/d_acc [8]), .A2(\pool/pool/pe_b/peij_3_1/n18 ), .ZN(\pool/pool/pe_b/peij_3_1/n3 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_1/U4  ( .A1(
        \pool/pool/pe_b/peij_3_1/d_acc [9]), .A2(\pool/pool/pe_b/peij_3_1/n18 ), .ZN(\pool/pool/pe_b/peij_3_1/n2 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_1/U3  ( .A1(
        \pool/pool/pe_b/peij_3_1/d_acc [10]), .A2(
        \pool/pool/pe_b/peij_3_1/n18 ), .ZN(\pool/pool/pe_b/peij_3_1/n1 ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_1/q_acc_reg[10]  ( .D(
        \pool/pool/pe_b/peij_3_1/n1 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_1/n16 ), .Q(\pool/pool/pe_b_o_data[3][32] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_1/q_acc_reg[9]  ( .D(
        \pool/pool/pe_b/peij_3_1/n2 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_1/n16 ), .Q(\pool/pool/pe_b_o_data[3][31] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_1/q_acc_reg[8]  ( .D(
        \pool/pool/pe_b/peij_3_1/n3 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_1/n16 ), .Q(\pool/pool/pe_b_o_data[3][30] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_1/q_acc_reg[7]  ( .D(
        \pool/pool/pe_b/peij_3_1/n4 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_1/n16 ), .Q(\pool/pool/pe_b_o_data[3][29] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_1/q_acc_reg[6]  ( .D(
        \pool/pool/pe_b/peij_3_1/n5 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_1/n16 ), .Q(\pool/pool/pe_b_o_data[3][28] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_1/q_acc_reg[5]  ( .D(
        \pool/pool/pe_b/peij_3_1/n6 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_1/n16 ), .Q(\pool/pool/pe_b_o_data[3][27] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_1/q_acc_reg[4]  ( .D(
        \pool/pool/pe_b/peij_3_1/n7 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_1/n16 ), .Q(\pool/pool/pe_b_o_data[3][26] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_1/q_acc_reg[3]  ( .D(
        \pool/pool/pe_b/peij_3_1/n8 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_1/n16 ), .Q(\pool/pool/pe_b_o_data[3][25] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_1/q_acc_reg[2]  ( .D(
        \pool/pool/pe_b/peij_3_1/n9 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_1/n16 ), .Q(\pool/pool/pe_b_o_data[3][24] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_1/q_acc_reg[1]  ( .D(
        \pool/pool/pe_b/peij_3_1/n10 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_1/n16 ), .Q(\pool/pool/pe_b_o_data[3][23] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_1/q_acc_reg[0]  ( .D(
        \pool/pool/pe_b/peij_3_1/n11 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_1/n16 ), .Q(\pool/pool/pe_b_o_data[3][22] ) );
  INV_X2 \pool/pool/pe_b/peij_3_1/U21  ( .A(\pool/sync_clr ), .ZN(
        \pool/pool/pe_b/peij_3_1/n18 ) );
  AND3_X2 \pool/pool/pe_b/peij_3_1/U20  ( .A1(\pool/pool/pe_b/int_pe_en[3][1] ), .A2(\pool/pool/pe_b/peij_3_1/n18 ), .A3(1'b1), .ZN(
        \pool/pool/pe_b/peij_3_1/n17 ) );
  AND2_X2 \pool/pool/pe_b/peij_3_1/U19  ( .A1(\pool/pool/pe_b_i_data[3][8] ), 
        .A2(\pool/pool/pe_b/peij_3_1/n17 ), .ZN(\pool/pool/pe_b/peij_3_1/N33 )
         );
  AND2_X2 \pool/pool/pe_b/peij_3_1/U18  ( .A1(\pool/pool/pe_b_i_data[3][9] ), 
        .A2(\pool/pool/pe_b/peij_3_1/n17 ), .ZN(\pool/pool/pe_b/peij_3_1/N34 )
         );
  AND2_X2 \pool/pool/pe_b/peij_3_1/U17  ( .A1(\pool/pool/pe_b_i_data[3][10] ), 
        .A2(\pool/pool/pe_b/peij_3_1/n17 ), .ZN(\pool/pool/pe_b/peij_3_1/N35 )
         );
  AND4_X4 \pool/pool/pe_b/peij_3_1/U16  ( .A1(1'b1), .A2(
        \pool/pool/pe_b_i_data[3][11] ), .A3(\pool/pool/pe_b/int_pe_en[3][1] ), 
        .A4(\pool/pool/pe_b/peij_3_1/n18 ), .ZN(\pool/pool/pe_b/peij_3_1/N36 )
         );
  DFFR_X1 \pool/pool/pe_b/peij_3_1/q_im_reg[0]  ( .D(
        \pool/pool/pe_b/peij_3_1/N33 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_1/n12 ), .Q(\pool/pool/pe_b/peij_3_1/sgnext [0]) );
  DFFR_X1 \pool/pool/pe_b/peij_3_1/q_im_reg[1]  ( .D(
        \pool/pool/pe_b/peij_3_1/N34 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_1/n12 ), .Q(\pool/pool/pe_b/peij_3_1/sgnext [1]) );
  DFFR_X1 \pool/pool/pe_b/peij_3_1/q_im_reg[2]  ( .D(
        \pool/pool/pe_b/peij_3_1/N35 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_1/n12 ), .Q(\pool/pool/pe_b/peij_3_1/sgnext [2]) );
  DFFR_X1 \pool/pool/pe_b/peij_3_1/q_im_reg[3]  ( .D(
        \pool/pool/pe_b/peij_3_1/N36 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_1/n12 ), .Q(\pool/pool/pe_b/peij_3_1/sgnext_10 ) );
  SDFFR_X1 \pool/pool/pe_b/peij_3_1/q_k_reg  ( .D(1'b0), .SI(
        \pool/pool/pe_b/peij_3_1/n18 ), .SE(1'b0), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_1/n12 ), .Q(\pool/pool/pe_b/peij_3_1/q_k ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/U11  ( .A(
        \pool/pool/pe_b/peij_3_1/sgnext [0]), .B(\pool/pool/pe_b/peij_3_1/q_k ), .Z(\pool/pool/pe_b/peij_3_1/add/notb [0]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/U10  ( .A(
        \pool/pool/pe_b/peij_3_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_1/q_k ), .Z(\pool/pool/pe_b/peij_3_1/add/notb [10]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/U9  ( .A(
        \pool/pool/pe_b/peij_3_1/sgnext [1]), .B(\pool/pool/pe_b/peij_3_1/q_k ), .Z(\pool/pool/pe_b/peij_3_1/add/notb [1]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/U8  ( .A(
        \pool/pool/pe_b/peij_3_1/sgnext [2]), .B(\pool/pool/pe_b/peij_3_1/q_k ), .Z(\pool/pool/pe_b/peij_3_1/add/notb [2]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/U7  ( .A(
        \pool/pool/pe_b/peij_3_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_1/q_k ), .Z(\pool/pool/pe_b/peij_3_1/add/notb [3]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/U6  ( .A(
        \pool/pool/pe_b/peij_3_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_1/q_k ), .Z(\pool/pool/pe_b/peij_3_1/add/notb [4]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/U5  ( .A(
        \pool/pool/pe_b/peij_3_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_1/q_k ), .Z(\pool/pool/pe_b/peij_3_1/add/notb [5]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/U4  ( .A(
        \pool/pool/pe_b/peij_3_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_1/q_k ), .Z(\pool/pool/pe_b/peij_3_1/add/notb [6]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/U3  ( .A(
        \pool/pool/pe_b/peij_3_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_1/q_k ), .Z(\pool/pool/pe_b/peij_3_1/add/notb [7]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/U2  ( .A(
        \pool/pool/pe_b/peij_3_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_1/q_k ), .Z(\pool/pool/pe_b/peij_3_1/add/notb [8]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/U1  ( .A(
        \pool/pool/pe_b/peij_3_1/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_1/q_k ), .Z(\pool/pool/pe_b/peij_3_1/add/notb [9]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_0/U4  ( .A(
        \pool/pool/pe_b_o_data[3][22] ), .B(
        \pool/pool/pe_b/peij_3_1/add/notb [0]), .Z(
        \pool/pool/pe_b/peij_3_1/add/fai_0/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_0/U3  ( .A(
        \pool/pool/pe_b/peij_3_1/q_k ), .B(
        \pool/pool/pe_b/peij_3_1/add/fai_0/n3 ), .Z(
        \pool/pool/pe_b/peij_3_1/d_acc [0]) );
  INV_X2 \pool/pool/pe_b/peij_3_1/add/fai_0/U2  ( .A(
        \pool/pool/pe_b/peij_3_1/add/fai_0/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_1/add/cprop [1]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_1/add/fai_0/U1  ( .A1(
        \pool/pool/pe_b/peij_3_1/add/notb [0]), .A2(
        \pool/pool/pe_b_o_data[3][22] ), .B1(
        \pool/pool/pe_b/peij_3_1/add/fai_0/n3 ), .B2(
        \pool/pool/pe_b/peij_3_1/q_k ), .ZN(
        \pool/pool/pe_b/peij_3_1/add/fai_0/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_1/U4  ( .A(
        \pool/pool/pe_b_o_data[3][23] ), .B(
        \pool/pool/pe_b/peij_3_1/add/notb [1]), .Z(
        \pool/pool/pe_b/peij_3_1/add/fai_1/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_1/U3  ( .A(
        \pool/pool/pe_b/peij_3_1/add/cprop [1]), .B(
        \pool/pool/pe_b/peij_3_1/add/fai_1/n3 ), .Z(
        \pool/pool/pe_b/peij_3_1/d_acc [1]) );
  INV_X2 \pool/pool/pe_b/peij_3_1/add/fai_1/U2  ( .A(
        \pool/pool/pe_b/peij_3_1/add/fai_1/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_1/add/cprop [2]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_1/add/fai_1/U1  ( .A1(
        \pool/pool/pe_b/peij_3_1/add/notb [1]), .A2(
        \pool/pool/pe_b_o_data[3][23] ), .B1(
        \pool/pool/pe_b/peij_3_1/add/fai_1/n3 ), .B2(
        \pool/pool/pe_b/peij_3_1/add/cprop [1]), .ZN(
        \pool/pool/pe_b/peij_3_1/add/fai_1/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_2/U4  ( .A(
        \pool/pool/pe_b_o_data[3][24] ), .B(
        \pool/pool/pe_b/peij_3_1/add/notb [2]), .Z(
        \pool/pool/pe_b/peij_3_1/add/fai_2/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_2/U3  ( .A(
        \pool/pool/pe_b/peij_3_1/add/cprop [2]), .B(
        \pool/pool/pe_b/peij_3_1/add/fai_2/n3 ), .Z(
        \pool/pool/pe_b/peij_3_1/d_acc [2]) );
  INV_X2 \pool/pool/pe_b/peij_3_1/add/fai_2/U2  ( .A(
        \pool/pool/pe_b/peij_3_1/add/fai_2/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_1/add/cprop [3]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_1/add/fai_2/U1  ( .A1(
        \pool/pool/pe_b/peij_3_1/add/notb [2]), .A2(
        \pool/pool/pe_b_o_data[3][24] ), .B1(
        \pool/pool/pe_b/peij_3_1/add/fai_2/n3 ), .B2(
        \pool/pool/pe_b/peij_3_1/add/cprop [2]), .ZN(
        \pool/pool/pe_b/peij_3_1/add/fai_2/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_3/U4  ( .A(
        \pool/pool/pe_b_o_data[3][25] ), .B(
        \pool/pool/pe_b/peij_3_1/add/notb [3]), .Z(
        \pool/pool/pe_b/peij_3_1/add/fai_3/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_3/U3  ( .A(
        \pool/pool/pe_b/peij_3_1/add/cprop [3]), .B(
        \pool/pool/pe_b/peij_3_1/add/fai_3/n3 ), .Z(
        \pool/pool/pe_b/peij_3_1/d_acc [3]) );
  INV_X2 \pool/pool/pe_b/peij_3_1/add/fai_3/U2  ( .A(
        \pool/pool/pe_b/peij_3_1/add/fai_3/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_1/add/cprop [4]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_1/add/fai_3/U1  ( .A1(
        \pool/pool/pe_b/peij_3_1/add/notb [3]), .A2(
        \pool/pool/pe_b_o_data[3][25] ), .B1(
        \pool/pool/pe_b/peij_3_1/add/fai_3/n3 ), .B2(
        \pool/pool/pe_b/peij_3_1/add/cprop [3]), .ZN(
        \pool/pool/pe_b/peij_3_1/add/fai_3/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_4/U4  ( .A(
        \pool/pool/pe_b_o_data[3][26] ), .B(
        \pool/pool/pe_b/peij_3_1/add/notb [4]), .Z(
        \pool/pool/pe_b/peij_3_1/add/fai_4/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_4/U3  ( .A(
        \pool/pool/pe_b/peij_3_1/add/cprop [4]), .B(
        \pool/pool/pe_b/peij_3_1/add/fai_4/n3 ), .Z(
        \pool/pool/pe_b/peij_3_1/d_acc [4]) );
  INV_X2 \pool/pool/pe_b/peij_3_1/add/fai_4/U2  ( .A(
        \pool/pool/pe_b/peij_3_1/add/fai_4/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_1/add/cprop [5]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_1/add/fai_4/U1  ( .A1(
        \pool/pool/pe_b/peij_3_1/add/notb [4]), .A2(
        \pool/pool/pe_b_o_data[3][26] ), .B1(
        \pool/pool/pe_b/peij_3_1/add/fai_4/n3 ), .B2(
        \pool/pool/pe_b/peij_3_1/add/cprop [4]), .ZN(
        \pool/pool/pe_b/peij_3_1/add/fai_4/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_5/U4  ( .A(
        \pool/pool/pe_b_o_data[3][27] ), .B(
        \pool/pool/pe_b/peij_3_1/add/notb [5]), .Z(
        \pool/pool/pe_b/peij_3_1/add/fai_5/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_5/U3  ( .A(
        \pool/pool/pe_b/peij_3_1/add/cprop [5]), .B(
        \pool/pool/pe_b/peij_3_1/add/fai_5/n3 ), .Z(
        \pool/pool/pe_b/peij_3_1/d_acc [5]) );
  INV_X2 \pool/pool/pe_b/peij_3_1/add/fai_5/U2  ( .A(
        \pool/pool/pe_b/peij_3_1/add/fai_5/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_1/add/cprop [6]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_1/add/fai_5/U1  ( .A1(
        \pool/pool/pe_b/peij_3_1/add/notb [5]), .A2(
        \pool/pool/pe_b_o_data[3][27] ), .B1(
        \pool/pool/pe_b/peij_3_1/add/fai_5/n3 ), .B2(
        \pool/pool/pe_b/peij_3_1/add/cprop [5]), .ZN(
        \pool/pool/pe_b/peij_3_1/add/fai_5/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_6/U4  ( .A(
        \pool/pool/pe_b_o_data[3][28] ), .B(
        \pool/pool/pe_b/peij_3_1/add/notb [6]), .Z(
        \pool/pool/pe_b/peij_3_1/add/fai_6/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_6/U3  ( .A(
        \pool/pool/pe_b/peij_3_1/add/cprop [6]), .B(
        \pool/pool/pe_b/peij_3_1/add/fai_6/n3 ), .Z(
        \pool/pool/pe_b/peij_3_1/d_acc [6]) );
  INV_X2 \pool/pool/pe_b/peij_3_1/add/fai_6/U2  ( .A(
        \pool/pool/pe_b/peij_3_1/add/fai_6/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_1/add/cprop [7]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_1/add/fai_6/U1  ( .A1(
        \pool/pool/pe_b/peij_3_1/add/notb [6]), .A2(
        \pool/pool/pe_b_o_data[3][28] ), .B1(
        \pool/pool/pe_b/peij_3_1/add/fai_6/n3 ), .B2(
        \pool/pool/pe_b/peij_3_1/add/cprop [6]), .ZN(
        \pool/pool/pe_b/peij_3_1/add/fai_6/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_7/U4  ( .A(
        \pool/pool/pe_b_o_data[3][29] ), .B(
        \pool/pool/pe_b/peij_3_1/add/notb [7]), .Z(
        \pool/pool/pe_b/peij_3_1/add/fai_7/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_7/U3  ( .A(
        \pool/pool/pe_b/peij_3_1/add/cprop [7]), .B(
        \pool/pool/pe_b/peij_3_1/add/fai_7/n3 ), .Z(
        \pool/pool/pe_b/peij_3_1/d_acc [7]) );
  INV_X2 \pool/pool/pe_b/peij_3_1/add/fai_7/U2  ( .A(
        \pool/pool/pe_b/peij_3_1/add/fai_7/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_1/add/cprop [8]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_1/add/fai_7/U1  ( .A1(
        \pool/pool/pe_b/peij_3_1/add/notb [7]), .A2(
        \pool/pool/pe_b_o_data[3][29] ), .B1(
        \pool/pool/pe_b/peij_3_1/add/fai_7/n3 ), .B2(
        \pool/pool/pe_b/peij_3_1/add/cprop [7]), .ZN(
        \pool/pool/pe_b/peij_3_1/add/fai_7/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_8/U4  ( .A(
        \pool/pool/pe_b_o_data[3][30] ), .B(
        \pool/pool/pe_b/peij_3_1/add/notb [8]), .Z(
        \pool/pool/pe_b/peij_3_1/add/fai_8/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_8/U3  ( .A(
        \pool/pool/pe_b/peij_3_1/add/cprop [8]), .B(
        \pool/pool/pe_b/peij_3_1/add/fai_8/n3 ), .Z(
        \pool/pool/pe_b/peij_3_1/d_acc [8]) );
  INV_X2 \pool/pool/pe_b/peij_3_1/add/fai_8/U2  ( .A(
        \pool/pool/pe_b/peij_3_1/add/fai_8/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_1/add/cprop [9]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_1/add/fai_8/U1  ( .A1(
        \pool/pool/pe_b/peij_3_1/add/notb [8]), .A2(
        \pool/pool/pe_b_o_data[3][30] ), .B1(
        \pool/pool/pe_b/peij_3_1/add/fai_8/n3 ), .B2(
        \pool/pool/pe_b/peij_3_1/add/cprop [8]), .ZN(
        \pool/pool/pe_b/peij_3_1/add/fai_8/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_9/U4  ( .A(
        \pool/pool/pe_b_o_data[3][31] ), .B(
        \pool/pool/pe_b/peij_3_1/add/notb [9]), .Z(
        \pool/pool/pe_b/peij_3_1/add/fai_9/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_9/U3  ( .A(
        \pool/pool/pe_b/peij_3_1/add/cprop [9]), .B(
        \pool/pool/pe_b/peij_3_1/add/fai_9/n3 ), .Z(
        \pool/pool/pe_b/peij_3_1/d_acc [9]) );
  INV_X2 \pool/pool/pe_b/peij_3_1/add/fai_9/U2  ( .A(
        \pool/pool/pe_b/peij_3_1/add/fai_9/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_1/add/cprop [10]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_1/add/fai_9/U1  ( .A1(
        \pool/pool/pe_b/peij_3_1/add/notb [9]), .A2(
        \pool/pool/pe_b_o_data[3][31] ), .B1(
        \pool/pool/pe_b/peij_3_1/add/fai_9/n3 ), .B2(
        \pool/pool/pe_b/peij_3_1/add/cprop [9]), .ZN(
        \pool/pool/pe_b/peij_3_1/add/fai_9/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_10/U4  ( .A(
        \pool/pool/pe_b_o_data[3][32] ), .B(
        \pool/pool/pe_b/peij_3_1/add/notb [10]), .Z(
        \pool/pool/pe_b/peij_3_1/add/fai_10/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_1/add/fai_10/U3  ( .A(
        \pool/pool/pe_b/peij_3_1/add/cprop [10]), .B(
        \pool/pool/pe_b/peij_3_1/add/fai_10/n3 ), .Z(
        \pool/pool/pe_b/peij_3_1/d_acc [10]) );
  INV_X2 \pool/pool/pe_b/peij_3_1/add/fai_10/U2  ( .A(
        \pool/pool/pe_b/peij_3_1/add/fai_10/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_1/add/c_out ) );
  AOI22_X2 \pool/pool/pe_b/peij_3_1/add/fai_10/U1  ( .A1(
        \pool/pool/pe_b/peij_3_1/add/notb [10]), .A2(
        \pool/pool/pe_b_o_data[3][32] ), .B1(
        \pool/pool/pe_b/peij_3_1/add/fai_10/n3 ), .B2(
        \pool/pool/pe_b/peij_3_1/add/cprop [10]), .ZN(
        \pool/pool/pe_b/peij_3_1/add/fai_10/n1 ) );
  INV_X1 \pool/pool/pe_b/peij_3_2/U22  ( .A(\pool/pool/pe_b/n7 ), .ZN(
        \pool/pool/pe_b/peij_3_2/n17 ) );
  INV_X1 \pool/pool/pe_b/peij_3_2/U17  ( .A(\pool/pool/pe_b/n7 ), .ZN(
        \pool/pool/pe_b/peij_3_2/n16 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_2/U14  ( .A1(
        \pool/pool/pe_b/peij_3_2/d_acc [0]), .A2(\pool/pool/pe_b/peij_3_2/n19 ), .ZN(\pool/pool/pe_b/peij_3_2/n12 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_2/U13  ( .A1(
        \pool/pool/pe_b/peij_3_2/d_acc [1]), .A2(\pool/pool/pe_b/peij_3_2/n19 ), .ZN(\pool/pool/pe_b/peij_3_2/n11 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_2/U12  ( .A1(
        \pool/pool/pe_b/peij_3_2/d_acc [2]), .A2(\pool/pool/pe_b/peij_3_2/n19 ), .ZN(\pool/pool/pe_b/peij_3_2/n10 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_2/U11  ( .A1(
        \pool/pool/pe_b/peij_3_2/d_acc [3]), .A2(\pool/pool/pe_b/peij_3_2/n19 ), .ZN(\pool/pool/pe_b/peij_3_2/n9 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_2/U10  ( .A1(
        \pool/pool/pe_b/peij_3_2/d_acc [4]), .A2(\pool/pool/pe_b/peij_3_2/n19 ), .ZN(\pool/pool/pe_b/peij_3_2/n8 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_2/U9  ( .A1(
        \pool/pool/pe_b/peij_3_2/d_acc [5]), .A2(\pool/pool/pe_b/peij_3_2/n19 ), .ZN(\pool/pool/pe_b/peij_3_2/n7 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_2/U8  ( .A1(
        \pool/pool/pe_b/peij_3_2/d_acc [6]), .A2(\pool/pool/pe_b/peij_3_2/n19 ), .ZN(\pool/pool/pe_b/peij_3_2/n6 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_2/U7  ( .A1(
        \pool/pool/pe_b/peij_3_2/d_acc [7]), .A2(\pool/pool/pe_b/peij_3_2/n19 ), .ZN(\pool/pool/pe_b/peij_3_2/n5 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_2/U6  ( .A1(
        \pool/pool/pe_b/peij_3_2/d_acc [8]), .A2(\pool/pool/pe_b/peij_3_2/n19 ), .ZN(\pool/pool/pe_b/peij_3_2/n4 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_2/U5  ( .A1(
        \pool/pool/pe_b/peij_3_2/d_acc [9]), .A2(\pool/pool/pe_b/peij_3_2/n19 ), .ZN(\pool/pool/pe_b/peij_3_2/n3 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_2/U4  ( .A1(
        \pool/pool/pe_b/peij_3_2/d_acc [10]), .A2(
        \pool/pool/pe_b/peij_3_2/n19 ), .ZN(\pool/pool/pe_b/peij_3_2/n2 ) );
  SDFFR_X1 \pool/pool/pe_b/peij_3_2/q_im_reg[2]  ( .D(1'b0), .SI(
        \pool/pool/pe_b/peij_3_2/n18 ), .SE(\pool/pool/pe_b_i_data[3][6] ), 
        .CK(clk), .RN(\pool/pool/pe_b/peij_3_2/n17 ), .Q(
        \pool/pool/pe_b/peij_3_2/sgnext [2]) );
  DFFR_X1 \pool/pool/pe_b/peij_3_2/q_acc_reg[10]  ( .D(
        \pool/pool/pe_b/peij_3_2/n2 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_2/n17 ), .Q(\pool/pool/pe_b_o_data[3][21] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_2/q_acc_reg[9]  ( .D(
        \pool/pool/pe_b/peij_3_2/n3 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_2/n17 ), .Q(\pool/pool/pe_b_o_data[3][20] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_2/q_acc_reg[8]  ( .D(
        \pool/pool/pe_b/peij_3_2/n4 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_2/n17 ), .Q(\pool/pool/pe_b_o_data[3][19] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_2/q_acc_reg[7]  ( .D(
        \pool/pool/pe_b/peij_3_2/n5 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_2/n17 ), .Q(\pool/pool/pe_b_o_data[3][18] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_2/q_acc_reg[6]  ( .D(
        \pool/pool/pe_b/peij_3_2/n6 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_2/n17 ), .Q(\pool/pool/pe_b_o_data[3][17] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_2/q_acc_reg[5]  ( .D(
        \pool/pool/pe_b/peij_3_2/n7 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_2/n17 ), .Q(\pool/pool/pe_b_o_data[3][16] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_2/q_acc_reg[4]  ( .D(
        \pool/pool/pe_b/peij_3_2/n8 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_2/n17 ), .Q(\pool/pool/pe_b_o_data[3][15] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_2/q_acc_reg[3]  ( .D(
        \pool/pool/pe_b/peij_3_2/n9 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_2/n17 ), .Q(\pool/pool/pe_b_o_data[3][14] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_2/q_acc_reg[2]  ( .D(
        \pool/pool/pe_b/peij_3_2/n10 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_2/n17 ), .Q(\pool/pool/pe_b_o_data[3][13] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_2/q_acc_reg[1]  ( .D(
        \pool/pool/pe_b/peij_3_2/n11 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_2/n17 ), .Q(\pool/pool/pe_b_o_data[3][12] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_2/q_acc_reg[0]  ( .D(
        \pool/pool/pe_b/peij_3_2/n12 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_2/n17 ), .Q(\pool/pool/pe_b_o_data[3][11] ) );
  INV_X2 \pool/pool/pe_b/peij_3_2/U21  ( .A(\pool/sync_clr ), .ZN(
        \pool/pool/pe_b/peij_3_2/n19 ) );
  AND3_X2 \pool/pool/pe_b/peij_3_2/U20  ( .A1(\pool/pool/pe_b/int_pe_en[3][2] ), .A2(\pool/pool/pe_b/peij_3_2/n19 ), .A3(1'b1), .ZN(
        \pool/pool/pe_b/peij_3_2/n18 ) );
  AND2_X2 \pool/pool/pe_b/peij_3_2/U19  ( .A1(\pool/pool/pe_b_i_data[3][4] ), 
        .A2(\pool/pool/pe_b/peij_3_2/n18 ), .ZN(\pool/pool/pe_b/peij_3_2/N33 )
         );
  AND2_X2 \pool/pool/pe_b/peij_3_2/U18  ( .A1(\pool/pool/pe_b_i_data[3][5] ), 
        .A2(\pool/pool/pe_b/peij_3_2/n18 ), .ZN(\pool/pool/pe_b/peij_3_2/N34 )
         );
  AND4_X4 \pool/pool/pe_b/peij_3_2/U16  ( .A1(1'b1), .A2(
        \pool/pool/pe_b_i_data[3][7] ), .A3(\pool/pool/pe_b/int_pe_en[3][2] ), 
        .A4(\pool/pool/pe_b/peij_3_2/n19 ), .ZN(\pool/pool/pe_b/peij_3_2/N36 )
         );
  DFFR_X1 \pool/pool/pe_b/peij_3_2/q_im_reg[0]  ( .D(
        \pool/pool/pe_b/peij_3_2/N33 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_2/n16 ), .Q(\pool/pool/pe_b/peij_3_2/sgnext [0]) );
  DFFR_X1 \pool/pool/pe_b/peij_3_2/q_im_reg[1]  ( .D(
        \pool/pool/pe_b/peij_3_2/N34 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_2/n16 ), .Q(\pool/pool/pe_b/peij_3_2/sgnext [1]) );
  DFFR_X1 \pool/pool/pe_b/peij_3_2/q_im_reg[3]  ( .D(
        \pool/pool/pe_b/peij_3_2/N36 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_2/n16 ), .Q(\pool/pool/pe_b/peij_3_2/sgnext_10 ) );
  SDFFR_X1 \pool/pool/pe_b/peij_3_2/q_k_reg  ( .D(1'b0), .SI(
        \pool/pool/pe_b/peij_3_2/n19 ), .SE(1'b0), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_2/n16 ), .Q(\pool/pool/pe_b/peij_3_2/q_k ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/U11  ( .A(
        \pool/pool/pe_b/peij_3_2/sgnext [0]), .B(\pool/pool/pe_b/peij_3_2/q_k ), .Z(\pool/pool/pe_b/peij_3_2/add/notb [0]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/U10  ( .A(
        \pool/pool/pe_b/peij_3_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_2/q_k ), .Z(\pool/pool/pe_b/peij_3_2/add/notb [10]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/U9  ( .A(
        \pool/pool/pe_b/peij_3_2/sgnext [1]), .B(\pool/pool/pe_b/peij_3_2/q_k ), .Z(\pool/pool/pe_b/peij_3_2/add/notb [1]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/U8  ( .A(
        \pool/pool/pe_b/peij_3_2/sgnext [2]), .B(\pool/pool/pe_b/peij_3_2/q_k ), .Z(\pool/pool/pe_b/peij_3_2/add/notb [2]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/U7  ( .A(
        \pool/pool/pe_b/peij_3_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_2/q_k ), .Z(\pool/pool/pe_b/peij_3_2/add/notb [3]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/U6  ( .A(
        \pool/pool/pe_b/peij_3_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_2/q_k ), .Z(\pool/pool/pe_b/peij_3_2/add/notb [4]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/U5  ( .A(
        \pool/pool/pe_b/peij_3_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_2/q_k ), .Z(\pool/pool/pe_b/peij_3_2/add/notb [5]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/U4  ( .A(
        \pool/pool/pe_b/peij_3_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_2/q_k ), .Z(\pool/pool/pe_b/peij_3_2/add/notb [6]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/U3  ( .A(
        \pool/pool/pe_b/peij_3_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_2/q_k ), .Z(\pool/pool/pe_b/peij_3_2/add/notb [7]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/U2  ( .A(
        \pool/pool/pe_b/peij_3_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_2/q_k ), .Z(\pool/pool/pe_b/peij_3_2/add/notb [8]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/U1  ( .A(
        \pool/pool/pe_b/peij_3_2/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_2/q_k ), .Z(\pool/pool/pe_b/peij_3_2/add/notb [9]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_0/U4  ( .A(
        \pool/pool/pe_b_o_data[3][11] ), .B(
        \pool/pool/pe_b/peij_3_2/add/notb [0]), .Z(
        \pool/pool/pe_b/peij_3_2/add/fai_0/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_0/U3  ( .A(
        \pool/pool/pe_b/peij_3_2/q_k ), .B(
        \pool/pool/pe_b/peij_3_2/add/fai_0/n3 ), .Z(
        \pool/pool/pe_b/peij_3_2/d_acc [0]) );
  INV_X2 \pool/pool/pe_b/peij_3_2/add/fai_0/U2  ( .A(
        \pool/pool/pe_b/peij_3_2/add/fai_0/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_2/add/cprop [1]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_2/add/fai_0/U1  ( .A1(
        \pool/pool/pe_b/peij_3_2/add/notb [0]), .A2(
        \pool/pool/pe_b_o_data[3][11] ), .B1(
        \pool/pool/pe_b/peij_3_2/add/fai_0/n3 ), .B2(
        \pool/pool/pe_b/peij_3_2/q_k ), .ZN(
        \pool/pool/pe_b/peij_3_2/add/fai_0/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_1/U4  ( .A(
        \pool/pool/pe_b_o_data[3][12] ), .B(
        \pool/pool/pe_b/peij_3_2/add/notb [1]), .Z(
        \pool/pool/pe_b/peij_3_2/add/fai_1/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_1/U3  ( .A(
        \pool/pool/pe_b/peij_3_2/add/cprop [1]), .B(
        \pool/pool/pe_b/peij_3_2/add/fai_1/n3 ), .Z(
        \pool/pool/pe_b/peij_3_2/d_acc [1]) );
  INV_X2 \pool/pool/pe_b/peij_3_2/add/fai_1/U2  ( .A(
        \pool/pool/pe_b/peij_3_2/add/fai_1/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_2/add/cprop [2]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_2/add/fai_1/U1  ( .A1(
        \pool/pool/pe_b/peij_3_2/add/notb [1]), .A2(
        \pool/pool/pe_b_o_data[3][12] ), .B1(
        \pool/pool/pe_b/peij_3_2/add/fai_1/n3 ), .B2(
        \pool/pool/pe_b/peij_3_2/add/cprop [1]), .ZN(
        \pool/pool/pe_b/peij_3_2/add/fai_1/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_2/U4  ( .A(
        \pool/pool/pe_b_o_data[3][13] ), .B(
        \pool/pool/pe_b/peij_3_2/add/notb [2]), .Z(
        \pool/pool/pe_b/peij_3_2/add/fai_2/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_2/U3  ( .A(
        \pool/pool/pe_b/peij_3_2/add/cprop [2]), .B(
        \pool/pool/pe_b/peij_3_2/add/fai_2/n3 ), .Z(
        \pool/pool/pe_b/peij_3_2/d_acc [2]) );
  INV_X2 \pool/pool/pe_b/peij_3_2/add/fai_2/U2  ( .A(
        \pool/pool/pe_b/peij_3_2/add/fai_2/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_2/add/cprop [3]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_2/add/fai_2/U1  ( .A1(
        \pool/pool/pe_b/peij_3_2/add/notb [2]), .A2(
        \pool/pool/pe_b_o_data[3][13] ), .B1(
        \pool/pool/pe_b/peij_3_2/add/fai_2/n3 ), .B2(
        \pool/pool/pe_b/peij_3_2/add/cprop [2]), .ZN(
        \pool/pool/pe_b/peij_3_2/add/fai_2/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_3/U4  ( .A(
        \pool/pool/pe_b_o_data[3][14] ), .B(
        \pool/pool/pe_b/peij_3_2/add/notb [3]), .Z(
        \pool/pool/pe_b/peij_3_2/add/fai_3/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_3/U3  ( .A(
        \pool/pool/pe_b/peij_3_2/add/cprop [3]), .B(
        \pool/pool/pe_b/peij_3_2/add/fai_3/n3 ), .Z(
        \pool/pool/pe_b/peij_3_2/d_acc [3]) );
  INV_X2 \pool/pool/pe_b/peij_3_2/add/fai_3/U2  ( .A(
        \pool/pool/pe_b/peij_3_2/add/fai_3/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_2/add/cprop [4]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_2/add/fai_3/U1  ( .A1(
        \pool/pool/pe_b/peij_3_2/add/notb [3]), .A2(
        \pool/pool/pe_b_o_data[3][14] ), .B1(
        \pool/pool/pe_b/peij_3_2/add/fai_3/n3 ), .B2(
        \pool/pool/pe_b/peij_3_2/add/cprop [3]), .ZN(
        \pool/pool/pe_b/peij_3_2/add/fai_3/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_4/U4  ( .A(
        \pool/pool/pe_b_o_data[3][15] ), .B(
        \pool/pool/pe_b/peij_3_2/add/notb [4]), .Z(
        \pool/pool/pe_b/peij_3_2/add/fai_4/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_4/U3  ( .A(
        \pool/pool/pe_b/peij_3_2/add/cprop [4]), .B(
        \pool/pool/pe_b/peij_3_2/add/fai_4/n3 ), .Z(
        \pool/pool/pe_b/peij_3_2/d_acc [4]) );
  INV_X2 \pool/pool/pe_b/peij_3_2/add/fai_4/U2  ( .A(
        \pool/pool/pe_b/peij_3_2/add/fai_4/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_2/add/cprop [5]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_2/add/fai_4/U1  ( .A1(
        \pool/pool/pe_b/peij_3_2/add/notb [4]), .A2(
        \pool/pool/pe_b_o_data[3][15] ), .B1(
        \pool/pool/pe_b/peij_3_2/add/fai_4/n3 ), .B2(
        \pool/pool/pe_b/peij_3_2/add/cprop [4]), .ZN(
        \pool/pool/pe_b/peij_3_2/add/fai_4/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_5/U4  ( .A(
        \pool/pool/pe_b_o_data[3][16] ), .B(
        \pool/pool/pe_b/peij_3_2/add/notb [5]), .Z(
        \pool/pool/pe_b/peij_3_2/add/fai_5/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_5/U3  ( .A(
        \pool/pool/pe_b/peij_3_2/add/cprop [5]), .B(
        \pool/pool/pe_b/peij_3_2/add/fai_5/n3 ), .Z(
        \pool/pool/pe_b/peij_3_2/d_acc [5]) );
  INV_X2 \pool/pool/pe_b/peij_3_2/add/fai_5/U2  ( .A(
        \pool/pool/pe_b/peij_3_2/add/fai_5/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_2/add/cprop [6]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_2/add/fai_5/U1  ( .A1(
        \pool/pool/pe_b/peij_3_2/add/notb [5]), .A2(
        \pool/pool/pe_b_o_data[3][16] ), .B1(
        \pool/pool/pe_b/peij_3_2/add/fai_5/n3 ), .B2(
        \pool/pool/pe_b/peij_3_2/add/cprop [5]), .ZN(
        \pool/pool/pe_b/peij_3_2/add/fai_5/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_6/U4  ( .A(
        \pool/pool/pe_b_o_data[3][17] ), .B(
        \pool/pool/pe_b/peij_3_2/add/notb [6]), .Z(
        \pool/pool/pe_b/peij_3_2/add/fai_6/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_6/U3  ( .A(
        \pool/pool/pe_b/peij_3_2/add/cprop [6]), .B(
        \pool/pool/pe_b/peij_3_2/add/fai_6/n3 ), .Z(
        \pool/pool/pe_b/peij_3_2/d_acc [6]) );
  INV_X2 \pool/pool/pe_b/peij_3_2/add/fai_6/U2  ( .A(
        \pool/pool/pe_b/peij_3_2/add/fai_6/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_2/add/cprop [7]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_2/add/fai_6/U1  ( .A1(
        \pool/pool/pe_b/peij_3_2/add/notb [6]), .A2(
        \pool/pool/pe_b_o_data[3][17] ), .B1(
        \pool/pool/pe_b/peij_3_2/add/fai_6/n3 ), .B2(
        \pool/pool/pe_b/peij_3_2/add/cprop [6]), .ZN(
        \pool/pool/pe_b/peij_3_2/add/fai_6/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_7/U4  ( .A(
        \pool/pool/pe_b_o_data[3][18] ), .B(
        \pool/pool/pe_b/peij_3_2/add/notb [7]), .Z(
        \pool/pool/pe_b/peij_3_2/add/fai_7/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_7/U3  ( .A(
        \pool/pool/pe_b/peij_3_2/add/cprop [7]), .B(
        \pool/pool/pe_b/peij_3_2/add/fai_7/n3 ), .Z(
        \pool/pool/pe_b/peij_3_2/d_acc [7]) );
  INV_X2 \pool/pool/pe_b/peij_3_2/add/fai_7/U2  ( .A(
        \pool/pool/pe_b/peij_3_2/add/fai_7/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_2/add/cprop [8]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_2/add/fai_7/U1  ( .A1(
        \pool/pool/pe_b/peij_3_2/add/notb [7]), .A2(
        \pool/pool/pe_b_o_data[3][18] ), .B1(
        \pool/pool/pe_b/peij_3_2/add/fai_7/n3 ), .B2(
        \pool/pool/pe_b/peij_3_2/add/cprop [7]), .ZN(
        \pool/pool/pe_b/peij_3_2/add/fai_7/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_8/U4  ( .A(
        \pool/pool/pe_b_o_data[3][19] ), .B(
        \pool/pool/pe_b/peij_3_2/add/notb [8]), .Z(
        \pool/pool/pe_b/peij_3_2/add/fai_8/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_8/U3  ( .A(
        \pool/pool/pe_b/peij_3_2/add/cprop [8]), .B(
        \pool/pool/pe_b/peij_3_2/add/fai_8/n3 ), .Z(
        \pool/pool/pe_b/peij_3_2/d_acc [8]) );
  INV_X2 \pool/pool/pe_b/peij_3_2/add/fai_8/U2  ( .A(
        \pool/pool/pe_b/peij_3_2/add/fai_8/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_2/add/cprop [9]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_2/add/fai_8/U1  ( .A1(
        \pool/pool/pe_b/peij_3_2/add/notb [8]), .A2(
        \pool/pool/pe_b_o_data[3][19] ), .B1(
        \pool/pool/pe_b/peij_3_2/add/fai_8/n3 ), .B2(
        \pool/pool/pe_b/peij_3_2/add/cprop [8]), .ZN(
        \pool/pool/pe_b/peij_3_2/add/fai_8/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_9/U4  ( .A(
        \pool/pool/pe_b_o_data[3][20] ), .B(
        \pool/pool/pe_b/peij_3_2/add/notb [9]), .Z(
        \pool/pool/pe_b/peij_3_2/add/fai_9/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_9/U3  ( .A(
        \pool/pool/pe_b/peij_3_2/add/cprop [9]), .B(
        \pool/pool/pe_b/peij_3_2/add/fai_9/n3 ), .Z(
        \pool/pool/pe_b/peij_3_2/d_acc [9]) );
  INV_X2 \pool/pool/pe_b/peij_3_2/add/fai_9/U2  ( .A(
        \pool/pool/pe_b/peij_3_2/add/fai_9/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_2/add/cprop [10]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_2/add/fai_9/U1  ( .A1(
        \pool/pool/pe_b/peij_3_2/add/notb [9]), .A2(
        \pool/pool/pe_b_o_data[3][20] ), .B1(
        \pool/pool/pe_b/peij_3_2/add/fai_9/n3 ), .B2(
        \pool/pool/pe_b/peij_3_2/add/cprop [9]), .ZN(
        \pool/pool/pe_b/peij_3_2/add/fai_9/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_10/U4  ( .A(
        \pool/pool/pe_b_o_data[3][21] ), .B(
        \pool/pool/pe_b/peij_3_2/add/notb [10]), .Z(
        \pool/pool/pe_b/peij_3_2/add/fai_10/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_2/add/fai_10/U3  ( .A(
        \pool/pool/pe_b/peij_3_2/add/cprop [10]), .B(
        \pool/pool/pe_b/peij_3_2/add/fai_10/n3 ), .Z(
        \pool/pool/pe_b/peij_3_2/d_acc [10]) );
  INV_X2 \pool/pool/pe_b/peij_3_2/add/fai_10/U2  ( .A(
        \pool/pool/pe_b/peij_3_2/add/fai_10/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_2/add/c_out ) );
  AOI22_X2 \pool/pool/pe_b/peij_3_2/add/fai_10/U1  ( .A1(
        \pool/pool/pe_b/peij_3_2/add/notb [10]), .A2(
        \pool/pool/pe_b_o_data[3][21] ), .B1(
        \pool/pool/pe_b/peij_3_2/add/fai_10/n3 ), .B2(
        \pool/pool/pe_b/peij_3_2/add/cprop [10]), .ZN(
        \pool/pool/pe_b/peij_3_2/add/fai_10/n1 ) );
  INV_X1 \pool/pool/pe_b/peij_3_3/U22  ( .A(\pool/pool/pe_b/n7 ), .ZN(
        \pool/pool/pe_b/peij_3_3/n16 ) );
  INV_X1 \pool/pool/pe_b/peij_3_3/U14  ( .A(\pool/pool/pe_b/n7 ), .ZN(
        \pool/pool/pe_b/peij_3_3/n12 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_3/U13  ( .A1(
        \pool/pool/pe_b/peij_3_3/d_acc [0]), .A2(\pool/pool/pe_b/peij_3_3/n18 ), .ZN(\pool/pool/pe_b/peij_3_3/n11 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_3/U12  ( .A1(
        \pool/pool/pe_b/peij_3_3/d_acc [1]), .A2(\pool/pool/pe_b/peij_3_3/n18 ), .ZN(\pool/pool/pe_b/peij_3_3/n10 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_3/U11  ( .A1(
        \pool/pool/pe_b/peij_3_3/d_acc [2]), .A2(\pool/pool/pe_b/peij_3_3/n18 ), .ZN(\pool/pool/pe_b/peij_3_3/n9 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_3/U10  ( .A1(
        \pool/pool/pe_b/peij_3_3/d_acc [3]), .A2(\pool/pool/pe_b/peij_3_3/n18 ), .ZN(\pool/pool/pe_b/peij_3_3/n8 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_3/U9  ( .A1(
        \pool/pool/pe_b/peij_3_3/d_acc [4]), .A2(\pool/pool/pe_b/peij_3_3/n18 ), .ZN(\pool/pool/pe_b/peij_3_3/n7 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_3/U8  ( .A1(
        \pool/pool/pe_b/peij_3_3/d_acc [5]), .A2(\pool/pool/pe_b/peij_3_3/n18 ), .ZN(\pool/pool/pe_b/peij_3_3/n6 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_3/U7  ( .A1(
        \pool/pool/pe_b/peij_3_3/d_acc [6]), .A2(\pool/pool/pe_b/peij_3_3/n18 ), .ZN(\pool/pool/pe_b/peij_3_3/n5 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_3/U6  ( .A1(
        \pool/pool/pe_b/peij_3_3/d_acc [7]), .A2(\pool/pool/pe_b/peij_3_3/n18 ), .ZN(\pool/pool/pe_b/peij_3_3/n4 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_3/U5  ( .A1(
        \pool/pool/pe_b/peij_3_3/d_acc [8]), .A2(\pool/pool/pe_b/peij_3_3/n18 ), .ZN(\pool/pool/pe_b/peij_3_3/n3 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_3/U4  ( .A1(
        \pool/pool/pe_b/peij_3_3/d_acc [9]), .A2(\pool/pool/pe_b/peij_3_3/n18 ), .ZN(\pool/pool/pe_b/peij_3_3/n2 ) );
  AND2_X1 \pool/pool/pe_b/peij_3_3/U3  ( .A1(
        \pool/pool/pe_b/peij_3_3/d_acc [10]), .A2(
        \pool/pool/pe_b/peij_3_3/n18 ), .ZN(\pool/pool/pe_b/peij_3_3/n1 ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_3/q_acc_reg[10]  ( .D(
        \pool/pool/pe_b/peij_3_3/n1 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_3/n16 ), .Q(\pool/pool/pe_b_o_data[3][10] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_3/q_acc_reg[9]  ( .D(
        \pool/pool/pe_b/peij_3_3/n2 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_3/n16 ), .Q(\pool/pool/pe_b_o_data[3][9] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_3/q_acc_reg[8]  ( .D(
        \pool/pool/pe_b/peij_3_3/n3 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_3/n16 ), .Q(\pool/pool/pe_b_o_data[3][8] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_3/q_acc_reg[7]  ( .D(
        \pool/pool/pe_b/peij_3_3/n4 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_3/n16 ), .Q(\pool/pool/pe_b_o_data[3][7] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_3/q_acc_reg[6]  ( .D(
        \pool/pool/pe_b/peij_3_3/n5 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_3/n16 ), .Q(\pool/pool/pe_b_o_data[3][6] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_3/q_acc_reg[5]  ( .D(
        \pool/pool/pe_b/peij_3_3/n6 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_3/n16 ), .Q(\pool/pool/pe_b_o_data[3][5] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_3/q_acc_reg[4]  ( .D(
        \pool/pool/pe_b/peij_3_3/n7 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_3/n16 ), .Q(\pool/pool/pe_b_o_data[3][4] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_3/q_acc_reg[3]  ( .D(
        \pool/pool/pe_b/peij_3_3/n8 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_3/n16 ), .Q(\pool/pool/pe_b_o_data[3][3] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_3/q_acc_reg[2]  ( .D(
        \pool/pool/pe_b/peij_3_3/n9 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_3/n16 ), .Q(\pool/pool/pe_b_o_data[3][2] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_3/q_acc_reg[1]  ( .D(
        \pool/pool/pe_b/peij_3_3/n10 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_3/n16 ), .Q(\pool/pool/pe_b_o_data[3][1] ) );
  DFFR_X1 \pool/pool/pe_b/peij_3_3/q_acc_reg[0]  ( .D(
        \pool/pool/pe_b/peij_3_3/n11 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_3/n16 ), .Q(\pool/pool/pe_b_o_data[3][0] ) );
  INV_X2 \pool/pool/pe_b/peij_3_3/U21  ( .A(\pool/sync_clr ), .ZN(
        \pool/pool/pe_b/peij_3_3/n18 ) );
  AND3_X2 \pool/pool/pe_b/peij_3_3/U20  ( .A1(\pool/pool/pe_b/int_pe_en[3][3] ), .A2(\pool/pool/pe_b/peij_3_3/n18 ), .A3(1'b1), .ZN(
        \pool/pool/pe_b/peij_3_3/n17 ) );
  AND2_X2 \pool/pool/pe_b/peij_3_3/U19  ( .A1(\pool/pool/pe_b_i_data[3][0] ), 
        .A2(\pool/pool/pe_b/peij_3_3/n17 ), .ZN(\pool/pool/pe_b/peij_3_3/N33 )
         );
  AND2_X2 \pool/pool/pe_b/peij_3_3/U18  ( .A1(\pool/pool/pe_b_i_data[3][1] ), 
        .A2(\pool/pool/pe_b/peij_3_3/n17 ), .ZN(\pool/pool/pe_b/peij_3_3/N34 )
         );
  AND2_X2 \pool/pool/pe_b/peij_3_3/U17  ( .A1(\pool/pool/pe_b_i_data[3][2] ), 
        .A2(\pool/pool/pe_b/peij_3_3/n17 ), .ZN(\pool/pool/pe_b/peij_3_3/N35 )
         );
  AND4_X4 \pool/pool/pe_b/peij_3_3/U16  ( .A1(1'b1), .A2(
        \pool/pool/pe_b_i_data[3][3] ), .A3(\pool/pool/pe_b/int_pe_en[3][3] ), 
        .A4(\pool/pool/pe_b/peij_3_3/n18 ), .ZN(\pool/pool/pe_b/peij_3_3/N36 )
         );
  DFFR_X1 \pool/pool/pe_b/peij_3_3/q_im_reg[0]  ( .D(
        \pool/pool/pe_b/peij_3_3/N33 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_3/n12 ), .Q(\pool/pool/pe_b/peij_3_3/sgnext [0]) );
  DFFR_X1 \pool/pool/pe_b/peij_3_3/q_im_reg[1]  ( .D(
        \pool/pool/pe_b/peij_3_3/N34 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_3/n12 ), .Q(\pool/pool/pe_b/peij_3_3/sgnext [1]) );
  DFFR_X1 \pool/pool/pe_b/peij_3_3/q_im_reg[2]  ( .D(
        \pool/pool/pe_b/peij_3_3/N35 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_3/n12 ), .Q(\pool/pool/pe_b/peij_3_3/sgnext [2]) );
  DFFR_X1 \pool/pool/pe_b/peij_3_3/q_im_reg[3]  ( .D(
        \pool/pool/pe_b/peij_3_3/N36 ), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_3/n12 ), .Q(\pool/pool/pe_b/peij_3_3/sgnext_10 ) );
  SDFFR_X1 \pool/pool/pe_b/peij_3_3/q_k_reg  ( .D(1'b0), .SI(
        \pool/pool/pe_b/peij_3_3/n18 ), .SE(1'b0), .CK(clk), .RN(
        \pool/pool/pe_b/peij_3_3/n12 ), .Q(\pool/pool/pe_b/peij_3_3/q_k ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/U11  ( .A(
        \pool/pool/pe_b/peij_3_3/sgnext [0]), .B(\pool/pool/pe_b/peij_3_3/q_k ), .Z(\pool/pool/pe_b/peij_3_3/add/notb [0]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/U10  ( .A(
        \pool/pool/pe_b/peij_3_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_3/q_k ), .Z(\pool/pool/pe_b/peij_3_3/add/notb [10]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/U9  ( .A(
        \pool/pool/pe_b/peij_3_3/sgnext [1]), .B(\pool/pool/pe_b/peij_3_3/q_k ), .Z(\pool/pool/pe_b/peij_3_3/add/notb [1]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/U8  ( .A(
        \pool/pool/pe_b/peij_3_3/sgnext [2]), .B(\pool/pool/pe_b/peij_3_3/q_k ), .Z(\pool/pool/pe_b/peij_3_3/add/notb [2]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/U7  ( .A(
        \pool/pool/pe_b/peij_3_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_3/q_k ), .Z(\pool/pool/pe_b/peij_3_3/add/notb [3]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/U6  ( .A(
        \pool/pool/pe_b/peij_3_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_3/q_k ), .Z(\pool/pool/pe_b/peij_3_3/add/notb [4]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/U5  ( .A(
        \pool/pool/pe_b/peij_3_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_3/q_k ), .Z(\pool/pool/pe_b/peij_3_3/add/notb [5]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/U4  ( .A(
        \pool/pool/pe_b/peij_3_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_3/q_k ), .Z(\pool/pool/pe_b/peij_3_3/add/notb [6]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/U3  ( .A(
        \pool/pool/pe_b/peij_3_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_3/q_k ), .Z(\pool/pool/pe_b/peij_3_3/add/notb [7]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/U2  ( .A(
        \pool/pool/pe_b/peij_3_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_3/q_k ), .Z(\pool/pool/pe_b/peij_3_3/add/notb [8]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/U1  ( .A(
        \pool/pool/pe_b/peij_3_3/sgnext_10 ), .B(\pool/pool/pe_b/peij_3_3/q_k ), .Z(\pool/pool/pe_b/peij_3_3/add/notb [9]) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_0/U4  ( .A(
        \pool/pool/pe_b_o_data[3][0] ), .B(
        \pool/pool/pe_b/peij_3_3/add/notb [0]), .Z(
        \pool/pool/pe_b/peij_3_3/add/fai_0/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_0/U3  ( .A(
        \pool/pool/pe_b/peij_3_3/q_k ), .B(
        \pool/pool/pe_b/peij_3_3/add/fai_0/n3 ), .Z(
        \pool/pool/pe_b/peij_3_3/d_acc [0]) );
  INV_X2 \pool/pool/pe_b/peij_3_3/add/fai_0/U2  ( .A(
        \pool/pool/pe_b/peij_3_3/add/fai_0/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_3/add/cprop [1]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_3/add/fai_0/U1  ( .A1(
        \pool/pool/pe_b/peij_3_3/add/notb [0]), .A2(
        \pool/pool/pe_b_o_data[3][0] ), .B1(
        \pool/pool/pe_b/peij_3_3/add/fai_0/n3 ), .B2(
        \pool/pool/pe_b/peij_3_3/q_k ), .ZN(
        \pool/pool/pe_b/peij_3_3/add/fai_0/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_1/U4  ( .A(
        \pool/pool/pe_b_o_data[3][1] ), .B(
        \pool/pool/pe_b/peij_3_3/add/notb [1]), .Z(
        \pool/pool/pe_b/peij_3_3/add/fai_1/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_1/U3  ( .A(
        \pool/pool/pe_b/peij_3_3/add/cprop [1]), .B(
        \pool/pool/pe_b/peij_3_3/add/fai_1/n3 ), .Z(
        \pool/pool/pe_b/peij_3_3/d_acc [1]) );
  INV_X2 \pool/pool/pe_b/peij_3_3/add/fai_1/U2  ( .A(
        \pool/pool/pe_b/peij_3_3/add/fai_1/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_3/add/cprop [2]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_3/add/fai_1/U1  ( .A1(
        \pool/pool/pe_b/peij_3_3/add/notb [1]), .A2(
        \pool/pool/pe_b_o_data[3][1] ), .B1(
        \pool/pool/pe_b/peij_3_3/add/fai_1/n3 ), .B2(
        \pool/pool/pe_b/peij_3_3/add/cprop [1]), .ZN(
        \pool/pool/pe_b/peij_3_3/add/fai_1/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_2/U4  ( .A(
        \pool/pool/pe_b_o_data[3][2] ), .B(
        \pool/pool/pe_b/peij_3_3/add/notb [2]), .Z(
        \pool/pool/pe_b/peij_3_3/add/fai_2/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_2/U3  ( .A(
        \pool/pool/pe_b/peij_3_3/add/cprop [2]), .B(
        \pool/pool/pe_b/peij_3_3/add/fai_2/n3 ), .Z(
        \pool/pool/pe_b/peij_3_3/d_acc [2]) );
  INV_X2 \pool/pool/pe_b/peij_3_3/add/fai_2/U2  ( .A(
        \pool/pool/pe_b/peij_3_3/add/fai_2/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_3/add/cprop [3]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_3/add/fai_2/U1  ( .A1(
        \pool/pool/pe_b/peij_3_3/add/notb [2]), .A2(
        \pool/pool/pe_b_o_data[3][2] ), .B1(
        \pool/pool/pe_b/peij_3_3/add/fai_2/n3 ), .B2(
        \pool/pool/pe_b/peij_3_3/add/cprop [2]), .ZN(
        \pool/pool/pe_b/peij_3_3/add/fai_2/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_3/U4  ( .A(
        \pool/pool/pe_b_o_data[3][3] ), .B(
        \pool/pool/pe_b/peij_3_3/add/notb [3]), .Z(
        \pool/pool/pe_b/peij_3_3/add/fai_3/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_3/U3  ( .A(
        \pool/pool/pe_b/peij_3_3/add/cprop [3]), .B(
        \pool/pool/pe_b/peij_3_3/add/fai_3/n3 ), .Z(
        \pool/pool/pe_b/peij_3_3/d_acc [3]) );
  INV_X2 \pool/pool/pe_b/peij_3_3/add/fai_3/U2  ( .A(
        \pool/pool/pe_b/peij_3_3/add/fai_3/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_3/add/cprop [4]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_3/add/fai_3/U1  ( .A1(
        \pool/pool/pe_b/peij_3_3/add/notb [3]), .A2(
        \pool/pool/pe_b_o_data[3][3] ), .B1(
        \pool/pool/pe_b/peij_3_3/add/fai_3/n3 ), .B2(
        \pool/pool/pe_b/peij_3_3/add/cprop [3]), .ZN(
        \pool/pool/pe_b/peij_3_3/add/fai_3/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_4/U4  ( .A(
        \pool/pool/pe_b_o_data[3][4] ), .B(
        \pool/pool/pe_b/peij_3_3/add/notb [4]), .Z(
        \pool/pool/pe_b/peij_3_3/add/fai_4/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_4/U3  ( .A(
        \pool/pool/pe_b/peij_3_3/add/cprop [4]), .B(
        \pool/pool/pe_b/peij_3_3/add/fai_4/n3 ), .Z(
        \pool/pool/pe_b/peij_3_3/d_acc [4]) );
  INV_X2 \pool/pool/pe_b/peij_3_3/add/fai_4/U2  ( .A(
        \pool/pool/pe_b/peij_3_3/add/fai_4/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_3/add/cprop [5]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_3/add/fai_4/U1  ( .A1(
        \pool/pool/pe_b/peij_3_3/add/notb [4]), .A2(
        \pool/pool/pe_b_o_data[3][4] ), .B1(
        \pool/pool/pe_b/peij_3_3/add/fai_4/n3 ), .B2(
        \pool/pool/pe_b/peij_3_3/add/cprop [4]), .ZN(
        \pool/pool/pe_b/peij_3_3/add/fai_4/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_5/U4  ( .A(
        \pool/pool/pe_b_o_data[3][5] ), .B(
        \pool/pool/pe_b/peij_3_3/add/notb [5]), .Z(
        \pool/pool/pe_b/peij_3_3/add/fai_5/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_5/U3  ( .A(
        \pool/pool/pe_b/peij_3_3/add/cprop [5]), .B(
        \pool/pool/pe_b/peij_3_3/add/fai_5/n3 ), .Z(
        \pool/pool/pe_b/peij_3_3/d_acc [5]) );
  INV_X2 \pool/pool/pe_b/peij_3_3/add/fai_5/U2  ( .A(
        \pool/pool/pe_b/peij_3_3/add/fai_5/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_3/add/cprop [6]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_3/add/fai_5/U1  ( .A1(
        \pool/pool/pe_b/peij_3_3/add/notb [5]), .A2(
        \pool/pool/pe_b_o_data[3][5] ), .B1(
        \pool/pool/pe_b/peij_3_3/add/fai_5/n3 ), .B2(
        \pool/pool/pe_b/peij_3_3/add/cprop [5]), .ZN(
        \pool/pool/pe_b/peij_3_3/add/fai_5/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_6/U4  ( .A(
        \pool/pool/pe_b_o_data[3][6] ), .B(
        \pool/pool/pe_b/peij_3_3/add/notb [6]), .Z(
        \pool/pool/pe_b/peij_3_3/add/fai_6/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_6/U3  ( .A(
        \pool/pool/pe_b/peij_3_3/add/cprop [6]), .B(
        \pool/pool/pe_b/peij_3_3/add/fai_6/n3 ), .Z(
        \pool/pool/pe_b/peij_3_3/d_acc [6]) );
  INV_X2 \pool/pool/pe_b/peij_3_3/add/fai_6/U2  ( .A(
        \pool/pool/pe_b/peij_3_3/add/fai_6/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_3/add/cprop [7]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_3/add/fai_6/U1  ( .A1(
        \pool/pool/pe_b/peij_3_3/add/notb [6]), .A2(
        \pool/pool/pe_b_o_data[3][6] ), .B1(
        \pool/pool/pe_b/peij_3_3/add/fai_6/n3 ), .B2(
        \pool/pool/pe_b/peij_3_3/add/cprop [6]), .ZN(
        \pool/pool/pe_b/peij_3_3/add/fai_6/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_7/U4  ( .A(
        \pool/pool/pe_b_o_data[3][7] ), .B(
        \pool/pool/pe_b/peij_3_3/add/notb [7]), .Z(
        \pool/pool/pe_b/peij_3_3/add/fai_7/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_7/U3  ( .A(
        \pool/pool/pe_b/peij_3_3/add/cprop [7]), .B(
        \pool/pool/pe_b/peij_3_3/add/fai_7/n3 ), .Z(
        \pool/pool/pe_b/peij_3_3/d_acc [7]) );
  INV_X2 \pool/pool/pe_b/peij_3_3/add/fai_7/U2  ( .A(
        \pool/pool/pe_b/peij_3_3/add/fai_7/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_3/add/cprop [8]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_3/add/fai_7/U1  ( .A1(
        \pool/pool/pe_b/peij_3_3/add/notb [7]), .A2(
        \pool/pool/pe_b_o_data[3][7] ), .B1(
        \pool/pool/pe_b/peij_3_3/add/fai_7/n3 ), .B2(
        \pool/pool/pe_b/peij_3_3/add/cprop [7]), .ZN(
        \pool/pool/pe_b/peij_3_3/add/fai_7/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_8/U4  ( .A(
        \pool/pool/pe_b_o_data[3][8] ), .B(
        \pool/pool/pe_b/peij_3_3/add/notb [8]), .Z(
        \pool/pool/pe_b/peij_3_3/add/fai_8/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_8/U3  ( .A(
        \pool/pool/pe_b/peij_3_3/add/cprop [8]), .B(
        \pool/pool/pe_b/peij_3_3/add/fai_8/n3 ), .Z(
        \pool/pool/pe_b/peij_3_3/d_acc [8]) );
  INV_X2 \pool/pool/pe_b/peij_3_3/add/fai_8/U2  ( .A(
        \pool/pool/pe_b/peij_3_3/add/fai_8/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_3/add/cprop [9]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_3/add/fai_8/U1  ( .A1(
        \pool/pool/pe_b/peij_3_3/add/notb [8]), .A2(
        \pool/pool/pe_b_o_data[3][8] ), .B1(
        \pool/pool/pe_b/peij_3_3/add/fai_8/n3 ), .B2(
        \pool/pool/pe_b/peij_3_3/add/cprop [8]), .ZN(
        \pool/pool/pe_b/peij_3_3/add/fai_8/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_9/U4  ( .A(
        \pool/pool/pe_b_o_data[3][9] ), .B(
        \pool/pool/pe_b/peij_3_3/add/notb [9]), .Z(
        \pool/pool/pe_b/peij_3_3/add/fai_9/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_9/U3  ( .A(
        \pool/pool/pe_b/peij_3_3/add/cprop [9]), .B(
        \pool/pool/pe_b/peij_3_3/add/fai_9/n3 ), .Z(
        \pool/pool/pe_b/peij_3_3/d_acc [9]) );
  INV_X2 \pool/pool/pe_b/peij_3_3/add/fai_9/U2  ( .A(
        \pool/pool/pe_b/peij_3_3/add/fai_9/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_3/add/cprop [10]) );
  AOI22_X2 \pool/pool/pe_b/peij_3_3/add/fai_9/U1  ( .A1(
        \pool/pool/pe_b/peij_3_3/add/notb [9]), .A2(
        \pool/pool/pe_b_o_data[3][9] ), .B1(
        \pool/pool/pe_b/peij_3_3/add/fai_9/n3 ), .B2(
        \pool/pool/pe_b/peij_3_3/add/cprop [9]), .ZN(
        \pool/pool/pe_b/peij_3_3/add/fai_9/n1 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_10/U4  ( .A(
        \pool/pool/pe_b_o_data[3][10] ), .B(
        \pool/pool/pe_b/peij_3_3/add/notb [10]), .Z(
        \pool/pool/pe_b/peij_3_3/add/fai_10/n3 ) );
  XOR2_X1 \pool/pool/pe_b/peij_3_3/add/fai_10/U3  ( .A(
        \pool/pool/pe_b/peij_3_3/add/cprop [10]), .B(
        \pool/pool/pe_b/peij_3_3/add/fai_10/n3 ), .Z(
        \pool/pool/pe_b/peij_3_3/d_acc [10]) );
  INV_X2 \pool/pool/pe_b/peij_3_3/add/fai_10/U2  ( .A(
        \pool/pool/pe_b/peij_3_3/add/fai_10/n1 ), .ZN(
        \pool/pool/pe_b/peij_3_3/add/c_out ) );
  AOI22_X2 \pool/pool/pe_b/peij_3_3/add/fai_10/U1  ( .A1(
        \pool/pool/pe_b/peij_3_3/add/notb [10]), .A2(
        \pool/pool/pe_b_o_data[3][10] ), .B1(
        \pool/pool/pe_b/peij_3_3/add/fai_10/n3 ), .B2(
        \pool/pool/pe_b/peij_3_3/add/cprop [10]), .ZN(
        \pool/pool/pe_b/peij_3_3/add/fai_10/n1 ) );
  DFFR_X1 \pool/pool/count/cnt_out_reg[1]  ( .D(\pool/pool/count/n15 ), .CK(
        clk), .RN(\pool/pool/count/n16 ), .Q(\pool/pool/cnt[1] ), .QN(
        \pool/pool/count/n4 ) );
  DFFR_X1 \pool/pool/count/cnt_out_reg[0]  ( .D(\pool/pool/count/n17 ), .CK(
        clk), .RN(\pool/pool/count/n16 ), .Q(\pool/pool/cnt[0] ), .QN(
        \pool/pool/count/n7 ) );
  DFFR_X1 \pool/pool/count/terminal_cnt_reg  ( .D(\pool/pool/count/n18 ), .CK(
        clk), .RN(\pool/pool/count/n16 ), .Q(\pool/tc ), .QN(
        \pool/pool/count/n10 ) );
  INV_X1 \pool/pool/count/U18  ( .A(1'b1), .ZN(\pool/pool/count/n12 ) );
  XOR2_X1 \pool/pool/count/U17  ( .A(\pool/pool/cnt[1] ), .B(1'b1), .Z(
        \pool/pool/count/n13 ) );
  INV_X1 \pool/pool/count/U15  ( .A(\pool/pool/count/n13 ), .ZN(
        \pool/pool/count/n14 ) );
  OAI33_X1 \pool/pool/count/U14  ( .A1(\pool/pool/count/n12 ), .A2(
        \pool/pool/cnt[0] ), .A3(\pool/pool/count/n13 ), .B1(
        \pool/pool/count/n7 ), .B2(1'b1), .B3(\pool/pool/count/n14 ), .ZN(
        \pool/pool/count/n11 ) );
  INV_X1 \pool/pool/count/U13  ( .A(\pool/pool/count/n11 ), .ZN(
        \pool/pool/count/n9 ) );
  NAND2_X1 \pool/pool/count/U11  ( .A1(\pool/en_cnt ), .A2(
        \pool/pool/count/n10 ), .ZN(\pool/pool/count/n6 ) );
  OAI22_X1 \pool/pool/count/U10  ( .A1(\pool/pool/count/n9 ), .A2(
        \pool/pool/count/n6 ), .B1(\pool/en_cnt ), .B2(\pool/pool/count/n10 ), 
        .ZN(\pool/pool/count/n18 ) );
  OAI22_X1 \pool/pool/count/U9  ( .A1(\pool/en_cnt ), .A2(\pool/pool/count/n7 ), .B1(\pool/pool/cnt[0] ), .B2(\pool/pool/count/n6 ), .ZN(
        \pool/pool/count/n17 ) );
  INV_X1 \pool/pool/count/U8  ( .A(\pool/rst_cnt ), .ZN(\pool/pool/count/n16 )
         );
  OAI21_X1 \pool/pool/count/U7  ( .B1(\pool/pool/cnt[0] ), .B2(\pool/tc ), .A(
        \pool/en_cnt ), .ZN(\pool/pool/count/n8 ) );
  INV_X1 \pool/pool/count/U6  ( .A(\pool/pool/count/n8 ), .ZN(
        \pool/pool/count/n3 ) );
  OR3_X1 \pool/pool/count/U4  ( .A1(\pool/pool/count/n6 ), .A2(
        \pool/pool/cnt[1] ), .A3(\pool/pool/count/n7 ), .ZN(
        \pool/pool/count/n5 ) );
  OAI21_X1 \pool/pool/count/U3  ( .B1(\pool/pool/count/n3 ), .B2(
        \pool/pool/count/n4 ), .A(\pool/pool/count/n5 ), .ZN(
        \pool/pool/count/n15 ) );
  XOR2_X1 \pool/pool/shift_row0/U25  ( .A(\pool/pool/pe_b_o_data[0][35] ), .B(
        \pool/pool/pe_b_o_data[0][34] ), .Z(o_pool_1[12]) );
  XOR2_X1 \pool/pool/shift_row0/U24  ( .A(\pool/pool/shift_row0/n1 ), .B(
        \pool/pool/shift_row0/n12 ), .Z(o_pool_1[13]) );
  XOR2_X1 \pool/pool/shift_row0/U23  ( .A(\pool/pool/pe_b_o_data[0][37] ), .B(
        \pool/pool/shift_row0/n11 ), .Z(o_pool_1[14]) );
  XOR2_X1 \pool/pool/shift_row0/U22  ( .A(\pool/pool/pe_b_o_data[0][24] ), .B(
        \pool/pool/pe_b_o_data[0][23] ), .Z(o_pool_1[8]) );
  XOR2_X1 \pool/pool/shift_row0/U21  ( .A(\pool/pool/shift_row0/n2 ), .B(
        \pool/pool/shift_row0/n10 ), .Z(o_pool_1[9]) );
  XOR2_X1 \pool/pool/shift_row0/U20  ( .A(\pool/pool/pe_b_o_data[0][26] ), .B(
        \pool/pool/shift_row0/n9 ), .Z(o_pool_1[10]) );
  XOR2_X1 \pool/pool/shift_row0/U19  ( .A(\pool/pool/pe_b_o_data[0][13] ), .B(
        \pool/pool/pe_b_o_data[0][12] ), .Z(o_pool_1[4]) );
  XOR2_X1 \pool/pool/shift_row0/U18  ( .A(\pool/pool/shift_row0/n3 ), .B(
        \pool/pool/shift_row0/n8 ), .Z(o_pool_1[5]) );
  XOR2_X1 \pool/pool/shift_row0/U17  ( .A(\pool/pool/pe_b_o_data[0][15] ), .B(
        \pool/pool/shift_row0/n7 ), .Z(o_pool_1[6]) );
  XOR2_X1 \pool/pool/shift_row0/U16  ( .A(\pool/pool/pe_b_o_data[0][2] ), .B(
        \pool/pool/pe_b_o_data[0][1] ), .Z(o_pool_1[0]) );
  XOR2_X1 \pool/pool/shift_row0/U15  ( .A(\pool/pool/shift_row0/n4 ), .B(
        \pool/pool/shift_row0/n6 ), .Z(o_pool_1[1]) );
  XOR2_X1 \pool/pool/shift_row0/U14  ( .A(\pool/pool/pe_b_o_data[0][4] ), .B(
        \pool/pool/shift_row0/n5 ), .Z(o_pool_1[2]) );
  INV_X2 \pool/pool/shift_row0/U13  ( .A(\pool/pool/pe_b_o_data[0][3] ), .ZN(
        \pool/pool/shift_row0/n4 ) );
  INV_X2 \pool/pool/shift_row0/U12  ( .A(\pool/pool/pe_b_o_data[0][14] ), .ZN(
        \pool/pool/shift_row0/n3 ) );
  INV_X2 \pool/pool/shift_row0/U11  ( .A(\pool/pool/pe_b_o_data[0][25] ), .ZN(
        \pool/pool/shift_row0/n2 ) );
  INV_X2 \pool/pool/shift_row0/U10  ( .A(\pool/pool/pe_b_o_data[0][36] ), .ZN(
        \pool/pool/shift_row0/n1 ) );
  NAND2_X2 \pool/pool/shift_row0/U9  ( .A1(\pool/pool/pe_b_o_data[0][35] ), 
        .A2(\pool/pool/pe_b_o_data[0][34] ), .ZN(\pool/pool/shift_row0/n12 )
         );
  NOR2_X2 \pool/pool/shift_row0/U8  ( .A1(\pool/pool/shift_row0/n12 ), .A2(
        \pool/pool/shift_row0/n1 ), .ZN(\pool/pool/shift_row0/n11 ) );
  NAND2_X2 \pool/pool/shift_row0/U7  ( .A1(\pool/pool/pe_b_o_data[0][24] ), 
        .A2(\pool/pool/pe_b_o_data[0][23] ), .ZN(\pool/pool/shift_row0/n10 )
         );
  NOR2_X2 \pool/pool/shift_row0/U6  ( .A1(\pool/pool/shift_row0/n10 ), .A2(
        \pool/pool/shift_row0/n2 ), .ZN(\pool/pool/shift_row0/n9 ) );
  NAND2_X2 \pool/pool/shift_row0/U5  ( .A1(\pool/pool/pe_b_o_data[0][13] ), 
        .A2(\pool/pool/pe_b_o_data[0][12] ), .ZN(\pool/pool/shift_row0/n8 ) );
  NOR2_X2 \pool/pool/shift_row0/U4  ( .A1(\pool/pool/shift_row0/n8 ), .A2(
        \pool/pool/shift_row0/n3 ), .ZN(\pool/pool/shift_row0/n7 ) );
  NAND2_X2 \pool/pool/shift_row0/U3  ( .A1(\pool/pool/pe_b_o_data[0][2] ), 
        .A2(\pool/pool/pe_b_o_data[0][1] ), .ZN(\pool/pool/shift_row0/n6 ) );
  NOR2_X2 \pool/pool/shift_row0/U2  ( .A1(\pool/pool/shift_row0/n6 ), .A2(
        \pool/pool/shift_row0/n4 ), .ZN(\pool/pool/shift_row0/n5 ) );
  XOR2_X1 \pool/pool/shift_row1/U25  ( .A(\pool/pool/pe_b_o_data[1][35] ), .B(
        \pool/pool/pe_b_o_data[1][34] ), .Z(o_pool_2[12]) );
  XOR2_X1 \pool/pool/shift_row1/U24  ( .A(\pool/pool/shift_row1/n24 ), .B(
        \pool/pool/shift_row1/n13 ), .Z(o_pool_2[13]) );
  XOR2_X1 \pool/pool/shift_row1/U23  ( .A(\pool/pool/pe_b_o_data[1][37] ), .B(
        \pool/pool/shift_row1/n14 ), .Z(o_pool_2[14]) );
  XOR2_X1 \pool/pool/shift_row1/U22  ( .A(\pool/pool/pe_b_o_data[1][24] ), .B(
        \pool/pool/pe_b_o_data[1][23] ), .Z(o_pool_2[8]) );
  XOR2_X1 \pool/pool/shift_row1/U21  ( .A(\pool/pool/shift_row1/n23 ), .B(
        \pool/pool/shift_row1/n15 ), .Z(o_pool_2[9]) );
  XOR2_X1 \pool/pool/shift_row1/U20  ( .A(\pool/pool/pe_b_o_data[1][26] ), .B(
        \pool/pool/shift_row1/n16 ), .Z(o_pool_2[10]) );
  XOR2_X1 \pool/pool/shift_row1/U19  ( .A(\pool/pool/pe_b_o_data[1][13] ), .B(
        \pool/pool/pe_b_o_data[1][12] ), .Z(o_pool_2[4]) );
  XOR2_X1 \pool/pool/shift_row1/U18  ( .A(\pool/pool/shift_row1/n22 ), .B(
        \pool/pool/shift_row1/n17 ), .Z(o_pool_2[5]) );
  XOR2_X1 \pool/pool/shift_row1/U17  ( .A(\pool/pool/pe_b_o_data[1][15] ), .B(
        \pool/pool/shift_row1/n18 ), .Z(o_pool_2[6]) );
  XOR2_X1 \pool/pool/shift_row1/U16  ( .A(\pool/pool/pe_b_o_data[1][2] ), .B(
        \pool/pool/pe_b_o_data[1][1] ), .Z(o_pool_2[0]) );
  XOR2_X1 \pool/pool/shift_row1/U15  ( .A(\pool/pool/shift_row1/n21 ), .B(
        \pool/pool/shift_row1/n19 ), .Z(o_pool_2[1]) );
  XOR2_X1 \pool/pool/shift_row1/U14  ( .A(\pool/pool/pe_b_o_data[1][4] ), .B(
        \pool/pool/shift_row1/n20 ), .Z(o_pool_2[2]) );
  INV_X2 \pool/pool/shift_row1/U13  ( .A(\pool/pool/pe_b_o_data[1][3] ), .ZN(
        \pool/pool/shift_row1/n21 ) );
  INV_X2 \pool/pool/shift_row1/U12  ( .A(\pool/pool/pe_b_o_data[1][14] ), .ZN(
        \pool/pool/shift_row1/n22 ) );
  INV_X2 \pool/pool/shift_row1/U11  ( .A(\pool/pool/pe_b_o_data[1][25] ), .ZN(
        \pool/pool/shift_row1/n23 ) );
  INV_X2 \pool/pool/shift_row1/U10  ( .A(\pool/pool/pe_b_o_data[1][36] ), .ZN(
        \pool/pool/shift_row1/n24 ) );
  NAND2_X2 \pool/pool/shift_row1/U9  ( .A1(\pool/pool/pe_b_o_data[1][35] ), 
        .A2(\pool/pool/pe_b_o_data[1][34] ), .ZN(\pool/pool/shift_row1/n13 )
         );
  NOR2_X2 \pool/pool/shift_row1/U8  ( .A1(\pool/pool/shift_row1/n13 ), .A2(
        \pool/pool/shift_row1/n24 ), .ZN(\pool/pool/shift_row1/n14 ) );
  NAND2_X2 \pool/pool/shift_row1/U7  ( .A1(\pool/pool/pe_b_o_data[1][24] ), 
        .A2(\pool/pool/pe_b_o_data[1][23] ), .ZN(\pool/pool/shift_row1/n15 )
         );
  NOR2_X2 \pool/pool/shift_row1/U6  ( .A1(\pool/pool/shift_row1/n15 ), .A2(
        \pool/pool/shift_row1/n23 ), .ZN(\pool/pool/shift_row1/n16 ) );
  NAND2_X2 \pool/pool/shift_row1/U5  ( .A1(\pool/pool/pe_b_o_data[1][13] ), 
        .A2(\pool/pool/pe_b_o_data[1][12] ), .ZN(\pool/pool/shift_row1/n17 )
         );
  NOR2_X2 \pool/pool/shift_row1/U4  ( .A1(\pool/pool/shift_row1/n17 ), .A2(
        \pool/pool/shift_row1/n22 ), .ZN(\pool/pool/shift_row1/n18 ) );
  NAND2_X2 \pool/pool/shift_row1/U3  ( .A1(\pool/pool/pe_b_o_data[1][2] ), 
        .A2(\pool/pool/pe_b_o_data[1][1] ), .ZN(\pool/pool/shift_row1/n19 ) );
  NOR2_X2 \pool/pool/shift_row1/U2  ( .A1(\pool/pool/shift_row1/n19 ), .A2(
        \pool/pool/shift_row1/n21 ), .ZN(\pool/pool/shift_row1/n20 ) );
  XOR2_X1 \pool/pool/shift_row2/U25  ( .A(\pool/pool/pe_b_o_data[2][35] ), .B(
        \pool/pool/pe_b_o_data[2][34] ), .Z(o_pool_3[12]) );
  XOR2_X1 \pool/pool/shift_row2/U24  ( .A(\pool/pool/shift_row2/n24 ), .B(
        \pool/pool/shift_row2/n13 ), .Z(o_pool_3[13]) );
  XOR2_X1 \pool/pool/shift_row2/U23  ( .A(\pool/pool/pe_b_o_data[2][37] ), .B(
        \pool/pool/shift_row2/n14 ), .Z(o_pool_3[14]) );
  XOR2_X1 \pool/pool/shift_row2/U22  ( .A(\pool/pool/pe_b_o_data[2][24] ), .B(
        \pool/pool/pe_b_o_data[2][23] ), .Z(o_pool_3[8]) );
  XOR2_X1 \pool/pool/shift_row2/U21  ( .A(\pool/pool/shift_row2/n23 ), .B(
        \pool/pool/shift_row2/n15 ), .Z(o_pool_3[9]) );
  XOR2_X1 \pool/pool/shift_row2/U20  ( .A(\pool/pool/pe_b_o_data[2][26] ), .B(
        \pool/pool/shift_row2/n16 ), .Z(o_pool_3[10]) );
  XOR2_X1 \pool/pool/shift_row2/U19  ( .A(\pool/pool/pe_b_o_data[2][13] ), .B(
        \pool/pool/pe_b_o_data[2][12] ), .Z(o_pool_3[4]) );
  XOR2_X1 \pool/pool/shift_row2/U18  ( .A(\pool/pool/shift_row2/n22 ), .B(
        \pool/pool/shift_row2/n17 ), .Z(o_pool_3[5]) );
  XOR2_X1 \pool/pool/shift_row2/U17  ( .A(\pool/pool/pe_b_o_data[2][15] ), .B(
        \pool/pool/shift_row2/n18 ), .Z(o_pool_3[6]) );
  XOR2_X1 \pool/pool/shift_row2/U16  ( .A(\pool/pool/pe_b_o_data[2][2] ), .B(
        \pool/pool/pe_b_o_data[2][1] ), .Z(o_pool_3[0]) );
  XOR2_X1 \pool/pool/shift_row2/U15  ( .A(\pool/pool/shift_row2/n21 ), .B(
        \pool/pool/shift_row2/n19 ), .Z(o_pool_3[1]) );
  XOR2_X1 \pool/pool/shift_row2/U14  ( .A(\pool/pool/pe_b_o_data[2][4] ), .B(
        \pool/pool/shift_row2/n20 ), .Z(o_pool_3[2]) );
  INV_X2 \pool/pool/shift_row2/U13  ( .A(\pool/pool/pe_b_o_data[2][3] ), .ZN(
        \pool/pool/shift_row2/n21 ) );
  INV_X2 \pool/pool/shift_row2/U12  ( .A(\pool/pool/pe_b_o_data[2][14] ), .ZN(
        \pool/pool/shift_row2/n22 ) );
  INV_X2 \pool/pool/shift_row2/U11  ( .A(\pool/pool/pe_b_o_data[2][25] ), .ZN(
        \pool/pool/shift_row2/n23 ) );
  INV_X2 \pool/pool/shift_row2/U10  ( .A(\pool/pool/pe_b_o_data[2][36] ), .ZN(
        \pool/pool/shift_row2/n24 ) );
  NAND2_X2 \pool/pool/shift_row2/U9  ( .A1(\pool/pool/pe_b_o_data[2][35] ), 
        .A2(\pool/pool/pe_b_o_data[2][34] ), .ZN(\pool/pool/shift_row2/n13 )
         );
  NOR2_X2 \pool/pool/shift_row2/U8  ( .A1(\pool/pool/shift_row2/n13 ), .A2(
        \pool/pool/shift_row2/n24 ), .ZN(\pool/pool/shift_row2/n14 ) );
  NAND2_X2 \pool/pool/shift_row2/U7  ( .A1(\pool/pool/pe_b_o_data[2][24] ), 
        .A2(\pool/pool/pe_b_o_data[2][23] ), .ZN(\pool/pool/shift_row2/n15 )
         );
  NOR2_X2 \pool/pool/shift_row2/U6  ( .A1(\pool/pool/shift_row2/n15 ), .A2(
        \pool/pool/shift_row2/n23 ), .ZN(\pool/pool/shift_row2/n16 ) );
  NAND2_X2 \pool/pool/shift_row2/U5  ( .A1(\pool/pool/pe_b_o_data[2][13] ), 
        .A2(\pool/pool/pe_b_o_data[2][12] ), .ZN(\pool/pool/shift_row2/n17 )
         );
  NOR2_X2 \pool/pool/shift_row2/U4  ( .A1(\pool/pool/shift_row2/n17 ), .A2(
        \pool/pool/shift_row2/n22 ), .ZN(\pool/pool/shift_row2/n18 ) );
  NAND2_X2 \pool/pool/shift_row2/U3  ( .A1(\pool/pool/pe_b_o_data[2][2] ), 
        .A2(\pool/pool/pe_b_o_data[2][1] ), .ZN(\pool/pool/shift_row2/n19 ) );
  NOR2_X2 \pool/pool/shift_row2/U2  ( .A1(\pool/pool/shift_row2/n19 ), .A2(
        \pool/pool/shift_row2/n21 ), .ZN(\pool/pool/shift_row2/n20 ) );
  XOR2_X1 \pool/pool/shift_row3/U25  ( .A(\pool/pool/pe_b_o_data[3][35] ), .B(
        \pool/pool/pe_b_o_data[3][34] ), .Z(o_pool_4[12]) );
  XOR2_X1 \pool/pool/shift_row3/U24  ( .A(\pool/pool/shift_row3/n24 ), .B(
        \pool/pool/shift_row3/n13 ), .Z(o_pool_4[13]) );
  XOR2_X1 \pool/pool/shift_row3/U23  ( .A(\pool/pool/pe_b_o_data[3][37] ), .B(
        \pool/pool/shift_row3/n14 ), .Z(o_pool_4[14]) );
  XOR2_X1 \pool/pool/shift_row3/U22  ( .A(\pool/pool/pe_b_o_data[3][24] ), .B(
        \pool/pool/pe_b_o_data[3][23] ), .Z(o_pool_4[8]) );
  XOR2_X1 \pool/pool/shift_row3/U21  ( .A(\pool/pool/shift_row3/n23 ), .B(
        \pool/pool/shift_row3/n15 ), .Z(o_pool_4[9]) );
  XOR2_X1 \pool/pool/shift_row3/U20  ( .A(\pool/pool/pe_b_o_data[3][26] ), .B(
        \pool/pool/shift_row3/n16 ), .Z(o_pool_4[10]) );
  XOR2_X1 \pool/pool/shift_row3/U19  ( .A(\pool/pool/pe_b_o_data[3][13] ), .B(
        \pool/pool/pe_b_o_data[3][12] ), .Z(o_pool_4[4]) );
  XOR2_X1 \pool/pool/shift_row3/U18  ( .A(\pool/pool/shift_row3/n22 ), .B(
        \pool/pool/shift_row3/n17 ), .Z(o_pool_4[5]) );
  XOR2_X1 \pool/pool/shift_row3/U17  ( .A(\pool/pool/pe_b_o_data[3][15] ), .B(
        \pool/pool/shift_row3/n18 ), .Z(o_pool_4[6]) );
  XOR2_X1 \pool/pool/shift_row3/U16  ( .A(\pool/pool/pe_b_o_data[3][2] ), .B(
        \pool/pool/pe_b_o_data[3][1] ), .Z(o_pool_4[0]) );
  XOR2_X1 \pool/pool/shift_row3/U15  ( .A(\pool/pool/shift_row3/n21 ), .B(
        \pool/pool/shift_row3/n19 ), .Z(o_pool_4[1]) );
  XOR2_X1 \pool/pool/shift_row3/U14  ( .A(\pool/pool/pe_b_o_data[3][4] ), .B(
        \pool/pool/shift_row3/n20 ), .Z(o_pool_4[2]) );
  INV_X2 \pool/pool/shift_row3/U13  ( .A(\pool/pool/pe_b_o_data[3][3] ), .ZN(
        \pool/pool/shift_row3/n21 ) );
  INV_X2 \pool/pool/shift_row3/U12  ( .A(\pool/pool/pe_b_o_data[3][14] ), .ZN(
        \pool/pool/shift_row3/n22 ) );
  INV_X2 \pool/pool/shift_row3/U11  ( .A(\pool/pool/pe_b_o_data[3][25] ), .ZN(
        \pool/pool/shift_row3/n23 ) );
  INV_X2 \pool/pool/shift_row3/U10  ( .A(\pool/pool/pe_b_o_data[3][36] ), .ZN(
        \pool/pool/shift_row3/n24 ) );
  NAND2_X2 \pool/pool/shift_row3/U9  ( .A1(\pool/pool/pe_b_o_data[3][35] ), 
        .A2(\pool/pool/pe_b_o_data[3][34] ), .ZN(\pool/pool/shift_row3/n13 )
         );
  NOR2_X2 \pool/pool/shift_row3/U8  ( .A1(\pool/pool/shift_row3/n13 ), .A2(
        \pool/pool/shift_row3/n24 ), .ZN(\pool/pool/shift_row3/n14 ) );
  NAND2_X2 \pool/pool/shift_row3/U7  ( .A1(\pool/pool/pe_b_o_data[3][24] ), 
        .A2(\pool/pool/pe_b_o_data[3][23] ), .ZN(\pool/pool/shift_row3/n15 )
         );
  NOR2_X2 \pool/pool/shift_row3/U6  ( .A1(\pool/pool/shift_row3/n15 ), .A2(
        \pool/pool/shift_row3/n23 ), .ZN(\pool/pool/shift_row3/n16 ) );
  NAND2_X2 \pool/pool/shift_row3/U5  ( .A1(\pool/pool/pe_b_o_data[3][13] ), 
        .A2(\pool/pool/pe_b_o_data[3][12] ), .ZN(\pool/pool/shift_row3/n17 )
         );
  NOR2_X2 \pool/pool/shift_row3/U4  ( .A1(\pool/pool/shift_row3/n17 ), .A2(
        \pool/pool/shift_row3/n22 ), .ZN(\pool/pool/shift_row3/n18 ) );
  NAND2_X2 \pool/pool/shift_row3/U3  ( .A1(\pool/pool/pe_b_o_data[3][2] ), 
        .A2(\pool/pool/pe_b_o_data[3][1] ), .ZN(\pool/pool/shift_row3/n19 ) );
  NOR2_X2 \pool/pool/shift_row3/U2  ( .A1(\pool/pool/shift_row3/n19 ), .A2(
        \pool/pool/shift_row3/n21 ), .ZN(\pool/pool/shift_row3/n20 ) );
  INV_X1 \pool/fsm/U27  ( .A(\pool/fsm/N11 ), .ZN(\pool/fsm/n17 ) );
  INV_X1 \pool/fsm/U26  ( .A(\pool/fsm/n17 ), .ZN(\pool/ld_h ) );
  INV_X2 \pool/fsm/U20  ( .A(\pool/fsm/n18 ), .ZN(\pool/fsm/n4 ) );
  INV_X1 \pool/fsm/U16  ( .A(\pool/fsm/n4 ), .ZN(\pool/sel ) );
  NAND3_X1 \pool/fsm/U25  ( .A1(\pool/fsm/n8 ), .A2(\pool/fsm/n6 ), .A3(
        \pool/fsm/current_state[0] ), .ZN(\pool/fsm/n12 ) );
  NAND3_X1 \pool/fsm/U24  ( .A1(\pool/fsm/n9 ), .A2(\pool/fsm/n8 ), .A3(
        \pool/fsm/current_state[2] ), .ZN(\pool/fsm/n15 ) );
  NAND3_X1 \pool/fsm/U23  ( .A1(\pool/fsm/n12 ), .A2(\pool/fsm/n15 ), .A3(
        \pool/fsm/n5 ), .ZN(\pool/fsm/N29 ) );
  NAND3_X1 \pool/fsm/U22  ( .A1(\pool/sel ), .A2(\pool/fsm/n10 ), .A3(
        \pool/tc ), .ZN(\pool/fsm/n13 ) );
  INV_X2 \pool/fsm/U21  ( .A(done), .ZN(\pool/fsm/n10 ) );
  INV_X2 \pool/fsm/U19  ( .A(\pool/fsm/n16 ), .ZN(\pool/fsm/n5 ) );
  INV_X2 \pool/fsm/U18  ( .A(\pool/fsm/n11 ), .ZN(\pool/rst_cnt ) );
  INV_X2 \pool/fsm/U17  ( .A(\pool/sync_clr ), .ZN(\pool/fsm/n3 ) );
  NOR3_X2 \pool/fsm/U15  ( .A1(\pool/fsm/current_state[1] ), .A2(
        \pool/fsm/current_state[2] ), .A3(\pool/fsm/current_state[0] ), .ZN(
        \pool/fsm/N11 ) );
  NOR3_X2 \pool/fsm/U14  ( .A1(\pool/fsm/n9 ), .A2(\pool/fsm/current_state[2] ), .A3(\pool/fsm/n8 ), .ZN(\pool/fsm/n16 ) );
  NAND2_X2 \pool/fsm/U13  ( .A1(\pool/fsm/n17 ), .A2(\pool/fsm/n15 ), .ZN(
        \pool/sync_clr ) );
  NOR2_X2 \pool/fsm/U12  ( .A1(\pool/fsm/n16 ), .A2(\pool/sync_clr ), .ZN(
        \pool/fsm/n11 ) );
  NAND2_X2 \pool/fsm/U11  ( .A1(\pool/fsm/n12 ), .A2(\pool/fsm/n11 ), .ZN(
        \pool/fsm/N28 ) );
  OR2_X2 \pool/fsm/U10  ( .A1(start), .A2(\pool/fsm/n17 ), .ZN(\pool/fsm/N31 )
         );
  NOR3_X2 \pool/fsm/U9  ( .A1(\pool/fsm/current_state[0] ), .A2(
        \pool/fsm/current_state[2] ), .A3(\pool/fsm/n8 ), .ZN(\pool/fsm/n18 )
         );
  NAND2_X2 \pool/fsm/U8  ( .A1(\pool/fsm/n12 ), .A2(\pool/fsm/n4 ), .ZN(
        \pool/en_cnt ) );
  AND2_X2 \pool/fsm/U7  ( .A1(\pool/tc ), .A2(done), .ZN(\pool/fsm/n14 ) );
  OAI21_X2 \pool/fsm/U6  ( .B1(\pool/fsm/n14 ), .B2(\pool/fsm/n4 ), .A(
        \pool/fsm/n3 ), .ZN(\pool/fsm/next_state [0]) );
  NAND2_X2 \pool/fsm/U5  ( .A1(\pool/fsm/n12 ), .A2(\pool/fsm/n13 ), .ZN(
        \pool/fsm/next_state [1]) );
  OR2_X2 \pool/fsm/U4  ( .A1(\pool/sel ), .A2(\pool/fsm/N29 ), .ZN(
        \pool/rst_cnt_c ) );
  INV_X1 \pool/fsm/U3  ( .A(rst_fsm), .ZN(\pool/fsm/n1 ) );
  DLH_X1 \pool/fsm/rst_cnt_r_reg  ( .G(\pool/fsm/N28 ), .D(\pool/fsm/N29 ), 
        .Q(\pool/rst_cnt_r ) );
  DFFR_X1 \pool/fsm/current_state_reg[2]  ( .D(\pool/fsm/n16 ), .CK(
        \pool/fsm/net468 ), .RN(\pool/fsm/n1 ), .Q(\pool/fsm/current_state[2] ), .QN(\pool/fsm/n6 ) );
  DFFR_X1 \pool/fsm/current_state_reg[1]  ( .D(\pool/fsm/next_state [1]), .CK(
        \pool/fsm/net468 ), .RN(\pool/fsm/n1 ), .Q(\pool/fsm/current_state[1] ), .QN(\pool/fsm/n8 ) );
  DFFR_X1 \pool/fsm/current_state_reg[0]  ( .D(\pool/fsm/next_state [0]), .CK(
        \pool/fsm/net468 ), .RN(\pool/fsm/n1 ), .Q(\pool/fsm/current_state[0] ), .QN(\pool/fsm/n9 ) );
  SNPS_CLOCK_GATE_HIGH_avr_pooling_fsm \pool/fsm/clk_gate_current_state_reg  ( 
        .CLK(clk), .EN(\pool/fsm/N31 ), .ENCLK(\pool/fsm/net468 ), .TE(1'b0)
         );
  INV_X1 \pool/gate_clk/U37  ( .A(\pool/ld_h ), .ZN(\pool/gate_clk/n32 ) );
  INV_X1 \pool/gate_clk/U36  ( .A(\pool/ld_h ), .ZN(\pool/gate_clk/n31 ) );
  INV_X1 \pool/gate_clk/U35  ( .A(\pool/gate_clk/n32 ), .ZN(
        \pool/gate_clk/n30 ) );
  INV_X1 \pool/gate_clk/U32  ( .A(\pool/ld_h ), .ZN(\pool/gate_clk/n14 ) );
  INV_X1 \pool/gate_clk/U31  ( .A(\pool/gate_clk/n14 ), .ZN(
        \pool/gate_clk/n13 ) );
  AND2_X1 \pool/gate_clk/U4  ( .A1(\pool/gate_clk/del_tc_r ), .A2(
        \pool/gate_clk/n14 ), .ZN(\pool/gate_clk/n2 ) );
  AND2_X1 \pool/gate_clk/U3  ( .A1(\pool/gate_clk/del_0_tc ), .A2(
        \pool/gate_clk/n14 ), .ZN(\pool/gate_clk/n1 ) );
  DFF_X1 \pool/gate_clk/del_1_tc_reg  ( .D(\pool/gate_clk/n1 ), .CK(clk), .Q(
        \pool/gate_clk/del_1_tc ) );
  DFF_X1 \pool/gate_clk/del_tc_r_1_reg  ( .D(\pool/gate_clk/n2 ), .CK(clk), 
        .Q(\pool/gate_clk/del_tc_r_1 ) );
  NAND3_X1 \pool/gate_clk/U34  ( .A1(\pool/gate_clk/cnt_c_out[1] ), .A2(
        \pool/gate_clk/n32 ), .A3(\pool/gate_clk/cnt_c_out[0] ), .ZN(
        \pool/gate_clk/n23 ) );
  INV_X2 \pool/gate_clk/U33  ( .A(\pool/rst_cnt_c ), .ZN(\pool/gate_clk/n15 )
         );
  INV_X2 \pool/gate_clk/U30  ( .A(\pool/tc ), .ZN(\pool/gate_clk/n12 ) );
  INV_X2 \pool/gate_clk/U29  ( .A(\pool/gate_clk/tc_c ), .ZN(
        \pool/gate_clk/n8 ) );
  INV_X2 \pool/gate_clk/U28  ( .A(\pool/gate_clk/n21 ), .ZN(\pool/gate_clk/n7 ) );
  INV_X2 \pool/gate_clk/U27  ( .A(\pool/gate_clk/pool_size[4] ), .ZN(
        \pool/gate_clk/n6 ) );
  INV_X2 \pool/gate_clk/U26  ( .A(\pool/gate_clk/pool_size[3] ), .ZN(
        \pool/gate_clk/n5 ) );
  INV_X2 \pool/gate_clk/U25  ( .A(\pool/gate_clk/pool_size[0] ), .ZN(
        \pool/gate_clk/n4 ) );
  INV_X2 \pool/gate_clk/U24  ( .A(\pool/gate_clk/dec_out[1] ), .ZN(
        \pool/gate_clk/n3 ) );
  NOR2_X2 \pool/gate_clk/U23  ( .A1(\pool/gate_clk/n13 ), .A2(
        \pool/gate_clk/n12 ), .ZN(\pool/gate_clk/N21 ) );
  NOR3_X2 \pool/gate_clk/U22  ( .A1(\pool/gate_clk/cnt_r_out[0] ), .A2(
        \pool/gate_clk/n13 ), .A3(\pool/gate_clk/cnt_r_out[1] ), .ZN(
        \pool/gate_clk/N45 ) );
  NOR2_X2 \pool/gate_clk/U21  ( .A1(\pool/gate_clk/pool_size[2] ), .A2(
        \pool/gate_clk/n4 ), .ZN(\pool/gate_clk/dec_out[1] ) );
  OAI21_X2 \pool/gate_clk/U20  ( .B1(\pool/gate_clk/pool_size[1] ), .B2(
        \pool/gate_clk/n4 ), .A(\pool/gate_clk/n3 ), .ZN(
        \pool/gate_clk/dec_out[0] ) );
  NOR2_X2 \pool/gate_clk/U19  ( .A1(\pool/gate_clk/pool_size[1] ), .A2(
        \pool/gate_clk/n3 ), .ZN(\pool/gate_clk/dec_out[2] ) );
  NOR3_X2 \pool/gate_clk/U18  ( .A1(\pool/gate_clk/n30 ), .A2(
        \pool/gate_clk/del_1_tc ), .A3(\pool/gate_clk/n15 ), .ZN(
        \pool/gate_clk/n21 ) );
  AOI221_X2 \pool/gate_clk/U17  ( .B1(\pool/gate_clk/n10 ), .B2(
        \pool/gate_clk/n32 ), .C1(\pool/gate_clk/pool_size[3] ), .C2(
        \pool/gate_clk/n30 ), .A(\pool/gate_clk/n15 ), .ZN(\pool/gate_clk/n25 ) );
  OAI22_X2 \pool/gate_clk/U16  ( .A1(\pool/gate_clk/n10 ), .A2(
        \pool/gate_clk/n7 ), .B1(\pool/gate_clk/n21 ), .B2(\pool/gate_clk/n25 ), .ZN(\pool/gate_clk/n29 ) );
  NOR3_X2 \pool/gate_clk/U15  ( .A1(\pool/gate_clk/cnt_c_out[0] ), .A2(
        \pool/gate_clk/n30 ), .A3(\pool/gate_clk/cnt_c_out[1] ), .ZN(
        \pool/gate_clk/n24 ) );
  AOI211_X2 \pool/gate_clk/U14  ( .C1(\pool/gate_clk/pool_size[4] ), .C2(
        \pool/gate_clk/n30 ), .A(\pool/gate_clk/n15 ), .B(\pool/gate_clk/n24 ), 
        .ZN(\pool/gate_clk/n22 ) );
  OAI221_X2 \pool/gate_clk/U13  ( .B1(\pool/gate_clk/n21 ), .B2(
        \pool/gate_clk/n22 ), .C1(\pool/gate_clk/n9 ), .C2(\pool/gate_clk/n7 ), 
        .A(\pool/gate_clk/n23 ), .ZN(\pool/gate_clk/n28 ) );
  NOR2_X2 \pool/gate_clk/U12  ( .A1(\pool/gate_clk/cnt_c_out[0] ), .A2(
        \pool/gate_clk/cnt_c_out[1] ), .ZN(\pool/gate_clk/tc_c ) );
  NAND2_X2 \pool/gate_clk/U11  ( .A1(\pool/tc ), .A2(\pool/gate_clk/tc_c ), 
        .ZN(\pool/gate_clk/n19 ) );
  NOR3_X2 \pool/gate_clk/U10  ( .A1(\pool/gate_clk/n8 ), .A2(
        \pool/gate_clk/cnt_r_out[0] ), .A3(\pool/gate_clk/n12 ), .ZN(
        \pool/gate_clk/n18 ) );
  AOI21_X2 \pool/gate_clk/U9  ( .B1(\pool/gate_clk/cnt_r_out[0] ), .B2(
        \pool/gate_clk/n19 ), .A(\pool/gate_clk/n18 ), .ZN(\pool/gate_clk/n20 ) );
  OAI221_X2 \pool/gate_clk/U8  ( .B1(\pool/gate_clk/n31 ), .B2(
        \pool/gate_clk/n5 ), .C1(\pool/gate_clk/n30 ), .C2(\pool/gate_clk/n20 ), .A(\pool/rst_cnt_r ), .ZN(\pool/gate_clk/n27 ) );
  OR2_X2 \pool/gate_clk/U7  ( .A1(\pool/gate_clk/cnt_r_out[0] ), .A2(
        \pool/gate_clk/n19 ), .ZN(\pool/gate_clk/n17 ) );
  AOI22_X2 \pool/gate_clk/U6  ( .A1(\pool/gate_clk/cnt_r_out[1] ), .A2(
        \pool/gate_clk/n17 ), .B1(\pool/gate_clk/n18 ), .B2(
        \pool/gate_clk/n11 ), .ZN(\pool/gate_clk/n16 ) );
  OAI221_X2 \pool/gate_clk/U5  ( .B1(\pool/gate_clk/n31 ), .B2(
        \pool/gate_clk/n6 ), .C1(\pool/gate_clk/n30 ), .C2(\pool/gate_clk/n16 ), .A(\pool/rst_cnt_r ), .ZN(\pool/gate_clk/n26 ) );
  DFF_X1 \pool/gate_clk/del_tc_r_reg  ( .D(\pool/gate_clk/N45 ), .CK(clk), .Q(
        \pool/gate_clk/del_tc_r ) );
  DFF_X1 \pool/gate_clk/cnt_r_out_reg[1]  ( .D(\pool/gate_clk/n26 ), .CK(clk), 
        .Q(\pool/gate_clk/cnt_r_out[1] ), .QN(\pool/gate_clk/n11 ) );
  DFF_X1 \pool/gate_clk/cnt_r_out_reg[0]  ( .D(\pool/gate_clk/n27 ), .CK(clk), 
        .Q(\pool/gate_clk/cnt_r_out[0] ) );
  DFF_X1 \pool/gate_clk/cnt_c_out_reg[1]  ( .D(\pool/gate_clk/n28 ), .CK(clk), 
        .Q(\pool/gate_clk/cnt_c_out[1] ), .QN(\pool/gate_clk/n9 ) );
  DFF_X1 \pool/gate_clk/cnt_c_out_reg[0]  ( .D(\pool/gate_clk/n29 ), .CK(clk), 
        .Q(\pool/gate_clk/cnt_c_out[0] ), .QN(\pool/gate_clk/n10 ) );
  DFF_X1 \pool/gate_clk/del_0_tc_reg  ( .D(\pool/gate_clk/N21 ), .CK(clk), .Q(
        \pool/gate_clk/del_0_tc ) );
  INV_X2 \pool/gate_clk/mux_pool/U11  ( .A(pool_sel), .ZN(
        \pool/gate_clk/mux_pool/n6 ) );
  INV_X2 \pool/gate_clk/mux_pool/U10  ( .A(\pool/gate_clk/mux_pool/n11 ), .ZN(
        \pool/gate_clk/pool_size[0] ) );
  INV_X2 \pool/gate_clk/mux_pool/U9  ( .A(\pool/gate_clk/mux_pool/n10 ), .ZN(
        \pool/gate_clk/pool_size[1] ) );
  INV_X2 \pool/gate_clk/mux_pool/U8  ( .A(\pool/gate_clk/mux_pool/n9 ), .ZN(
        \pool/gate_clk/pool_size[2] ) );
  INV_X2 \pool/gate_clk/mux_pool/U7  ( .A(\pool/gate_clk/mux_pool/n8 ), .ZN(
        \pool/gate_clk/pool_size[3] ) );
  INV_X2 \pool/gate_clk/mux_pool/U6  ( .A(\pool/gate_clk/mux_pool/n7 ), .ZN(
        \pool/gate_clk/pool_size[4] ) );
  AOI22_X2 \pool/gate_clk/mux_pool/U5  ( .A1(size_1[0]), .A2(
        \pool/gate_clk/mux_pool/n6 ), .B1(size_2[0]), .B2(pool_sel), .ZN(
        \pool/gate_clk/mux_pool/n11 ) );
  AOI22_X2 \pool/gate_clk/mux_pool/U4  ( .A1(size_1[1]), .A2(
        \pool/gate_clk/mux_pool/n6 ), .B1(size_2[1]), .B2(pool_sel), .ZN(
        \pool/gate_clk/mux_pool/n10 ) );
  AOI22_X2 \pool/gate_clk/mux_pool/U3  ( .A1(size_1[2]), .A2(
        \pool/gate_clk/mux_pool/n6 ), .B1(size_2[2]), .B2(pool_sel), .ZN(
        \pool/gate_clk/mux_pool/n9 ) );
  AOI22_X2 \pool/gate_clk/mux_pool/U2  ( .A1(size_1[3]), .A2(
        \pool/gate_clk/mux_pool/n6 ), .B1(size_2[3]), .B2(pool_sel), .ZN(
        \pool/gate_clk/mux_pool/n8 ) );
  AOI22_X2 \pool/gate_clk/mux_pool/U1  ( .A1(size_1[4]), .A2(
        \pool/gate_clk/mux_pool/n6 ), .B1(pool_sel), .B2(size_2[4]), .ZN(
        \pool/gate_clk/mux_pool/n7 ) );
  INV_X2 \pool/gate_clk/mux_cmask/U9  ( .A(\pool/gate_clk/tc_c ), .ZN(
        \pool/gate_clk/mux_cmask/n5 ) );
  INV_X2 \pool/gate_clk/mux_cmask/U8  ( .A(\pool/gate_clk/mux_cmask/n9 ), .ZN(
        \pool/ckg_cmask [0]) );
  INV_X2 \pool/gate_clk/mux_cmask/U7  ( .A(\pool/gate_clk/mux_cmask/n8 ), .ZN(
        \pool/ckg_cmask [1]) );
  INV_X2 \pool/gate_clk/mux_cmask/U6  ( .A(\pool/gate_clk/mux_cmask/n7 ), .ZN(
        \pool/ckg_cmask [2]) );
  INV_X2 \pool/gate_clk/mux_cmask/U5  ( .A(\pool/gate_clk/mux_cmask/n6 ), .ZN(
        \pool/ckg_cmask [3]) );
  AOI22_X2 \pool/gate_clk/mux_cmask/U4  ( .A1(1'b0), .A2(
        \pool/gate_clk/mux_cmask/n5 ), .B1(\pool/gate_clk/dec_out[0] ), .B2(
        \pool/gate_clk/tc_c ), .ZN(\pool/gate_clk/mux_cmask/n9 ) );
  AOI22_X2 \pool/gate_clk/mux_cmask/U3  ( .A1(1'b0), .A2(
        \pool/gate_clk/mux_cmask/n5 ), .B1(\pool/gate_clk/dec_out[1] ), .B2(
        \pool/gate_clk/tc_c ), .ZN(\pool/gate_clk/mux_cmask/n8 ) );
  AOI22_X2 \pool/gate_clk/mux_cmask/U2  ( .A1(1'b0), .A2(
        \pool/gate_clk/mux_cmask/n5 ), .B1(\pool/gate_clk/dec_out[2] ), .B2(
        \pool/gate_clk/tc_c ), .ZN(\pool/gate_clk/mux_cmask/n7 ) );
  AOI22_X2 \pool/gate_clk/mux_cmask/U1  ( .A1(1'b0), .A2(
        \pool/gate_clk/mux_cmask/n5 ), .B1(\pool/gate_clk/tc_c ), .B2(1'b0), 
        .ZN(\pool/gate_clk/mux_cmask/n6 ) );
  INV_X2 \pool/gate_clk/mux_rmask/U9  ( .A(\pool/gate_clk/del_tc_r_1 ), .ZN(
        \pool/gate_clk/mux_rmask/n6 ) );
  INV_X2 \pool/gate_clk/mux_rmask/U8  ( .A(\pool/gate_clk/mux_rmask/n1 ), .ZN(
        \pool/ckg_rmask [0]) );
  INV_X2 \pool/gate_clk/mux_rmask/U7  ( .A(\pool/gate_clk/mux_rmask/n2 ), .ZN(
        \pool/ckg_rmask [1]) );
  INV_X2 \pool/gate_clk/mux_rmask/U6  ( .A(\pool/gate_clk/mux_rmask/n3 ), .ZN(
        \pool/ckg_rmask [2]) );
  INV_X2 \pool/gate_clk/mux_rmask/U5  ( .A(\pool/gate_clk/mux_rmask/n4 ), .ZN(
        \pool/ckg_rmask [3]) );
  AOI22_X2 \pool/gate_clk/mux_rmask/U4  ( .A1(1'b0), .A2(
        \pool/gate_clk/mux_rmask/n6 ), .B1(\pool/gate_clk/dec_out[0] ), .B2(
        \pool/gate_clk/del_tc_r_1 ), .ZN(\pool/gate_clk/mux_rmask/n1 ) );
  AOI22_X2 \pool/gate_clk/mux_rmask/U3  ( .A1(1'b0), .A2(
        \pool/gate_clk/mux_rmask/n6 ), .B1(\pool/gate_clk/dec_out[1] ), .B2(
        \pool/gate_clk/del_tc_r_1 ), .ZN(\pool/gate_clk/mux_rmask/n2 ) );
  AOI22_X2 \pool/gate_clk/mux_rmask/U2  ( .A1(1'b0), .A2(
        \pool/gate_clk/mux_rmask/n6 ), .B1(\pool/gate_clk/dec_out[2] ), .B2(
        \pool/gate_clk/del_tc_r_1 ), .ZN(\pool/gate_clk/mux_rmask/n3 ) );
  AOI22_X2 \pool/gate_clk/mux_rmask/U1  ( .A1(1'b0), .A2(
        \pool/gate_clk/mux_rmask/n6 ), .B1(\pool/gate_clk/del_tc_r_1 ), .B2(
        1'b0), .ZN(\pool/gate_clk/mux_rmask/n4 ) );
endmodule

