
module dp ( ck, rst, i_acth, i_actv, i_weight, arv_ckg, arv_k, arv_i_tile, 
        arv_o_tile, arv_ifmaps, arv_ofmaps, ctrl_en_npu, ctrl_ldh_v_n, 
        ctrl_en_hmode, ctrl_en_vmode, ctrl_wr_pipe, ctrl_en_p, ctrl_wr_mem, 
        s_tc_hmode, s_tc_vmode, s_tc_res, s_tc_npu_ptr, s_tc_tilev, s_tc_tileh, 
        s_tc_ifmaps, s_tc_ofmaps, i_weight_addr, i_data_ev_odd_n, 
        i_data_even_addr, i_data_odd_addr, o_data_ev_odd_n, o_data_even_addr, 
        o_data_odd_addr, o_data_wr, o_data_wrh_l_n, o_data, o_data_relu );
  input [15:0] i_acth;
  input [15:0] i_actv;
  input [1:0] i_weight;
  input [2:0] arv_ckg;
  input [2:0] arv_k;
  input [1:0] arv_i_tile;
  input [1:0] arv_o_tile;
  input [2:0] arv_ifmaps;
  input [3:0] arv_ofmaps;
  output [15:0] i_weight_addr;
  output [9:0] i_data_even_addr;
  output [9:0] i_data_odd_addr;
  output [9:0] o_data_even_addr;
  output [9:0] o_data_odd_addr;
  output [7:0] o_data;
  output [15:0] o_data_relu;
  input ck, rst, ctrl_en_npu, ctrl_ldh_v_n, ctrl_en_hmode, ctrl_en_vmode,
         ctrl_wr_pipe, ctrl_en_p, ctrl_wr_mem;
  output s_tc_hmode, s_tc_vmode, s_tc_res, s_tc_npu_ptr, s_tc_tilev,
         s_tc_tileh, s_tc_ifmaps, s_tc_ofmaps, i_data_ev_odd_n,
         o_data_ev_odd_n, o_data_wr, o_data_wrh_l_n;
  wire   ps_ctrl_en_npu, ps_ctrl_ldh_v_n, ps_ctrl_wr_pipe, ps_ctrl_en_p,
         int_en_hmode, int_en_vmode, int_en_npu_ptr, int_en_tilev_ptr,
         int_en_ofmaps_ptr, int_tileh_ptr_1_, int_c_i_en_weight_addr,
         int_c_i_en_even, int_c_i_en_odd, ps_int_s_tc_res, ps_int_s_tc_tilev,
         ps_int_s_tc_tileh, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N100, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123,
         N124, N125, net2747, net2753, net2758, net2763, n16, n19, n21, n26,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         wrap_act_buffer_inst_n2, wrap_act_buffer_inst_n1,
         wrap_act_buffer_inst_net4501,
         wrap_act_buffer_inst_act_buffer_inst_n267,
         wrap_act_buffer_inst_act_buffer_inst_n266,
         wrap_act_buffer_inst_act_buffer_inst_n265,
         wrap_act_buffer_inst_act_buffer_inst_n264,
         wrap_act_buffer_inst_act_buffer_inst_n263,
         wrap_act_buffer_inst_act_buffer_inst_n262,
         wrap_act_buffer_inst_act_buffer_inst_n261,
         wrap_act_buffer_inst_act_buffer_inst_n260,
         wrap_act_buffer_inst_act_buffer_inst_n259,
         wrap_act_buffer_inst_act_buffer_inst_n258,
         wrap_act_buffer_inst_act_buffer_inst_n257,
         wrap_act_buffer_inst_act_buffer_inst_n256,
         wrap_act_buffer_inst_act_buffer_inst_n255,
         wrap_act_buffer_inst_act_buffer_inst_n254,
         wrap_act_buffer_inst_act_buffer_inst_n253,
         wrap_act_buffer_inst_act_buffer_inst_n252,
         wrap_act_buffer_inst_act_buffer_inst_n251,
         wrap_act_buffer_inst_act_buffer_inst_n250,
         wrap_act_buffer_inst_act_buffer_inst_n249,
         wrap_act_buffer_inst_act_buffer_inst_n248,
         wrap_act_buffer_inst_act_buffer_inst_n247,
         wrap_act_buffer_inst_act_buffer_inst_n246,
         wrap_act_buffer_inst_act_buffer_inst_n245,
         wrap_act_buffer_inst_act_buffer_inst_n244,
         wrap_act_buffer_inst_act_buffer_inst_n243,
         wrap_act_buffer_inst_act_buffer_inst_n242,
         wrap_act_buffer_inst_act_buffer_inst_n241,
         wrap_act_buffer_inst_act_buffer_inst_n240,
         wrap_act_buffer_inst_act_buffer_inst_n239,
         wrap_act_buffer_inst_act_buffer_inst_n238,
         wrap_act_buffer_inst_act_buffer_inst_n237,
         wrap_act_buffer_inst_act_buffer_inst_n236,
         wrap_act_buffer_inst_act_buffer_inst_n235,
         wrap_act_buffer_inst_act_buffer_inst_n234,
         wrap_act_buffer_inst_act_buffer_inst_n233,
         wrap_act_buffer_inst_act_buffer_inst_n232,
         wrap_act_buffer_inst_act_buffer_inst_n231,
         wrap_act_buffer_inst_act_buffer_inst_n230,
         wrap_act_buffer_inst_act_buffer_inst_n229,
         wrap_act_buffer_inst_act_buffer_inst_n228,
         wrap_act_buffer_inst_act_buffer_inst_n227,
         wrap_act_buffer_inst_act_buffer_inst_n226,
         wrap_act_buffer_inst_act_buffer_inst_n225,
         wrap_act_buffer_inst_act_buffer_inst_n224,
         wrap_act_buffer_inst_act_buffer_inst_n223,
         wrap_act_buffer_inst_act_buffer_inst_n222,
         wrap_act_buffer_inst_act_buffer_inst_n221,
         wrap_act_buffer_inst_act_buffer_inst_n220,
         wrap_act_buffer_inst_act_buffer_inst_n219,
         wrap_act_buffer_inst_act_buffer_inst_n218,
         wrap_act_buffer_inst_act_buffer_inst_n217,
         wrap_act_buffer_inst_act_buffer_inst_n216,
         wrap_act_buffer_inst_act_buffer_inst_n215,
         wrap_act_buffer_inst_act_buffer_inst_n214,
         wrap_act_buffer_inst_act_buffer_inst_n213,
         wrap_act_buffer_inst_act_buffer_inst_n212,
         wrap_act_buffer_inst_act_buffer_inst_n211,
         wrap_act_buffer_inst_act_buffer_inst_n210,
         wrap_act_buffer_inst_act_buffer_inst_n209,
         wrap_act_buffer_inst_act_buffer_inst_n208,
         wrap_act_buffer_inst_act_buffer_inst_n207,
         wrap_act_buffer_inst_act_buffer_inst_n206,
         wrap_act_buffer_inst_act_buffer_inst_n205,
         wrap_act_buffer_inst_act_buffer_inst_n204,
         wrap_act_buffer_inst_act_buffer_inst_n203,
         wrap_act_buffer_inst_act_buffer_inst_n202,
         wrap_act_buffer_inst_act_buffer_inst_n201,
         wrap_act_buffer_inst_act_buffer_inst_n200,
         wrap_act_buffer_inst_act_buffer_inst_n199,
         wrap_act_buffer_inst_act_buffer_inst_n198,
         wrap_act_buffer_inst_act_buffer_inst_n197,
         wrap_act_buffer_inst_act_buffer_inst_n196,
         wrap_act_buffer_inst_act_buffer_inst_n195,
         wrap_act_buffer_inst_act_buffer_inst_n194,
         wrap_act_buffer_inst_act_buffer_inst_n193,
         wrap_act_buffer_inst_act_buffer_inst_n192,
         wrap_act_buffer_inst_act_buffer_inst_n191,
         wrap_act_buffer_inst_act_buffer_inst_n190,
         wrap_act_buffer_inst_act_buffer_inst_n189,
         wrap_act_buffer_inst_act_buffer_inst_n188,
         wrap_act_buffer_inst_act_buffer_inst_n187,
         wrap_act_buffer_inst_act_buffer_inst_n186,
         wrap_act_buffer_inst_act_buffer_inst_n185,
         wrap_act_buffer_inst_act_buffer_inst_n184,
         wrap_act_buffer_inst_act_buffer_inst_n183,
         wrap_act_buffer_inst_act_buffer_inst_n182,
         wrap_act_buffer_inst_act_buffer_inst_n181,
         wrap_act_buffer_inst_act_buffer_inst_n180,
         wrap_act_buffer_inst_act_buffer_inst_n179,
         wrap_act_buffer_inst_act_buffer_inst_n178,
         wrap_act_buffer_inst_act_buffer_inst_n177,
         wrap_act_buffer_inst_act_buffer_inst_n176,
         wrap_act_buffer_inst_act_buffer_inst_n175,
         wrap_act_buffer_inst_act_buffer_inst_n174,
         wrap_act_buffer_inst_act_buffer_inst_n173,
         wrap_act_buffer_inst_act_buffer_inst_n172,
         wrap_act_buffer_inst_act_buffer_inst_n171,
         wrap_act_buffer_inst_act_buffer_inst_n170,
         wrap_act_buffer_inst_act_buffer_inst_n169,
         wrap_act_buffer_inst_act_buffer_inst_n168,
         wrap_act_buffer_inst_act_buffer_inst_n167,
         wrap_act_buffer_inst_act_buffer_inst_n166,
         wrap_act_buffer_inst_act_buffer_inst_n165,
         wrap_act_buffer_inst_act_buffer_inst_n164,
         wrap_act_buffer_inst_act_buffer_inst_n163,
         wrap_act_buffer_inst_act_buffer_inst_n162,
         wrap_act_buffer_inst_act_buffer_inst_n161,
         wrap_act_buffer_inst_act_buffer_inst_n160,
         wrap_act_buffer_inst_act_buffer_inst_n159,
         wrap_act_buffer_inst_act_buffer_inst_n9,
         wrap_act_buffer_inst_act_buffer_inst_n8,
         wrap_act_buffer_inst_act_buffer_inst_n7,
         wrap_act_buffer_inst_act_buffer_inst_n6,
         wrap_act_buffer_inst_act_buffer_inst_n5,
         wrap_act_buffer_inst_act_buffer_inst_n4,
         wrap_act_buffer_inst_act_buffer_inst_n3,
         wrap_act_buffer_inst_act_buffer_inst_n2,
         wrap_act_buffer_inst_act_buffer_inst_n1,
         wrap_act_buffer_inst_act_buffer_inst_n158,
         wrap_act_buffer_inst_act_buffer_inst_n157,
         wrap_act_buffer_inst_act_buffer_inst_n156,
         wrap_act_buffer_inst_act_buffer_inst_n155,
         wrap_act_buffer_inst_act_buffer_inst_n154,
         wrap_act_buffer_inst_act_buffer_inst_n153,
         wrap_act_buffer_inst_act_buffer_inst_n152,
         wrap_act_buffer_inst_act_buffer_inst_n151,
         wrap_act_buffer_inst_act_buffer_inst_n150,
         wrap_act_buffer_inst_act_buffer_inst_n149,
         wrap_act_buffer_inst_act_buffer_inst_n148,
         wrap_act_buffer_inst_act_buffer_inst_n147,
         wrap_act_buffer_inst_act_buffer_inst_n146,
         wrap_act_buffer_inst_act_buffer_inst_n145,
         wrap_act_buffer_inst_act_buffer_inst_n144,
         wrap_act_buffer_inst_act_buffer_inst_n143,
         wrap_act_buffer_inst_act_buffer_inst_n142,
         wrap_act_buffer_inst_act_buffer_inst_n141,
         wrap_act_buffer_inst_act_buffer_inst_n140,
         wrap_act_buffer_inst_act_buffer_inst_n139,
         wrap_act_buffer_inst_act_buffer_inst_n138,
         wrap_act_buffer_inst_act_buffer_inst_n137,
         wrap_act_buffer_inst_act_buffer_inst_n136,
         wrap_act_buffer_inst_act_buffer_inst_n135,
         wrap_act_buffer_inst_act_buffer_inst_n134,
         wrap_act_buffer_inst_act_buffer_inst_n133,
         wrap_act_buffer_inst_act_buffer_inst_n132,
         wrap_act_buffer_inst_act_buffer_inst_n131,
         wrap_act_buffer_inst_act_buffer_inst_n130,
         wrap_act_buffer_inst_act_buffer_inst_n129,
         wrap_act_buffer_inst_act_buffer_inst_n128,
         wrap_act_buffer_inst_act_buffer_inst_n127,
         wrap_act_buffer_inst_act_buffer_inst_n126,
         wrap_act_buffer_inst_act_buffer_inst_n125,
         wrap_act_buffer_inst_act_buffer_inst_n124,
         wrap_act_buffer_inst_act_buffer_inst_n123,
         wrap_act_buffer_inst_act_buffer_inst_n122,
         wrap_act_buffer_inst_act_buffer_inst_n121,
         wrap_act_buffer_inst_act_buffer_inst_n120,
         wrap_act_buffer_inst_act_buffer_inst_n119,
         wrap_act_buffer_inst_act_buffer_inst_n118,
         wrap_act_buffer_inst_act_buffer_inst_n117,
         wrap_act_buffer_inst_act_buffer_inst_n116,
         wrap_act_buffer_inst_act_buffer_inst_n115,
         wrap_act_buffer_inst_act_buffer_inst_n114,
         wrap_act_buffer_inst_act_buffer_inst_n113,
         wrap_act_buffer_inst_act_buffer_inst_n112,
         wrap_act_buffer_inst_act_buffer_inst_n111,
         wrap_act_buffer_inst_act_buffer_inst_n110,
         wrap_act_buffer_inst_act_buffer_inst_n109,
         wrap_act_buffer_inst_act_buffer_inst_n108,
         wrap_act_buffer_inst_act_buffer_inst_n107,
         wrap_act_buffer_inst_act_buffer_inst_n106,
         wrap_act_buffer_inst_act_buffer_inst_n105,
         wrap_act_buffer_inst_act_buffer_inst_n104,
         wrap_act_buffer_inst_act_buffer_inst_n103,
         wrap_act_buffer_inst_act_buffer_inst_n102,
         wrap_act_buffer_inst_act_buffer_inst_n101,
         wrap_act_buffer_inst_act_buffer_inst_n100,
         wrap_act_buffer_inst_act_buffer_inst_n99,
         wrap_act_buffer_inst_act_buffer_inst_n98,
         wrap_act_buffer_inst_act_buffer_inst_n97,
         wrap_act_buffer_inst_act_buffer_inst_n96,
         wrap_act_buffer_inst_act_buffer_inst_n95,
         wrap_act_buffer_inst_act_buffer_inst_n94,
         wrap_act_buffer_inst_act_buffer_inst_n93,
         wrap_act_buffer_inst_act_buffer_inst_n92,
         wrap_act_buffer_inst_act_buffer_inst_n91,
         wrap_act_buffer_inst_act_buffer_inst_n90,
         wrap_act_buffer_inst_act_buffer_inst_n89,
         wrap_act_buffer_inst_act_buffer_inst_n88,
         wrap_act_buffer_inst_act_buffer_inst_n87,
         wrap_act_buffer_inst_act_buffer_inst_n86,
         wrap_act_buffer_inst_act_buffer_inst_n85,
         wrap_act_buffer_inst_act_buffer_inst_n84,
         wrap_act_buffer_inst_act_buffer_inst_n83,
         wrap_act_buffer_inst_act_buffer_inst_n82,
         wrap_act_buffer_inst_act_buffer_inst_n81,
         wrap_act_buffer_inst_act_buffer_inst_n80,
         wrap_act_buffer_inst_act_buffer_inst_n79,
         wrap_act_buffer_inst_act_buffer_inst_n78,
         wrap_act_buffer_inst_act_buffer_inst_n77,
         wrap_act_buffer_inst_act_buffer_inst_n76,
         wrap_act_buffer_inst_act_buffer_inst_n75,
         wrap_act_buffer_inst_act_buffer_inst_n74,
         wrap_act_buffer_inst_act_buffer_inst_n73,
         wrap_act_buffer_inst_act_buffer_inst_n72,
         wrap_act_buffer_inst_act_buffer_inst_n71,
         wrap_act_buffer_inst_act_buffer_inst_n70,
         wrap_act_buffer_inst_act_buffer_inst_n69,
         wrap_act_buffer_inst_act_buffer_inst_n68,
         wrap_act_buffer_inst_act_buffer_inst_n67,
         wrap_act_buffer_inst_act_buffer_inst_n66,
         wrap_act_buffer_inst_act_buffer_inst_n65,
         wrap_act_buffer_inst_act_buffer_inst_n64,
         wrap_act_buffer_inst_act_buffer_inst_n63,
         wrap_act_buffer_inst_act_buffer_inst_n62,
         wrap_act_buffer_inst_act_buffer_inst_n61,
         wrap_act_buffer_inst_act_buffer_inst_n60,
         wrap_act_buffer_inst_act_buffer_inst_n59,
         wrap_act_buffer_inst_act_buffer_inst_n58,
         wrap_act_buffer_inst_act_buffer_inst_n57,
         wrap_act_buffer_inst_act_buffer_inst_n56,
         wrap_act_buffer_inst_act_buffer_inst_n55,
         wrap_act_buffer_inst_act_buffer_inst_n54,
         wrap_act_buffer_inst_act_buffer_inst_n53,
         wrap_act_buffer_inst_act_buffer_inst_n52,
         wrap_act_buffer_inst_act_buffer_inst_n51,
         wrap_act_buffer_inst_act_buffer_inst_n50,
         wrap_act_buffer_inst_act_buffer_inst_n49,
         wrap_act_buffer_inst_act_buffer_inst_n48,
         wrap_act_buffer_inst_act_buffer_inst_n47,
         wrap_act_buffer_inst_act_buffer_inst_n46,
         wrap_act_buffer_inst_act_buffer_inst_n45,
         wrap_act_buffer_inst_act_buffer_inst_n44,
         wrap_act_buffer_inst_act_buffer_inst_n43,
         wrap_act_buffer_inst_act_buffer_inst_n42,
         wrap_act_buffer_inst_act_buffer_inst_n41,
         wrap_act_buffer_inst_act_buffer_inst_n40,
         wrap_act_buffer_inst_act_buffer_inst_n39,
         wrap_act_buffer_inst_act_buffer_inst_n38,
         wrap_act_buffer_inst_act_buffer_inst_n37,
         wrap_act_buffer_inst_act_buffer_inst_n36,
         wrap_act_buffer_inst_act_buffer_inst_n35,
         wrap_act_buffer_inst_act_buffer_inst_n34,
         wrap_act_buffer_inst_act_buffer_inst_n33,
         wrap_act_buffer_inst_act_buffer_inst_n32,
         wrap_act_buffer_inst_act_buffer_inst_n31,
         wrap_act_buffer_inst_act_buffer_inst_n30,
         wrap_act_buffer_inst_act_buffer_inst_n29,
         wrap_act_buffer_inst_act_buffer_inst_n28,
         wrap_act_buffer_inst_act_buffer_inst_n27,
         wrap_act_buffer_inst_act_buffer_inst_n26,
         wrap_act_buffer_inst_act_buffer_inst_n25,
         wrap_act_buffer_inst_act_buffer_inst_n24,
         wrap_act_buffer_inst_act_buffer_inst_n23,
         wrap_act_buffer_inst_act_buffer_inst_n22,
         wrap_act_buffer_inst_act_buffer_inst_n21,
         wrap_act_buffer_inst_act_buffer_inst_n20,
         wrap_act_buffer_inst_act_buffer_inst_n19,
         wrap_act_buffer_inst_act_buffer_inst_n18,
         wrap_act_buffer_inst_act_buffer_inst_n17,
         wrap_act_buffer_inst_act_buffer_inst_n16,
         wrap_act_buffer_inst_act_buffer_inst_n15,
         wrap_act_buffer_inst_act_buffer_inst_n14,
         wrap_act_buffer_inst_act_buffer_inst_n13,
         wrap_act_buffer_inst_act_buffer_inst_n12,
         wrap_act_buffer_inst_act_buffer_inst_n11,
         wrap_act_buffer_inst_act_buffer_inst_n10,
         wrap_act_buffer_inst_act_buffer_inst_net4755,
         wrap_act_buffer_inst_act_buffer_inst_net4750,
         wrap_act_buffer_inst_act_buffer_inst_net4745,
         wrap_act_buffer_inst_act_buffer_inst_net4740,
         wrap_act_buffer_inst_act_buffer_inst_net4735,
         wrap_act_buffer_inst_act_buffer_inst_net4730,
         wrap_act_buffer_inst_act_buffer_inst_net4725,
         wrap_act_buffer_inst_act_buffer_inst_net4720,
         wrap_act_buffer_inst_act_buffer_inst_net4715,
         wrap_act_buffer_inst_act_buffer_inst_net4710,
         wrap_act_buffer_inst_act_buffer_inst_net4705,
         wrap_act_buffer_inst_act_buffer_inst_net4700,
         wrap_act_buffer_inst_act_buffer_inst_net4695,
         wrap_act_buffer_inst_act_buffer_inst_net4690,
         wrap_act_buffer_inst_act_buffer_inst_net4685,
         wrap_act_buffer_inst_act_buffer_inst_net4680,
         wrap_act_buffer_inst_act_buffer_inst_net4675,
         wrap_act_buffer_inst_act_buffer_inst_net4670,
         wrap_act_buffer_inst_act_buffer_inst_net4665,
         wrap_act_buffer_inst_act_buffer_inst_net4660,
         wrap_act_buffer_inst_act_buffer_inst_net4655,
         wrap_act_buffer_inst_act_buffer_inst_net4650,
         wrap_act_buffer_inst_act_buffer_inst_net4645,
         wrap_act_buffer_inst_act_buffer_inst_net4640,
         wrap_act_buffer_inst_act_buffer_inst_net4635,
         wrap_act_buffer_inst_act_buffer_inst_net4630,
         wrap_act_buffer_inst_act_buffer_inst_net4625,
         wrap_act_buffer_inst_act_buffer_inst_net4620,
         wrap_act_buffer_inst_act_buffer_inst_net4615,
         wrap_act_buffer_inst_act_buffer_inst_net4610,
         wrap_act_buffer_inst_act_buffer_inst_net4605,
         wrap_act_buffer_inst_act_buffer_inst_net4600,
         wrap_act_buffer_inst_act_buffer_inst_net4595,
         wrap_act_buffer_inst_act_buffer_inst_net4590,
         wrap_act_buffer_inst_act_buffer_inst_net4585,
         wrap_act_buffer_inst_act_buffer_inst_net4580,
         wrap_act_buffer_inst_act_buffer_inst_net4575,
         wrap_act_buffer_inst_act_buffer_inst_net4570,
         wrap_act_buffer_inst_act_buffer_inst_net4565,
         wrap_act_buffer_inst_act_buffer_inst_net4560,
         wrap_act_buffer_inst_act_buffer_inst_net4555,
         wrap_act_buffer_inst_act_buffer_inst_net4550,
         wrap_act_buffer_inst_act_buffer_inst_net4545,
         wrap_act_buffer_inst_act_buffer_inst_net4540,
         wrap_act_buffer_inst_act_buffer_inst_net4535,
         wrap_act_buffer_inst_act_buffer_inst_net4530,
         wrap_act_buffer_inst_act_buffer_inst_net4525,
         wrap_act_buffer_inst_act_buffer_inst_net4519,
         wrap_act_buffer_inst_act_buffer_inst_N162,
         wrap_act_buffer_inst_act_buffer_inst_N161,
         wrap_act_buffer_inst_act_buffer_inst_N160,
         wrap_act_buffer_inst_act_buffer_inst_N159,
         wrap_act_buffer_inst_act_buffer_inst_N158,
         wrap_act_buffer_inst_act_buffer_inst_N157,
         wrap_act_buffer_inst_act_buffer_inst_N156,
         wrap_act_buffer_inst_act_buffer_inst_N155,
         wrap_act_buffer_inst_act_buffer_inst_N154,
         wrap_act_buffer_inst_act_buffer_inst_N153,
         wrap_act_buffer_inst_act_buffer_inst_N152,
         wrap_act_buffer_inst_act_buffer_inst_N151,
         wrap_act_buffer_inst_act_buffer_inst_N150,
         wrap_act_buffer_inst_act_buffer_inst_N149,
         wrap_act_buffer_inst_act_buffer_inst_N148,
         wrap_act_buffer_inst_act_buffer_inst_N147,
         wrap_act_buffer_inst_act_buffer_inst_N146,
         wrap_act_buffer_inst_act_buffer_inst_N145,
         wrap_act_buffer_inst_act_buffer_inst_N144,
         wrap_act_buffer_inst_act_buffer_inst_N143,
         wrap_act_buffer_inst_act_buffer_inst_N142,
         wrap_act_buffer_inst_act_buffer_inst_N141,
         wrap_act_buffer_inst_act_buffer_inst_N140,
         wrap_act_buffer_inst_act_buffer_inst_N139,
         wrap_act_buffer_inst_act_buffer_inst_N138,
         wrap_act_buffer_inst_act_buffer_inst_N137,
         wrap_act_buffer_inst_act_buffer_inst_N136,
         wrap_act_buffer_inst_act_buffer_inst_N135,
         wrap_act_buffer_inst_act_buffer_inst_N134,
         wrap_act_buffer_inst_act_buffer_inst_N133,
         wrap_act_buffer_inst_act_buffer_inst_N132,
         wrap_act_buffer_inst_act_buffer_inst_N131,
         wrap_act_buffer_inst_act_buffer_inst_N130,
         wrap_act_buffer_inst_act_buffer_inst_N129,
         wrap_act_buffer_inst_act_buffer_inst_N128,
         wrap_act_buffer_inst_act_buffer_inst_N127,
         wrap_act_buffer_inst_act_buffer_inst_N126,
         wrap_act_buffer_inst_act_buffer_inst_N125,
         wrap_act_buffer_inst_act_buffer_inst_N124,
         wrap_act_buffer_inst_act_buffer_inst_N123,
         wrap_act_buffer_inst_act_buffer_inst_N122,
         wrap_act_buffer_inst_act_buffer_inst_N121,
         wrap_act_buffer_inst_act_buffer_inst_N120,
         wrap_act_buffer_inst_act_buffer_inst_N119,
         wrap_act_buffer_inst_act_buffer_inst_N118,
         wrap_act_buffer_inst_act_buffer_inst_N117,
         wrap_act_buffer_inst_act_buffer_inst_N116,
         wrap_act_buffer_inst_act_buffer_inst_N115,
         wrap_act_buffer_inst_act_if_inst_n312,
         wrap_act_buffer_inst_act_if_inst_n311,
         wrap_act_buffer_inst_act_if_inst_n310,
         wrap_act_buffer_inst_act_if_inst_n309,
         wrap_act_buffer_inst_act_if_inst_n308,
         wrap_act_buffer_inst_act_if_inst_n307,
         wrap_act_buffer_inst_act_if_inst_n306,
         wrap_act_buffer_inst_act_if_inst_n305,
         wrap_act_buffer_inst_act_if_inst_n304,
         wrap_act_buffer_inst_act_if_inst_n303,
         wrap_act_buffer_inst_act_if_inst_n302,
         wrap_act_buffer_inst_act_if_inst_n301,
         wrap_act_buffer_inst_act_if_inst_n300,
         wrap_act_buffer_inst_act_if_inst_n299,
         wrap_act_buffer_inst_act_if_inst_n298,
         wrap_act_buffer_inst_act_if_inst_n297,
         wrap_act_buffer_inst_act_if_inst_n296,
         wrap_act_buffer_inst_act_if_inst_n295,
         wrap_act_buffer_inst_act_if_inst_n294,
         wrap_act_buffer_inst_act_if_inst_n293,
         wrap_act_buffer_inst_act_if_inst_n292,
         wrap_act_buffer_inst_act_if_inst_n291,
         wrap_act_buffer_inst_act_if_inst_n290,
         wrap_act_buffer_inst_act_if_inst_n289,
         wrap_act_buffer_inst_act_if_inst_n288,
         wrap_act_buffer_inst_act_if_inst_n287,
         wrap_act_buffer_inst_act_if_inst_n286,
         wrap_act_buffer_inst_act_if_inst_n285,
         wrap_act_buffer_inst_act_if_inst_n284,
         wrap_act_buffer_inst_act_if_inst_n283,
         wrap_act_buffer_inst_act_if_inst_n282,
         wrap_act_buffer_inst_act_if_inst_n281,
         wrap_act_buffer_inst_act_if_inst_n280,
         wrap_act_buffer_inst_act_if_inst_n279,
         wrap_act_buffer_inst_act_if_inst_n278,
         wrap_act_buffer_inst_act_if_inst_n277,
         wrap_act_buffer_inst_act_if_inst_n276,
         wrap_act_buffer_inst_act_if_inst_n275,
         wrap_act_buffer_inst_act_if_inst_n274,
         wrap_act_buffer_inst_act_if_inst_n273,
         wrap_act_buffer_inst_act_if_inst_n272,
         wrap_act_buffer_inst_act_if_inst_n271,
         wrap_act_buffer_inst_act_if_inst_n270,
         wrap_act_buffer_inst_act_if_inst_n269,
         wrap_act_buffer_inst_act_if_inst_n268,
         wrap_act_buffer_inst_act_if_inst_n267,
         wrap_act_buffer_inst_act_if_inst_n266,
         wrap_act_buffer_inst_act_if_inst_n265,
         wrap_act_buffer_inst_act_if_inst_n264,
         wrap_act_buffer_inst_act_if_inst_n263,
         wrap_act_buffer_inst_act_if_inst_n262,
         wrap_act_buffer_inst_act_if_inst_n261,
         wrap_act_buffer_inst_act_if_inst_n260,
         wrap_act_buffer_inst_act_if_inst_n259,
         wrap_act_buffer_inst_act_if_inst_n258,
         wrap_act_buffer_inst_act_if_inst_n257,
         wrap_act_buffer_inst_act_if_inst_n256,
         wrap_act_buffer_inst_act_if_inst_n255,
         wrap_act_buffer_inst_act_if_inst_n254,
         wrap_act_buffer_inst_act_if_inst_n253,
         wrap_act_buffer_inst_act_if_inst_n252,
         wrap_act_buffer_inst_act_if_inst_n251,
         wrap_act_buffer_inst_act_if_inst_n250,
         wrap_act_buffer_inst_act_if_inst_n249,
         wrap_act_buffer_inst_act_if_inst_n248,
         wrap_act_buffer_inst_act_if_inst_n247,
         wrap_act_buffer_inst_act_if_inst_n246,
         wrap_act_buffer_inst_act_if_inst_n245,
         wrap_act_buffer_inst_act_if_inst_n244,
         wrap_act_buffer_inst_act_if_inst_n243,
         wrap_act_buffer_inst_act_if_inst_n242,
         wrap_act_buffer_inst_act_if_inst_n241,
         wrap_act_buffer_inst_act_if_inst_n240,
         wrap_act_buffer_inst_act_if_inst_n239,
         wrap_act_buffer_inst_act_if_inst_n238,
         wrap_act_buffer_inst_act_if_inst_n237,
         wrap_act_buffer_inst_act_if_inst_n236,
         wrap_act_buffer_inst_act_if_inst_n235,
         wrap_act_buffer_inst_act_if_inst_n234,
         wrap_act_buffer_inst_act_if_inst_n233,
         wrap_act_buffer_inst_act_if_inst_n232,
         wrap_act_buffer_inst_act_if_inst_n231,
         wrap_act_buffer_inst_act_if_inst_n230,
         wrap_act_buffer_inst_act_if_inst_n229,
         wrap_act_buffer_inst_act_if_inst_n228,
         wrap_act_buffer_inst_act_if_inst_n227,
         wrap_act_buffer_inst_act_if_inst_n226,
         wrap_act_buffer_inst_act_if_inst_n225,
         wrap_act_buffer_inst_act_if_inst_n224,
         wrap_act_buffer_inst_act_if_inst_n223,
         wrap_act_buffer_inst_act_if_inst_n222,
         wrap_act_buffer_inst_act_if_inst_n221,
         wrap_act_buffer_inst_act_if_inst_n220,
         wrap_act_buffer_inst_act_if_inst_n219,
         wrap_act_buffer_inst_act_if_inst_n218,
         wrap_act_buffer_inst_act_if_inst_n217,
         wrap_act_buffer_inst_act_if_inst_n216,
         wrap_act_buffer_inst_act_if_inst_n215,
         wrap_act_buffer_inst_act_if_inst_n214,
         wrap_act_buffer_inst_act_if_inst_n213,
         wrap_act_buffer_inst_act_if_inst_n212,
         wrap_act_buffer_inst_act_if_inst_n211,
         wrap_act_buffer_inst_act_if_inst_n210,
         wrap_act_buffer_inst_act_if_inst_n209,
         wrap_act_buffer_inst_act_if_inst_n208,
         wrap_act_buffer_inst_act_if_inst_n207,
         wrap_act_buffer_inst_act_if_inst_n206,
         wrap_act_buffer_inst_act_if_inst_n205,
         wrap_act_buffer_inst_act_if_inst_n204,
         wrap_act_buffer_inst_act_if_inst_n203,
         wrap_act_buffer_inst_act_if_inst_n202,
         wrap_act_buffer_inst_act_if_inst_n201,
         wrap_act_buffer_inst_act_if_inst_n200,
         wrap_act_buffer_inst_act_if_inst_n199,
         wrap_act_buffer_inst_act_if_inst_n198,
         wrap_act_buffer_inst_act_if_inst_n197,
         wrap_act_buffer_inst_act_if_inst_n196,
         wrap_act_buffer_inst_act_if_inst_n195,
         wrap_act_buffer_inst_act_if_inst_n194,
         wrap_act_buffer_inst_act_if_inst_n193,
         wrap_act_buffer_inst_act_if_inst_n192,
         wrap_act_buffer_inst_act_if_inst_n191,
         wrap_act_buffer_inst_act_if_inst_n190,
         wrap_act_buffer_inst_act_if_inst_n189,
         wrap_act_buffer_inst_act_if_inst_n188,
         wrap_act_buffer_inst_act_if_inst_n187,
         wrap_act_buffer_inst_act_if_inst_n186,
         wrap_act_buffer_inst_act_if_inst_n185,
         wrap_act_buffer_inst_act_if_inst_n184,
         wrap_act_buffer_inst_act_if_inst_n183,
         wrap_act_buffer_inst_act_if_inst_n182,
         wrap_act_buffer_inst_act_if_inst_n181,
         wrap_act_buffer_inst_act_if_inst_n180,
         wrap_act_buffer_inst_act_if_inst_n179,
         wrap_act_buffer_inst_act_if_inst_n178,
         wrap_act_buffer_inst_act_if_inst_n177,
         wrap_act_buffer_inst_act_if_inst_n176,
         wrap_act_buffer_inst_act_if_inst_n175,
         wrap_act_buffer_inst_act_if_inst_n174,
         wrap_act_buffer_inst_act_if_inst_n173,
         wrap_act_buffer_inst_act_if_inst_n172,
         wrap_act_buffer_inst_act_if_inst_n171,
         wrap_act_buffer_inst_act_if_inst_n170,
         wrap_act_buffer_inst_act_if_inst_n169,
         wrap_act_buffer_inst_act_if_inst_n168,
         wrap_act_buffer_inst_act_if_inst_n167,
         wrap_act_buffer_inst_act_if_inst_n166,
         wrap_act_buffer_inst_act_if_inst_n165,
         wrap_act_buffer_inst_act_if_inst_n164,
         wrap_act_buffer_inst_act_if_inst_n163,
         wrap_act_buffer_inst_act_if_inst_n162,
         wrap_act_buffer_inst_act_if_inst_n161,
         wrap_act_buffer_inst_act_if_inst_n160,
         wrap_act_buffer_inst_act_if_inst_n159,
         wrap_act_buffer_inst_act_if_inst_n158,
         wrap_act_buffer_inst_act_if_inst_n157,
         wrap_act_buffer_inst_act_if_inst_n156,
         wrap_act_buffer_inst_act_if_inst_n155,
         wrap_act_buffer_inst_act_if_inst_n154,
         wrap_act_buffer_inst_act_if_inst_n153,
         wrap_act_buffer_inst_act_if_inst_n152,
         wrap_act_buffer_inst_act_if_inst_n151,
         wrap_act_buffer_inst_act_if_inst_n150,
         wrap_act_buffer_inst_act_if_inst_n149,
         wrap_act_buffer_inst_act_if_inst_n148,
         wrap_act_buffer_inst_act_if_inst_n147,
         wrap_act_buffer_inst_act_if_inst_n146,
         wrap_act_buffer_inst_act_if_inst_n145,
         wrap_act_buffer_inst_act_if_inst_n144,
         wrap_act_buffer_inst_act_if_inst_n143,
         wrap_act_buffer_inst_act_if_inst_n142,
         wrap_act_buffer_inst_act_if_inst_n141,
         wrap_act_buffer_inst_act_if_inst_n140,
         wrap_act_buffer_inst_act_if_inst_n139,
         wrap_act_buffer_inst_act_if_inst_n138,
         wrap_act_buffer_inst_act_if_inst_n137,
         wrap_act_buffer_inst_act_if_inst_n136,
         wrap_act_buffer_inst_act_if_inst_n135,
         wrap_act_buffer_inst_act_if_inst_n134,
         wrap_act_buffer_inst_act_if_inst_n133,
         wrap_act_buffer_inst_act_if_inst_n132,
         wrap_act_buffer_inst_act_if_inst_n131,
         wrap_act_buffer_inst_act_if_inst_n130,
         wrap_act_buffer_inst_act_if_inst_n129,
         wrap_act_buffer_inst_act_if_inst_n128,
         wrap_act_buffer_inst_act_if_inst_n127,
         wrap_act_buffer_inst_act_if_inst_n126,
         wrap_act_buffer_inst_act_if_inst_n125,
         wrap_act_buffer_inst_act_if_inst_n124,
         wrap_act_buffer_inst_act_if_inst_n123,
         wrap_act_buffer_inst_act_if_inst_n122,
         wrap_act_buffer_inst_act_if_inst_n121,
         wrap_act_buffer_inst_act_if_inst_n120,
         wrap_act_buffer_inst_act_if_inst_n119,
         wrap_act_buffer_inst_act_if_inst_n118,
         wrap_act_buffer_inst_act_if_inst_n117,
         wrap_act_buffer_inst_act_if_inst_n116,
         wrap_act_buffer_inst_act_if_inst_n115,
         wrap_act_buffer_inst_act_if_inst_n114,
         wrap_act_buffer_inst_act_if_inst_n113,
         wrap_act_buffer_inst_act_if_inst_n112,
         wrap_act_buffer_inst_act_if_inst_n111,
         wrap_act_buffer_inst_act_if_inst_n110,
         wrap_act_buffer_inst_act_if_inst_n109,
         wrap_act_buffer_inst_act_if_inst_n108,
         wrap_act_buffer_inst_act_if_inst_n107,
         wrap_act_buffer_inst_act_if_inst_n106,
         wrap_act_buffer_inst_act_if_inst_n105,
         wrap_act_buffer_inst_act_if_inst_n104,
         wrap_act_buffer_inst_act_if_inst_n103,
         wrap_act_buffer_inst_act_if_inst_n102,
         wrap_act_buffer_inst_act_if_inst_n101,
         wrap_act_buffer_inst_act_if_inst_n100,
         wrap_act_buffer_inst_act_if_inst_n99,
         wrap_act_buffer_inst_act_if_inst_n98,
         wrap_act_buffer_inst_act_if_inst_n97,
         wrap_act_buffer_inst_act_if_inst_n96,
         wrap_act_buffer_inst_act_if_inst_n95,
         wrap_act_buffer_inst_act_if_inst_n94,
         wrap_act_buffer_inst_act_if_inst_n93,
         wrap_act_buffer_inst_act_if_inst_n92,
         wrap_act_buffer_inst_act_if_inst_n91,
         wrap_act_buffer_inst_act_if_inst_n90,
         wrap_act_buffer_inst_act_if_inst_n89,
         wrap_act_buffer_inst_act_if_inst_n88,
         wrap_act_buffer_inst_act_if_inst_n87,
         wrap_act_buffer_inst_act_if_inst_n86,
         wrap_act_buffer_inst_act_if_inst_n85,
         wrap_act_buffer_inst_act_if_inst_n84,
         wrap_act_buffer_inst_act_if_inst_n83,
         wrap_act_buffer_inst_act_if_inst_n82,
         wrap_act_buffer_inst_act_if_inst_n81,
         wrap_act_buffer_inst_act_if_inst_n80,
         wrap_act_buffer_inst_act_if_inst_n79,
         wrap_act_buffer_inst_act_if_inst_n78,
         wrap_act_buffer_inst_act_if_inst_n77,
         wrap_act_buffer_inst_act_if_inst_n76,
         wrap_act_buffer_inst_act_if_inst_n75,
         wrap_act_buffer_inst_act_if_inst_n74,
         wrap_act_buffer_inst_act_if_inst_n73,
         wrap_act_buffer_inst_act_if_inst_n72,
         wrap_act_buffer_inst_act_if_inst_n71,
         wrap_act_buffer_inst_act_if_inst_n70,
         wrap_act_buffer_inst_act_if_inst_n69,
         wrap_act_buffer_inst_act_if_inst_n68,
         wrap_act_buffer_inst_act_if_inst_n67,
         wrap_act_buffer_inst_act_if_inst_n66,
         wrap_act_buffer_inst_act_if_inst_n65,
         wrap_act_buffer_inst_act_if_inst_n64,
         wrap_act_buffer_inst_act_if_inst_n63,
         wrap_act_buffer_inst_act_if_inst_n62,
         wrap_act_buffer_inst_act_if_inst_n61,
         wrap_act_buffer_inst_act_if_inst_n60,
         wrap_act_buffer_inst_act_if_inst_n59,
         wrap_act_buffer_inst_act_if_inst_n58,
         wrap_act_buffer_inst_act_if_inst_n57,
         wrap_act_buffer_inst_act_if_inst_n56,
         wrap_act_buffer_inst_act_if_inst_n55,
         wrap_act_buffer_inst_act_if_inst_n54,
         wrap_act_buffer_inst_act_if_inst_n53,
         wrap_act_buffer_inst_act_if_inst_n52,
         wrap_act_buffer_inst_act_if_inst_n51,
         wrap_act_buffer_inst_act_if_inst_n50,
         wrap_act_buffer_inst_act_if_inst_n49,
         wrap_act_buffer_inst_act_if_inst_n48,
         wrap_act_buffer_inst_act_if_inst_n47,
         wrap_act_buffer_inst_act_if_inst_n46,
         wrap_act_buffer_inst_act_if_inst_n45,
         wrap_act_buffer_inst_act_if_inst_n44,
         wrap_act_buffer_inst_act_if_inst_n43,
         wrap_act_buffer_inst_act_if_inst_n42,
         wrap_act_buffer_inst_act_if_inst_n41,
         wrap_act_buffer_inst_act_if_inst_n40,
         wrap_act_buffer_inst_act_if_inst_n39,
         wrap_act_buffer_inst_act_if_inst_n2,
         wrap_act_buffer_inst_act_if_inst_n1,
         wrap_act_buffer_inst_act_if_inst_n38,
         wrap_act_buffer_inst_act_if_inst_n37,
         wrap_act_buffer_inst_act_if_inst_n36,
         wrap_act_buffer_inst_act_if_inst_n35,
         wrap_act_buffer_inst_act_if_inst_n34,
         wrap_act_buffer_inst_act_if_inst_n33,
         wrap_act_buffer_inst_act_if_inst_n32,
         wrap_act_buffer_inst_act_if_inst_n31,
         wrap_act_buffer_inst_act_if_inst_n30,
         wrap_act_buffer_inst_act_if_inst_n29,
         wrap_act_buffer_inst_act_if_inst_n28,
         wrap_act_buffer_inst_act_if_inst_n27,
         wrap_act_buffer_inst_act_if_inst_n26,
         wrap_act_buffer_inst_act_if_inst_n25,
         wrap_act_buffer_inst_act_if_inst_n24,
         wrap_act_buffer_inst_act_if_inst_n23,
         wrap_act_buffer_inst_act_if_inst_n22,
         wrap_act_buffer_inst_act_if_inst_n21,
         wrap_act_buffer_inst_act_if_inst_n20,
         wrap_act_buffer_inst_act_if_inst_n19,
         wrap_act_buffer_inst_act_if_inst_n18,
         wrap_act_buffer_inst_act_if_inst_n17,
         wrap_act_buffer_inst_act_if_inst_n16,
         wrap_act_buffer_inst_act_if_inst_n15,
         wrap_act_buffer_inst_act_if_inst_n14,
         wrap_act_buffer_inst_act_if_inst_n13,
         wrap_act_buffer_inst_act_if_inst_n12,
         wrap_act_buffer_inst_act_if_inst_n11,
         wrap_act_buffer_inst_act_if_inst_n10,
         wrap_act_buffer_inst_act_if_inst_n9,
         wrap_act_buffer_inst_act_if_inst_n8,
         wrap_act_buffer_inst_act_if_inst_n7,
         wrap_act_buffer_inst_act_if_inst_n6,
         wrap_act_buffer_inst_act_if_inst_n5,
         wrap_act_buffer_inst_act_if_inst_n4,
         wrap_act_buffer_inst_act_if_inst_n3, npu_inst_n125, npu_inst_n124,
         npu_inst_n123, npu_inst_n122, npu_inst_n121, npu_inst_n120,
         npu_inst_n119, npu_inst_n118, npu_inst_n117, npu_inst_n116,
         npu_inst_n115, npu_inst_n114, npu_inst_n113, npu_inst_n112,
         npu_inst_n111, npu_inst_n110, npu_inst_n109, npu_inst_n108,
         npu_inst_n107, npu_inst_n106, npu_inst_n105, npu_inst_n104,
         npu_inst_n103, npu_inst_n102, npu_inst_n101, npu_inst_n100,
         npu_inst_n99, npu_inst_n98, npu_inst_n97, npu_inst_n96, npu_inst_n95,
         npu_inst_n94, npu_inst_n93, npu_inst_n92, npu_inst_n91, npu_inst_n90,
         npu_inst_n89, npu_inst_n88, npu_inst_n87, npu_inst_n86, npu_inst_n85,
         npu_inst_n84, npu_inst_n83, npu_inst_n82, npu_inst_n81, npu_inst_n80,
         npu_inst_n79, npu_inst_n78, npu_inst_n77, npu_inst_n76, npu_inst_n75,
         npu_inst_n74, npu_inst_n73, npu_inst_n72, npu_inst_n71, npu_inst_n70,
         npu_inst_n69, npu_inst_n68, npu_inst_n67, npu_inst_n66, npu_inst_n65,
         npu_inst_n64, npu_inst_n63, npu_inst_n62, npu_inst_n61, npu_inst_n60,
         npu_inst_n59, npu_inst_n58, npu_inst_n57, npu_inst_n56, npu_inst_n55,
         npu_inst_n54, npu_inst_n53, npu_inst_n52, npu_inst_n51, npu_inst_n50,
         npu_inst_n49, npu_inst_n48, npu_inst_n47, npu_inst_n46, npu_inst_n45,
         npu_inst_n44, npu_inst_n43, npu_inst_n42, npu_inst_n41, npu_inst_n40,
         npu_inst_n39, npu_inst_n38, npu_inst_n37, npu_inst_n36, npu_inst_n35,
         npu_inst_n34, npu_inst_n33, npu_inst_n32, npu_inst_n31, npu_inst_n30,
         npu_inst_n29, npu_inst_n28, npu_inst_n27, npu_inst_n26, npu_inst_n25,
         npu_inst_n24, npu_inst_n23, npu_inst_n22, npu_inst_n21, npu_inst_n20,
         npu_inst_n19, npu_inst_n18, npu_inst_n17, npu_inst_n16, npu_inst_n15,
         npu_inst_n14, npu_inst_n13, npu_inst_n12, npu_inst_n11, npu_inst_n10,
         npu_inst_n9, npu_inst_n8, npu_inst_n7, npu_inst_n6, npu_inst_n5,
         npu_inst_n4, npu_inst_n3, npu_inst_n2, npu_inst_n1,
         npu_inst_int_data_res_7__7__0_, npu_inst_int_data_res_7__7__1_,
         npu_inst_int_data_res_7__7__2_, npu_inst_int_data_res_7__7__3_,
         npu_inst_int_data_res_7__7__4_, npu_inst_int_data_res_7__7__5_,
         npu_inst_int_data_res_7__7__6_, npu_inst_int_data_res_7__7__7_,
         npu_inst_int_data_res_7__6__0_, npu_inst_int_data_res_7__6__1_,
         npu_inst_int_data_res_7__6__2_, npu_inst_int_data_res_7__6__3_,
         npu_inst_int_data_res_7__6__4_, npu_inst_int_data_res_7__6__5_,
         npu_inst_int_data_res_7__6__6_, npu_inst_int_data_res_7__6__7_,
         npu_inst_int_data_res_7__5__0_, npu_inst_int_data_res_7__5__1_,
         npu_inst_int_data_res_7__5__2_, npu_inst_int_data_res_7__5__3_,
         npu_inst_int_data_res_7__5__4_, npu_inst_int_data_res_7__5__5_,
         npu_inst_int_data_res_7__5__6_, npu_inst_int_data_res_7__5__7_,
         npu_inst_int_data_res_7__4__0_, npu_inst_int_data_res_7__4__1_,
         npu_inst_int_data_res_7__4__2_, npu_inst_int_data_res_7__4__3_,
         npu_inst_int_data_res_7__4__4_, npu_inst_int_data_res_7__4__5_,
         npu_inst_int_data_res_7__4__6_, npu_inst_int_data_res_7__4__7_,
         npu_inst_int_data_res_7__3__0_, npu_inst_int_data_res_7__3__1_,
         npu_inst_int_data_res_7__3__2_, npu_inst_int_data_res_7__3__3_,
         npu_inst_int_data_res_7__3__4_, npu_inst_int_data_res_7__3__5_,
         npu_inst_int_data_res_7__3__6_, npu_inst_int_data_res_7__3__7_,
         npu_inst_int_data_res_7__2__0_, npu_inst_int_data_res_7__2__1_,
         npu_inst_int_data_res_7__2__2_, npu_inst_int_data_res_7__2__3_,
         npu_inst_int_data_res_7__2__4_, npu_inst_int_data_res_7__2__5_,
         npu_inst_int_data_res_7__2__6_, npu_inst_int_data_res_7__2__7_,
         npu_inst_int_data_res_7__1__0_, npu_inst_int_data_res_7__1__1_,
         npu_inst_int_data_res_7__1__2_, npu_inst_int_data_res_7__1__3_,
         npu_inst_int_data_res_7__1__4_, npu_inst_int_data_res_7__1__5_,
         npu_inst_int_data_res_7__1__6_, npu_inst_int_data_res_7__1__7_,
         npu_inst_int_data_res_7__0__0_, npu_inst_int_data_res_7__0__1_,
         npu_inst_int_data_res_7__0__2_, npu_inst_int_data_res_7__0__3_,
         npu_inst_int_data_res_7__0__4_, npu_inst_int_data_res_7__0__5_,
         npu_inst_int_data_res_7__0__6_, npu_inst_int_data_res_7__0__7_,
         npu_inst_int_data_res_6__7__0_, npu_inst_int_data_res_6__7__1_,
         npu_inst_int_data_res_6__7__2_, npu_inst_int_data_res_6__7__3_,
         npu_inst_int_data_res_6__7__4_, npu_inst_int_data_res_6__7__5_,
         npu_inst_int_data_res_6__7__6_, npu_inst_int_data_res_6__7__7_,
         npu_inst_int_data_res_6__6__0_, npu_inst_int_data_res_6__6__1_,
         npu_inst_int_data_res_6__6__2_, npu_inst_int_data_res_6__6__3_,
         npu_inst_int_data_res_6__6__4_, npu_inst_int_data_res_6__6__5_,
         npu_inst_int_data_res_6__6__6_, npu_inst_int_data_res_6__6__7_,
         npu_inst_int_data_res_6__5__0_, npu_inst_int_data_res_6__5__1_,
         npu_inst_int_data_res_6__5__2_, npu_inst_int_data_res_6__5__3_,
         npu_inst_int_data_res_6__5__4_, npu_inst_int_data_res_6__5__5_,
         npu_inst_int_data_res_6__5__6_, npu_inst_int_data_res_6__5__7_,
         npu_inst_int_data_res_6__4__0_, npu_inst_int_data_res_6__4__1_,
         npu_inst_int_data_res_6__4__2_, npu_inst_int_data_res_6__4__3_,
         npu_inst_int_data_res_6__4__4_, npu_inst_int_data_res_6__4__5_,
         npu_inst_int_data_res_6__4__6_, npu_inst_int_data_res_6__4__7_,
         npu_inst_int_data_res_6__3__0_, npu_inst_int_data_res_6__3__1_,
         npu_inst_int_data_res_6__3__2_, npu_inst_int_data_res_6__3__3_,
         npu_inst_int_data_res_6__3__4_, npu_inst_int_data_res_6__3__5_,
         npu_inst_int_data_res_6__3__6_, npu_inst_int_data_res_6__3__7_,
         npu_inst_int_data_res_6__2__0_, npu_inst_int_data_res_6__2__1_,
         npu_inst_int_data_res_6__2__2_, npu_inst_int_data_res_6__2__3_,
         npu_inst_int_data_res_6__2__4_, npu_inst_int_data_res_6__2__5_,
         npu_inst_int_data_res_6__2__6_, npu_inst_int_data_res_6__2__7_,
         npu_inst_int_data_res_6__1__0_, npu_inst_int_data_res_6__1__1_,
         npu_inst_int_data_res_6__1__2_, npu_inst_int_data_res_6__1__3_,
         npu_inst_int_data_res_6__1__4_, npu_inst_int_data_res_6__1__5_,
         npu_inst_int_data_res_6__1__6_, npu_inst_int_data_res_6__1__7_,
         npu_inst_int_data_res_6__0__0_, npu_inst_int_data_res_6__0__1_,
         npu_inst_int_data_res_6__0__2_, npu_inst_int_data_res_6__0__3_,
         npu_inst_int_data_res_6__0__4_, npu_inst_int_data_res_6__0__5_,
         npu_inst_int_data_res_6__0__6_, npu_inst_int_data_res_6__0__7_,
         npu_inst_int_data_res_5__7__0_, npu_inst_int_data_res_5__7__1_,
         npu_inst_int_data_res_5__7__2_, npu_inst_int_data_res_5__7__3_,
         npu_inst_int_data_res_5__7__4_, npu_inst_int_data_res_5__7__5_,
         npu_inst_int_data_res_5__7__6_, npu_inst_int_data_res_5__7__7_,
         npu_inst_int_data_res_5__6__0_, npu_inst_int_data_res_5__6__1_,
         npu_inst_int_data_res_5__6__2_, npu_inst_int_data_res_5__6__3_,
         npu_inst_int_data_res_5__6__4_, npu_inst_int_data_res_5__6__5_,
         npu_inst_int_data_res_5__6__6_, npu_inst_int_data_res_5__6__7_,
         npu_inst_int_data_res_5__5__0_, npu_inst_int_data_res_5__5__1_,
         npu_inst_int_data_res_5__5__2_, npu_inst_int_data_res_5__5__3_,
         npu_inst_int_data_res_5__5__4_, npu_inst_int_data_res_5__5__5_,
         npu_inst_int_data_res_5__5__6_, npu_inst_int_data_res_5__5__7_,
         npu_inst_int_data_res_5__4__0_, npu_inst_int_data_res_5__4__1_,
         npu_inst_int_data_res_5__4__2_, npu_inst_int_data_res_5__4__3_,
         npu_inst_int_data_res_5__4__4_, npu_inst_int_data_res_5__4__5_,
         npu_inst_int_data_res_5__4__6_, npu_inst_int_data_res_5__4__7_,
         npu_inst_int_data_res_5__3__0_, npu_inst_int_data_res_5__3__1_,
         npu_inst_int_data_res_5__3__2_, npu_inst_int_data_res_5__3__3_,
         npu_inst_int_data_res_5__3__4_, npu_inst_int_data_res_5__3__5_,
         npu_inst_int_data_res_5__3__6_, npu_inst_int_data_res_5__3__7_,
         npu_inst_int_data_res_5__2__0_, npu_inst_int_data_res_5__2__1_,
         npu_inst_int_data_res_5__2__2_, npu_inst_int_data_res_5__2__3_,
         npu_inst_int_data_res_5__2__4_, npu_inst_int_data_res_5__2__5_,
         npu_inst_int_data_res_5__2__6_, npu_inst_int_data_res_5__2__7_,
         npu_inst_int_data_res_5__1__0_, npu_inst_int_data_res_5__1__1_,
         npu_inst_int_data_res_5__1__2_, npu_inst_int_data_res_5__1__3_,
         npu_inst_int_data_res_5__1__4_, npu_inst_int_data_res_5__1__5_,
         npu_inst_int_data_res_5__1__6_, npu_inst_int_data_res_5__1__7_,
         npu_inst_int_data_res_5__0__0_, npu_inst_int_data_res_5__0__1_,
         npu_inst_int_data_res_5__0__2_, npu_inst_int_data_res_5__0__3_,
         npu_inst_int_data_res_5__0__4_, npu_inst_int_data_res_5__0__5_,
         npu_inst_int_data_res_5__0__6_, npu_inst_int_data_res_5__0__7_,
         npu_inst_int_data_res_4__7__0_, npu_inst_int_data_res_4__7__1_,
         npu_inst_int_data_res_4__7__2_, npu_inst_int_data_res_4__7__3_,
         npu_inst_int_data_res_4__7__4_, npu_inst_int_data_res_4__7__5_,
         npu_inst_int_data_res_4__7__6_, npu_inst_int_data_res_4__7__7_,
         npu_inst_int_data_res_4__6__0_, npu_inst_int_data_res_4__6__1_,
         npu_inst_int_data_res_4__6__2_, npu_inst_int_data_res_4__6__3_,
         npu_inst_int_data_res_4__6__4_, npu_inst_int_data_res_4__6__5_,
         npu_inst_int_data_res_4__6__6_, npu_inst_int_data_res_4__6__7_,
         npu_inst_int_data_res_4__5__0_, npu_inst_int_data_res_4__5__1_,
         npu_inst_int_data_res_4__5__2_, npu_inst_int_data_res_4__5__3_,
         npu_inst_int_data_res_4__5__4_, npu_inst_int_data_res_4__5__5_,
         npu_inst_int_data_res_4__5__6_, npu_inst_int_data_res_4__5__7_,
         npu_inst_int_data_res_4__4__0_, npu_inst_int_data_res_4__4__1_,
         npu_inst_int_data_res_4__4__2_, npu_inst_int_data_res_4__4__3_,
         npu_inst_int_data_res_4__4__4_, npu_inst_int_data_res_4__4__5_,
         npu_inst_int_data_res_4__4__6_, npu_inst_int_data_res_4__4__7_,
         npu_inst_int_data_res_4__3__0_, npu_inst_int_data_res_4__3__1_,
         npu_inst_int_data_res_4__3__2_, npu_inst_int_data_res_4__3__3_,
         npu_inst_int_data_res_4__3__4_, npu_inst_int_data_res_4__3__5_,
         npu_inst_int_data_res_4__3__6_, npu_inst_int_data_res_4__3__7_,
         npu_inst_int_data_res_4__2__0_, npu_inst_int_data_res_4__2__1_,
         npu_inst_int_data_res_4__2__2_, npu_inst_int_data_res_4__2__3_,
         npu_inst_int_data_res_4__2__4_, npu_inst_int_data_res_4__2__5_,
         npu_inst_int_data_res_4__2__6_, npu_inst_int_data_res_4__2__7_,
         npu_inst_int_data_res_4__1__0_, npu_inst_int_data_res_4__1__1_,
         npu_inst_int_data_res_4__1__2_, npu_inst_int_data_res_4__1__3_,
         npu_inst_int_data_res_4__1__4_, npu_inst_int_data_res_4__1__5_,
         npu_inst_int_data_res_4__1__6_, npu_inst_int_data_res_4__1__7_,
         npu_inst_int_data_res_4__0__0_, npu_inst_int_data_res_4__0__1_,
         npu_inst_int_data_res_4__0__2_, npu_inst_int_data_res_4__0__3_,
         npu_inst_int_data_res_4__0__4_, npu_inst_int_data_res_4__0__5_,
         npu_inst_int_data_res_4__0__6_, npu_inst_int_data_res_4__0__7_,
         npu_inst_int_data_res_3__7__0_, npu_inst_int_data_res_3__7__1_,
         npu_inst_int_data_res_3__7__2_, npu_inst_int_data_res_3__7__3_,
         npu_inst_int_data_res_3__7__4_, npu_inst_int_data_res_3__7__5_,
         npu_inst_int_data_res_3__7__6_, npu_inst_int_data_res_3__7__7_,
         npu_inst_int_data_res_3__6__0_, npu_inst_int_data_res_3__6__1_,
         npu_inst_int_data_res_3__6__2_, npu_inst_int_data_res_3__6__3_,
         npu_inst_int_data_res_3__6__4_, npu_inst_int_data_res_3__6__5_,
         npu_inst_int_data_res_3__6__6_, npu_inst_int_data_res_3__6__7_,
         npu_inst_int_data_res_3__5__0_, npu_inst_int_data_res_3__5__1_,
         npu_inst_int_data_res_3__5__2_, npu_inst_int_data_res_3__5__3_,
         npu_inst_int_data_res_3__5__4_, npu_inst_int_data_res_3__5__5_,
         npu_inst_int_data_res_3__5__6_, npu_inst_int_data_res_3__5__7_,
         npu_inst_int_data_res_3__4__0_, npu_inst_int_data_res_3__4__1_,
         npu_inst_int_data_res_3__4__2_, npu_inst_int_data_res_3__4__3_,
         npu_inst_int_data_res_3__4__4_, npu_inst_int_data_res_3__4__5_,
         npu_inst_int_data_res_3__4__6_, npu_inst_int_data_res_3__4__7_,
         npu_inst_int_data_res_3__3__0_, npu_inst_int_data_res_3__3__1_,
         npu_inst_int_data_res_3__3__2_, npu_inst_int_data_res_3__3__3_,
         npu_inst_int_data_res_3__3__4_, npu_inst_int_data_res_3__3__5_,
         npu_inst_int_data_res_3__3__6_, npu_inst_int_data_res_3__3__7_,
         npu_inst_int_data_res_3__2__0_, npu_inst_int_data_res_3__2__1_,
         npu_inst_int_data_res_3__2__2_, npu_inst_int_data_res_3__2__3_,
         npu_inst_int_data_res_3__2__4_, npu_inst_int_data_res_3__2__5_,
         npu_inst_int_data_res_3__2__6_, npu_inst_int_data_res_3__2__7_,
         npu_inst_int_data_res_3__1__0_, npu_inst_int_data_res_3__1__1_,
         npu_inst_int_data_res_3__1__2_, npu_inst_int_data_res_3__1__3_,
         npu_inst_int_data_res_3__1__4_, npu_inst_int_data_res_3__1__5_,
         npu_inst_int_data_res_3__1__6_, npu_inst_int_data_res_3__1__7_,
         npu_inst_int_data_res_3__0__0_, npu_inst_int_data_res_3__0__1_,
         npu_inst_int_data_res_3__0__2_, npu_inst_int_data_res_3__0__3_,
         npu_inst_int_data_res_3__0__4_, npu_inst_int_data_res_3__0__5_,
         npu_inst_int_data_res_3__0__6_, npu_inst_int_data_res_3__0__7_,
         npu_inst_int_data_res_2__7__0_, npu_inst_int_data_res_2__7__1_,
         npu_inst_int_data_res_2__7__2_, npu_inst_int_data_res_2__7__3_,
         npu_inst_int_data_res_2__7__4_, npu_inst_int_data_res_2__7__5_,
         npu_inst_int_data_res_2__7__6_, npu_inst_int_data_res_2__7__7_,
         npu_inst_int_data_res_2__6__0_, npu_inst_int_data_res_2__6__1_,
         npu_inst_int_data_res_2__6__2_, npu_inst_int_data_res_2__6__3_,
         npu_inst_int_data_res_2__6__4_, npu_inst_int_data_res_2__6__5_,
         npu_inst_int_data_res_2__6__6_, npu_inst_int_data_res_2__6__7_,
         npu_inst_int_data_res_2__5__0_, npu_inst_int_data_res_2__5__1_,
         npu_inst_int_data_res_2__5__2_, npu_inst_int_data_res_2__5__3_,
         npu_inst_int_data_res_2__5__4_, npu_inst_int_data_res_2__5__5_,
         npu_inst_int_data_res_2__5__6_, npu_inst_int_data_res_2__5__7_,
         npu_inst_int_data_res_2__4__0_, npu_inst_int_data_res_2__4__1_,
         npu_inst_int_data_res_2__4__2_, npu_inst_int_data_res_2__4__3_,
         npu_inst_int_data_res_2__4__4_, npu_inst_int_data_res_2__4__5_,
         npu_inst_int_data_res_2__4__6_, npu_inst_int_data_res_2__4__7_,
         npu_inst_int_data_res_2__3__0_, npu_inst_int_data_res_2__3__1_,
         npu_inst_int_data_res_2__3__2_, npu_inst_int_data_res_2__3__3_,
         npu_inst_int_data_res_2__3__4_, npu_inst_int_data_res_2__3__5_,
         npu_inst_int_data_res_2__3__6_, npu_inst_int_data_res_2__3__7_,
         npu_inst_int_data_res_2__2__0_, npu_inst_int_data_res_2__2__1_,
         npu_inst_int_data_res_2__2__2_, npu_inst_int_data_res_2__2__3_,
         npu_inst_int_data_res_2__2__4_, npu_inst_int_data_res_2__2__5_,
         npu_inst_int_data_res_2__2__6_, npu_inst_int_data_res_2__2__7_,
         npu_inst_int_data_res_2__1__0_, npu_inst_int_data_res_2__1__1_,
         npu_inst_int_data_res_2__1__2_, npu_inst_int_data_res_2__1__3_,
         npu_inst_int_data_res_2__1__4_, npu_inst_int_data_res_2__1__5_,
         npu_inst_int_data_res_2__1__6_, npu_inst_int_data_res_2__1__7_,
         npu_inst_int_data_res_2__0__0_, npu_inst_int_data_res_2__0__1_,
         npu_inst_int_data_res_2__0__2_, npu_inst_int_data_res_2__0__3_,
         npu_inst_int_data_res_2__0__4_, npu_inst_int_data_res_2__0__5_,
         npu_inst_int_data_res_2__0__6_, npu_inst_int_data_res_2__0__7_,
         npu_inst_int_data_res_1__7__0_, npu_inst_int_data_res_1__7__1_,
         npu_inst_int_data_res_1__7__2_, npu_inst_int_data_res_1__7__3_,
         npu_inst_int_data_res_1__7__4_, npu_inst_int_data_res_1__7__5_,
         npu_inst_int_data_res_1__7__6_, npu_inst_int_data_res_1__7__7_,
         npu_inst_int_data_res_1__6__0_, npu_inst_int_data_res_1__6__1_,
         npu_inst_int_data_res_1__6__2_, npu_inst_int_data_res_1__6__3_,
         npu_inst_int_data_res_1__6__4_, npu_inst_int_data_res_1__6__5_,
         npu_inst_int_data_res_1__6__6_, npu_inst_int_data_res_1__6__7_,
         npu_inst_int_data_res_1__5__0_, npu_inst_int_data_res_1__5__1_,
         npu_inst_int_data_res_1__5__2_, npu_inst_int_data_res_1__5__3_,
         npu_inst_int_data_res_1__5__4_, npu_inst_int_data_res_1__5__5_,
         npu_inst_int_data_res_1__5__6_, npu_inst_int_data_res_1__5__7_,
         npu_inst_int_data_res_1__4__0_, npu_inst_int_data_res_1__4__1_,
         npu_inst_int_data_res_1__4__2_, npu_inst_int_data_res_1__4__3_,
         npu_inst_int_data_res_1__4__4_, npu_inst_int_data_res_1__4__5_,
         npu_inst_int_data_res_1__4__6_, npu_inst_int_data_res_1__4__7_,
         npu_inst_int_data_res_1__3__0_, npu_inst_int_data_res_1__3__1_,
         npu_inst_int_data_res_1__3__2_, npu_inst_int_data_res_1__3__3_,
         npu_inst_int_data_res_1__3__4_, npu_inst_int_data_res_1__3__5_,
         npu_inst_int_data_res_1__3__6_, npu_inst_int_data_res_1__3__7_,
         npu_inst_int_data_res_1__2__0_, npu_inst_int_data_res_1__2__1_,
         npu_inst_int_data_res_1__2__2_, npu_inst_int_data_res_1__2__3_,
         npu_inst_int_data_res_1__2__4_, npu_inst_int_data_res_1__2__5_,
         npu_inst_int_data_res_1__2__6_, npu_inst_int_data_res_1__2__7_,
         npu_inst_int_data_res_1__1__0_, npu_inst_int_data_res_1__1__1_,
         npu_inst_int_data_res_1__1__2_, npu_inst_int_data_res_1__1__3_,
         npu_inst_int_data_res_1__1__4_, npu_inst_int_data_res_1__1__5_,
         npu_inst_int_data_res_1__1__6_, npu_inst_int_data_res_1__1__7_,
         npu_inst_int_data_res_1__0__0_, npu_inst_int_data_res_1__0__1_,
         npu_inst_int_data_res_1__0__2_, npu_inst_int_data_res_1__0__3_,
         npu_inst_int_data_res_1__0__4_, npu_inst_int_data_res_1__0__5_,
         npu_inst_int_data_res_1__0__6_, npu_inst_int_data_res_1__0__7_,
         npu_inst_int_data_y_7__7__0_, npu_inst_int_data_y_7__7__1_,
         npu_inst_int_data_y_7__6__0_, npu_inst_int_data_y_7__6__1_,
         npu_inst_int_data_y_7__5__0_, npu_inst_int_data_y_7__5__1_,
         npu_inst_int_data_y_7__4__0_, npu_inst_int_data_y_7__4__1_,
         npu_inst_int_data_y_7__3__0_, npu_inst_int_data_y_7__3__1_,
         npu_inst_int_data_y_7__2__0_, npu_inst_int_data_y_7__2__1_,
         npu_inst_int_data_y_7__1__0_, npu_inst_int_data_y_7__1__1_,
         npu_inst_int_data_y_7__0__0_, npu_inst_int_data_y_7__0__1_,
         npu_inst_int_data_y_6__7__0_, npu_inst_int_data_y_6__7__1_,
         npu_inst_int_data_y_6__6__0_, npu_inst_int_data_y_6__6__1_,
         npu_inst_int_data_y_6__5__0_, npu_inst_int_data_y_6__5__1_,
         npu_inst_int_data_y_6__4__0_, npu_inst_int_data_y_6__4__1_,
         npu_inst_int_data_y_6__3__0_, npu_inst_int_data_y_6__3__1_,
         npu_inst_int_data_y_6__2__0_, npu_inst_int_data_y_6__2__1_,
         npu_inst_int_data_y_6__1__0_, npu_inst_int_data_y_6__1__1_,
         npu_inst_int_data_y_6__0__0_, npu_inst_int_data_y_6__0__1_,
         npu_inst_int_data_y_5__7__0_, npu_inst_int_data_y_5__7__1_,
         npu_inst_int_data_y_5__6__0_, npu_inst_int_data_y_5__6__1_,
         npu_inst_int_data_y_5__5__0_, npu_inst_int_data_y_5__5__1_,
         npu_inst_int_data_y_5__4__0_, npu_inst_int_data_y_5__4__1_,
         npu_inst_int_data_y_5__3__0_, npu_inst_int_data_y_5__3__1_,
         npu_inst_int_data_y_5__2__0_, npu_inst_int_data_y_5__2__1_,
         npu_inst_int_data_y_5__1__0_, npu_inst_int_data_y_5__1__1_,
         npu_inst_int_data_y_5__0__0_, npu_inst_int_data_y_5__0__1_,
         npu_inst_int_data_y_4__7__0_, npu_inst_int_data_y_4__7__1_,
         npu_inst_int_data_y_4__6__0_, npu_inst_int_data_y_4__6__1_,
         npu_inst_int_data_y_4__5__0_, npu_inst_int_data_y_4__5__1_,
         npu_inst_int_data_y_4__4__0_, npu_inst_int_data_y_4__4__1_,
         npu_inst_int_data_y_4__3__0_, npu_inst_int_data_y_4__3__1_,
         npu_inst_int_data_y_4__2__0_, npu_inst_int_data_y_4__2__1_,
         npu_inst_int_data_y_4__1__0_, npu_inst_int_data_y_4__1__1_,
         npu_inst_int_data_y_4__0__0_, npu_inst_int_data_y_4__0__1_,
         npu_inst_int_data_y_3__7__0_, npu_inst_int_data_y_3__7__1_,
         npu_inst_int_data_y_3__6__0_, npu_inst_int_data_y_3__6__1_,
         npu_inst_int_data_y_3__5__0_, npu_inst_int_data_y_3__5__1_,
         npu_inst_int_data_y_3__4__0_, npu_inst_int_data_y_3__4__1_,
         npu_inst_int_data_y_3__3__0_, npu_inst_int_data_y_3__3__1_,
         npu_inst_int_data_y_3__2__0_, npu_inst_int_data_y_3__2__1_,
         npu_inst_int_data_y_3__1__0_, npu_inst_int_data_y_3__1__1_,
         npu_inst_int_data_y_3__0__0_, npu_inst_int_data_y_3__0__1_,
         npu_inst_int_data_y_2__7__0_, npu_inst_int_data_y_2__7__1_,
         npu_inst_int_data_y_2__6__0_, npu_inst_int_data_y_2__6__1_,
         npu_inst_int_data_y_2__5__0_, npu_inst_int_data_y_2__5__1_,
         npu_inst_int_data_y_2__4__0_, npu_inst_int_data_y_2__4__1_,
         npu_inst_int_data_y_2__3__0_, npu_inst_int_data_y_2__3__1_,
         npu_inst_int_data_y_2__2__0_, npu_inst_int_data_y_2__2__1_,
         npu_inst_int_data_y_2__1__0_, npu_inst_int_data_y_2__1__1_,
         npu_inst_int_data_y_2__0__0_, npu_inst_int_data_y_2__0__1_,
         npu_inst_int_data_y_1__7__0_, npu_inst_int_data_y_1__7__1_,
         npu_inst_int_data_y_1__6__0_, npu_inst_int_data_y_1__6__1_,
         npu_inst_int_data_y_1__5__0_, npu_inst_int_data_y_1__5__1_,
         npu_inst_int_data_y_1__4__0_, npu_inst_int_data_y_1__4__1_,
         npu_inst_int_data_y_1__3__0_, npu_inst_int_data_y_1__3__1_,
         npu_inst_int_data_y_1__2__0_, npu_inst_int_data_y_1__2__1_,
         npu_inst_int_data_y_1__1__0_, npu_inst_int_data_y_1__1__1_,
         npu_inst_int_data_y_1__0__0_, npu_inst_int_data_y_1__0__1_,
         npu_inst_int_data_x_7__7__0_, npu_inst_int_data_x_7__7__1_,
         npu_inst_int_data_x_7__6__0_, npu_inst_int_data_x_7__6__1_,
         npu_inst_int_data_x_7__5__0_, npu_inst_int_data_x_7__5__1_,
         npu_inst_int_data_x_7__4__0_, npu_inst_int_data_x_7__4__1_,
         npu_inst_int_data_x_7__3__0_, npu_inst_int_data_x_7__3__1_,
         npu_inst_int_data_x_7__2__0_, npu_inst_int_data_x_7__2__1_,
         npu_inst_int_data_x_7__1__0_, npu_inst_int_data_x_7__1__1_,
         npu_inst_int_data_x_6__7__0_, npu_inst_int_data_x_6__7__1_,
         npu_inst_int_data_x_6__6__0_, npu_inst_int_data_x_6__6__1_,
         npu_inst_int_data_x_6__5__0_, npu_inst_int_data_x_6__5__1_,
         npu_inst_int_data_x_6__4__0_, npu_inst_int_data_x_6__4__1_,
         npu_inst_int_data_x_6__3__0_, npu_inst_int_data_x_6__3__1_,
         npu_inst_int_data_x_6__2__0_, npu_inst_int_data_x_6__2__1_,
         npu_inst_int_data_x_6__1__0_, npu_inst_int_data_x_6__1__1_,
         npu_inst_int_data_x_5__7__0_, npu_inst_int_data_x_5__7__1_,
         npu_inst_int_data_x_5__6__0_, npu_inst_int_data_x_5__6__1_,
         npu_inst_int_data_x_5__5__0_, npu_inst_int_data_x_5__5__1_,
         npu_inst_int_data_x_5__4__0_, npu_inst_int_data_x_5__4__1_,
         npu_inst_int_data_x_5__3__0_, npu_inst_int_data_x_5__3__1_,
         npu_inst_int_data_x_5__2__0_, npu_inst_int_data_x_5__2__1_,
         npu_inst_int_data_x_5__1__0_, npu_inst_int_data_x_5__1__1_,
         npu_inst_int_data_x_4__7__0_, npu_inst_int_data_x_4__7__1_,
         npu_inst_int_data_x_4__6__0_, npu_inst_int_data_x_4__6__1_,
         npu_inst_int_data_x_4__5__0_, npu_inst_int_data_x_4__5__1_,
         npu_inst_int_data_x_4__4__0_, npu_inst_int_data_x_4__4__1_,
         npu_inst_int_data_x_4__3__0_, npu_inst_int_data_x_4__3__1_,
         npu_inst_int_data_x_4__2__0_, npu_inst_int_data_x_4__2__1_,
         npu_inst_int_data_x_4__1__0_, npu_inst_int_data_x_4__1__1_,
         npu_inst_int_data_x_3__7__0_, npu_inst_int_data_x_3__7__1_,
         npu_inst_int_data_x_3__6__0_, npu_inst_int_data_x_3__6__1_,
         npu_inst_int_data_x_3__5__0_, npu_inst_int_data_x_3__5__1_,
         npu_inst_int_data_x_3__4__0_, npu_inst_int_data_x_3__4__1_,
         npu_inst_int_data_x_3__3__0_, npu_inst_int_data_x_3__3__1_,
         npu_inst_int_data_x_3__2__0_, npu_inst_int_data_x_3__2__1_,
         npu_inst_int_data_x_3__1__0_, npu_inst_int_data_x_3__1__1_,
         npu_inst_int_data_x_2__7__0_, npu_inst_int_data_x_2__7__1_,
         npu_inst_int_data_x_2__6__0_, npu_inst_int_data_x_2__6__1_,
         npu_inst_int_data_x_2__5__0_, npu_inst_int_data_x_2__5__1_,
         npu_inst_int_data_x_2__4__0_, npu_inst_int_data_x_2__4__1_,
         npu_inst_int_data_x_2__3__0_, npu_inst_int_data_x_2__3__1_,
         npu_inst_int_data_x_2__2__0_, npu_inst_int_data_x_2__2__1_,
         npu_inst_int_data_x_2__1__0_, npu_inst_int_data_x_2__1__1_,
         npu_inst_int_data_x_1__7__0_, npu_inst_int_data_x_1__7__1_,
         npu_inst_int_data_x_1__6__0_, npu_inst_int_data_x_1__6__1_,
         npu_inst_int_data_x_1__5__0_, npu_inst_int_data_x_1__5__1_,
         npu_inst_int_data_x_1__4__0_, npu_inst_int_data_x_1__4__1_,
         npu_inst_int_data_x_1__3__0_, npu_inst_int_data_x_1__3__1_,
         npu_inst_int_data_x_1__2__0_, npu_inst_int_data_x_1__2__1_,
         npu_inst_int_data_x_1__1__0_, npu_inst_int_data_x_1__1__1_,
         npu_inst_int_data_x_0__7__0_, npu_inst_int_data_x_0__7__1_,
         npu_inst_int_data_x_0__6__0_, npu_inst_int_data_x_0__6__1_,
         npu_inst_int_data_x_0__5__0_, npu_inst_int_data_x_0__5__1_,
         npu_inst_int_data_x_0__4__0_, npu_inst_int_data_x_0__4__1_,
         npu_inst_int_data_x_0__3__0_, npu_inst_int_data_x_0__3__1_,
         npu_inst_int_data_x_0__2__0_, npu_inst_int_data_x_0__2__1_,
         npu_inst_int_data_x_0__1__0_, npu_inst_int_data_x_0__1__1_,
         npu_inst_pe_1_0_0_n116, npu_inst_pe_1_0_0_n115,
         npu_inst_pe_1_0_0_n114, npu_inst_pe_1_0_0_n113,
         npu_inst_pe_1_0_0_n112, npu_inst_pe_1_0_0_n111,
         npu_inst_pe_1_0_0_n110, npu_inst_pe_1_0_0_n109,
         npu_inst_pe_1_0_0_n108, npu_inst_pe_1_0_0_n107,
         npu_inst_pe_1_0_0_n106, npu_inst_pe_1_0_0_n105,
         npu_inst_pe_1_0_0_n104, npu_inst_pe_1_0_0_n103,
         npu_inst_pe_1_0_0_n102, npu_inst_pe_1_0_0_n101,
         npu_inst_pe_1_0_0_n100, npu_inst_pe_1_0_0_n99, npu_inst_pe_1_0_0_n98,
         npu_inst_pe_1_0_0_n36, npu_inst_pe_1_0_0_n35, npu_inst_pe_1_0_0_n34,
         npu_inst_pe_1_0_0_n33, npu_inst_pe_1_0_0_n32, npu_inst_pe_1_0_0_n31,
         npu_inst_pe_1_0_0_n30, npu_inst_pe_1_0_0_n29, npu_inst_pe_1_0_0_n28,
         npu_inst_pe_1_0_0_n25, npu_inst_pe_1_0_0_n24, npu_inst_pe_1_0_0_n23,
         npu_inst_pe_1_0_0_n22, npu_inst_pe_1_0_0_n21, npu_inst_pe_1_0_0_n20,
         npu_inst_pe_1_0_0_n19, npu_inst_pe_1_0_0_n18, npu_inst_pe_1_0_0_n17,
         npu_inst_pe_1_0_0_n16, npu_inst_pe_1_0_0_n15, npu_inst_pe_1_0_0_n14,
         npu_inst_pe_1_0_0_n13, npu_inst_pe_1_0_0_n12, npu_inst_pe_1_0_0_n11,
         npu_inst_pe_1_0_0_n10, npu_inst_pe_1_0_0_n9, npu_inst_pe_1_0_0_n8,
         npu_inst_pe_1_0_0_n7, npu_inst_pe_1_0_0_n6, npu_inst_pe_1_0_0_n5,
         npu_inst_pe_1_0_0_n4, npu_inst_pe_1_0_0_n3, npu_inst_pe_1_0_0_n2,
         npu_inst_pe_1_0_0_n1, npu_inst_pe_1_0_0_sub_77_carry_7_,
         npu_inst_pe_1_0_0_sub_77_carry_6_, npu_inst_pe_1_0_0_sub_77_carry_5_,
         npu_inst_pe_1_0_0_sub_77_carry_4_, npu_inst_pe_1_0_0_sub_77_carry_3_,
         npu_inst_pe_1_0_0_sub_77_carry_2_, npu_inst_pe_1_0_0_sub_77_carry_1_,
         npu_inst_pe_1_0_0_add_79_carry_7_, npu_inst_pe_1_0_0_add_79_carry_6_,
         npu_inst_pe_1_0_0_add_79_carry_5_, npu_inst_pe_1_0_0_add_79_carry_4_,
         npu_inst_pe_1_0_0_add_79_carry_3_, npu_inst_pe_1_0_0_add_79_carry_2_,
         npu_inst_pe_1_0_0_add_79_carry_1_, npu_inst_pe_1_0_0_n97,
         npu_inst_pe_1_0_0_n96, npu_inst_pe_1_0_0_n95, npu_inst_pe_1_0_0_n94,
         npu_inst_pe_1_0_0_n93, npu_inst_pe_1_0_0_n92, npu_inst_pe_1_0_0_n91,
         npu_inst_pe_1_0_0_n90, npu_inst_pe_1_0_0_n89, npu_inst_pe_1_0_0_n88,
         npu_inst_pe_1_0_0_n87, npu_inst_pe_1_0_0_n86, npu_inst_pe_1_0_0_n85,
         npu_inst_pe_1_0_0_n84, npu_inst_pe_1_0_0_n83, npu_inst_pe_1_0_0_n82,
         npu_inst_pe_1_0_0_n81, npu_inst_pe_1_0_0_n80, npu_inst_pe_1_0_0_n79,
         npu_inst_pe_1_0_0_n78, npu_inst_pe_1_0_0_n77, npu_inst_pe_1_0_0_n76,
         npu_inst_pe_1_0_0_n75, npu_inst_pe_1_0_0_n74, npu_inst_pe_1_0_0_n73,
         npu_inst_pe_1_0_0_n72, npu_inst_pe_1_0_0_n71, npu_inst_pe_1_0_0_n70,
         npu_inst_pe_1_0_0_n69, npu_inst_pe_1_0_0_n68, npu_inst_pe_1_0_0_n67,
         npu_inst_pe_1_0_0_n66, npu_inst_pe_1_0_0_n65, npu_inst_pe_1_0_0_n64,
         npu_inst_pe_1_0_0_n63, npu_inst_pe_1_0_0_n62, npu_inst_pe_1_0_0_n61,
         npu_inst_pe_1_0_0_n60, npu_inst_pe_1_0_0_n59, npu_inst_pe_1_0_0_n58,
         npu_inst_pe_1_0_0_n57, npu_inst_pe_1_0_0_n56, npu_inst_pe_1_0_0_n55,
         npu_inst_pe_1_0_0_n54, npu_inst_pe_1_0_0_n53, npu_inst_pe_1_0_0_n52,
         npu_inst_pe_1_0_0_n51, npu_inst_pe_1_0_0_n50, npu_inst_pe_1_0_0_n49,
         npu_inst_pe_1_0_0_n48, npu_inst_pe_1_0_0_n47, npu_inst_pe_1_0_0_n46,
         npu_inst_pe_1_0_0_n45, npu_inst_pe_1_0_0_n44, npu_inst_pe_1_0_0_n43,
         npu_inst_pe_1_0_0_n42, npu_inst_pe_1_0_0_n41, npu_inst_pe_1_0_0_n40,
         npu_inst_pe_1_0_0_n39, npu_inst_pe_1_0_0_n38, npu_inst_pe_1_0_0_n37,
         npu_inst_pe_1_0_0_n27, npu_inst_pe_1_0_0_n26,
         npu_inst_pe_1_0_0_net4484, npu_inst_pe_1_0_0_net4478,
         npu_inst_pe_1_0_0_N94, npu_inst_pe_1_0_0_N93, npu_inst_pe_1_0_0_N84,
         npu_inst_pe_1_0_0_N80, npu_inst_pe_1_0_0_N79, npu_inst_pe_1_0_0_N78,
         npu_inst_pe_1_0_0_N77, npu_inst_pe_1_0_0_N76, npu_inst_pe_1_0_0_N75,
         npu_inst_pe_1_0_0_N74, npu_inst_pe_1_0_0_N73, npu_inst_pe_1_0_0_N72,
         npu_inst_pe_1_0_0_N71, npu_inst_pe_1_0_0_N70, npu_inst_pe_1_0_0_N69,
         npu_inst_pe_1_0_0_N68, npu_inst_pe_1_0_0_N67, npu_inst_pe_1_0_0_N66,
         npu_inst_pe_1_0_0_N65, npu_inst_pe_1_0_0_int_data_0_,
         npu_inst_pe_1_0_0_int_data_1_, npu_inst_pe_1_0_0_int_q_weight_0_,
         npu_inst_pe_1_0_0_int_q_weight_1_,
         npu_inst_pe_1_0_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_0_int_q_reg_h_0__1_, npu_inst_pe_1_0_0_o_data_v_0_,
         npu_inst_pe_1_0_0_o_data_v_1_, npu_inst_pe_1_0_0_o_data_h_0_,
         npu_inst_pe_1_0_0_o_data_h_1_, npu_inst_pe_1_0_1_n116,
         npu_inst_pe_1_0_1_n115, npu_inst_pe_1_0_1_n114,
         npu_inst_pe_1_0_1_n113, npu_inst_pe_1_0_1_n112,
         npu_inst_pe_1_0_1_n111, npu_inst_pe_1_0_1_n110,
         npu_inst_pe_1_0_1_n109, npu_inst_pe_1_0_1_n108,
         npu_inst_pe_1_0_1_n107, npu_inst_pe_1_0_1_n106,
         npu_inst_pe_1_0_1_n105, npu_inst_pe_1_0_1_n104,
         npu_inst_pe_1_0_1_n103, npu_inst_pe_1_0_1_n102,
         npu_inst_pe_1_0_1_n101, npu_inst_pe_1_0_1_n100, npu_inst_pe_1_0_1_n99,
         npu_inst_pe_1_0_1_n98, npu_inst_pe_1_0_1_n36, npu_inst_pe_1_0_1_n35,
         npu_inst_pe_1_0_1_n34, npu_inst_pe_1_0_1_n33, npu_inst_pe_1_0_1_n32,
         npu_inst_pe_1_0_1_n31, npu_inst_pe_1_0_1_n30, npu_inst_pe_1_0_1_n29,
         npu_inst_pe_1_0_1_n28, npu_inst_pe_1_0_1_n25, npu_inst_pe_1_0_1_n24,
         npu_inst_pe_1_0_1_n23, npu_inst_pe_1_0_1_n22, npu_inst_pe_1_0_1_n21,
         npu_inst_pe_1_0_1_n20, npu_inst_pe_1_0_1_n19, npu_inst_pe_1_0_1_n18,
         npu_inst_pe_1_0_1_n17, npu_inst_pe_1_0_1_n16, npu_inst_pe_1_0_1_n15,
         npu_inst_pe_1_0_1_n14, npu_inst_pe_1_0_1_n13, npu_inst_pe_1_0_1_n12,
         npu_inst_pe_1_0_1_n11, npu_inst_pe_1_0_1_n10, npu_inst_pe_1_0_1_n9,
         npu_inst_pe_1_0_1_n8, npu_inst_pe_1_0_1_n7, npu_inst_pe_1_0_1_n6,
         npu_inst_pe_1_0_1_n5, npu_inst_pe_1_0_1_n4, npu_inst_pe_1_0_1_n3,
         npu_inst_pe_1_0_1_n2, npu_inst_pe_1_0_1_n1,
         npu_inst_pe_1_0_1_sub_77_carry_7_, npu_inst_pe_1_0_1_sub_77_carry_6_,
         npu_inst_pe_1_0_1_sub_77_carry_5_, npu_inst_pe_1_0_1_sub_77_carry_4_,
         npu_inst_pe_1_0_1_sub_77_carry_3_, npu_inst_pe_1_0_1_sub_77_carry_2_,
         npu_inst_pe_1_0_1_sub_77_carry_1_, npu_inst_pe_1_0_1_add_79_carry_7_,
         npu_inst_pe_1_0_1_add_79_carry_6_, npu_inst_pe_1_0_1_add_79_carry_5_,
         npu_inst_pe_1_0_1_add_79_carry_4_, npu_inst_pe_1_0_1_add_79_carry_3_,
         npu_inst_pe_1_0_1_add_79_carry_2_, npu_inst_pe_1_0_1_add_79_carry_1_,
         npu_inst_pe_1_0_1_n97, npu_inst_pe_1_0_1_n96, npu_inst_pe_1_0_1_n95,
         npu_inst_pe_1_0_1_n94, npu_inst_pe_1_0_1_n93, npu_inst_pe_1_0_1_n92,
         npu_inst_pe_1_0_1_n91, npu_inst_pe_1_0_1_n90, npu_inst_pe_1_0_1_n89,
         npu_inst_pe_1_0_1_n88, npu_inst_pe_1_0_1_n87, npu_inst_pe_1_0_1_n86,
         npu_inst_pe_1_0_1_n85, npu_inst_pe_1_0_1_n84, npu_inst_pe_1_0_1_n83,
         npu_inst_pe_1_0_1_n82, npu_inst_pe_1_0_1_n81, npu_inst_pe_1_0_1_n80,
         npu_inst_pe_1_0_1_n79, npu_inst_pe_1_0_1_n78, npu_inst_pe_1_0_1_n77,
         npu_inst_pe_1_0_1_n76, npu_inst_pe_1_0_1_n75, npu_inst_pe_1_0_1_n74,
         npu_inst_pe_1_0_1_n73, npu_inst_pe_1_0_1_n72, npu_inst_pe_1_0_1_n71,
         npu_inst_pe_1_0_1_n70, npu_inst_pe_1_0_1_n69, npu_inst_pe_1_0_1_n68,
         npu_inst_pe_1_0_1_n67, npu_inst_pe_1_0_1_n66, npu_inst_pe_1_0_1_n65,
         npu_inst_pe_1_0_1_n64, npu_inst_pe_1_0_1_n63, npu_inst_pe_1_0_1_n62,
         npu_inst_pe_1_0_1_n61, npu_inst_pe_1_0_1_n60, npu_inst_pe_1_0_1_n59,
         npu_inst_pe_1_0_1_n58, npu_inst_pe_1_0_1_n57, npu_inst_pe_1_0_1_n56,
         npu_inst_pe_1_0_1_n55, npu_inst_pe_1_0_1_n54, npu_inst_pe_1_0_1_n53,
         npu_inst_pe_1_0_1_n52, npu_inst_pe_1_0_1_n51, npu_inst_pe_1_0_1_n50,
         npu_inst_pe_1_0_1_n49, npu_inst_pe_1_0_1_n48, npu_inst_pe_1_0_1_n47,
         npu_inst_pe_1_0_1_n46, npu_inst_pe_1_0_1_n45, npu_inst_pe_1_0_1_n44,
         npu_inst_pe_1_0_1_n43, npu_inst_pe_1_0_1_n42, npu_inst_pe_1_0_1_n41,
         npu_inst_pe_1_0_1_n40, npu_inst_pe_1_0_1_n39, npu_inst_pe_1_0_1_n38,
         npu_inst_pe_1_0_1_n37, npu_inst_pe_1_0_1_n27, npu_inst_pe_1_0_1_n26,
         npu_inst_pe_1_0_1_net4461, npu_inst_pe_1_0_1_net4455,
         npu_inst_pe_1_0_1_N94, npu_inst_pe_1_0_1_N93, npu_inst_pe_1_0_1_N84,
         npu_inst_pe_1_0_1_N80, npu_inst_pe_1_0_1_N79, npu_inst_pe_1_0_1_N78,
         npu_inst_pe_1_0_1_N77, npu_inst_pe_1_0_1_N76, npu_inst_pe_1_0_1_N75,
         npu_inst_pe_1_0_1_N74, npu_inst_pe_1_0_1_N73, npu_inst_pe_1_0_1_N72,
         npu_inst_pe_1_0_1_N71, npu_inst_pe_1_0_1_N70, npu_inst_pe_1_0_1_N69,
         npu_inst_pe_1_0_1_N68, npu_inst_pe_1_0_1_N67, npu_inst_pe_1_0_1_N66,
         npu_inst_pe_1_0_1_N65, npu_inst_pe_1_0_1_int_data_0_,
         npu_inst_pe_1_0_1_int_data_1_, npu_inst_pe_1_0_1_int_q_weight_0_,
         npu_inst_pe_1_0_1_int_q_weight_1_,
         npu_inst_pe_1_0_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_1_int_q_reg_h_0__1_, npu_inst_pe_1_0_1_o_data_v_0_,
         npu_inst_pe_1_0_1_o_data_v_1_, npu_inst_pe_1_0_2_n117,
         npu_inst_pe_1_0_2_n116, npu_inst_pe_1_0_2_n115,
         npu_inst_pe_1_0_2_n114, npu_inst_pe_1_0_2_n113,
         npu_inst_pe_1_0_2_n112, npu_inst_pe_1_0_2_n111,
         npu_inst_pe_1_0_2_n110, npu_inst_pe_1_0_2_n109,
         npu_inst_pe_1_0_2_n108, npu_inst_pe_1_0_2_n107,
         npu_inst_pe_1_0_2_n106, npu_inst_pe_1_0_2_n105,
         npu_inst_pe_1_0_2_n104, npu_inst_pe_1_0_2_n103,
         npu_inst_pe_1_0_2_n102, npu_inst_pe_1_0_2_n101,
         npu_inst_pe_1_0_2_n100, npu_inst_pe_1_0_2_n99, npu_inst_pe_1_0_2_n98,
         npu_inst_pe_1_0_2_n36, npu_inst_pe_1_0_2_n35, npu_inst_pe_1_0_2_n34,
         npu_inst_pe_1_0_2_n33, npu_inst_pe_1_0_2_n32, npu_inst_pe_1_0_2_n31,
         npu_inst_pe_1_0_2_n30, npu_inst_pe_1_0_2_n29, npu_inst_pe_1_0_2_n28,
         npu_inst_pe_1_0_2_n25, npu_inst_pe_1_0_2_n24, npu_inst_pe_1_0_2_n23,
         npu_inst_pe_1_0_2_n22, npu_inst_pe_1_0_2_n21, npu_inst_pe_1_0_2_n20,
         npu_inst_pe_1_0_2_n19, npu_inst_pe_1_0_2_n18, npu_inst_pe_1_0_2_n17,
         npu_inst_pe_1_0_2_n16, npu_inst_pe_1_0_2_n15, npu_inst_pe_1_0_2_n14,
         npu_inst_pe_1_0_2_n13, npu_inst_pe_1_0_2_n12, npu_inst_pe_1_0_2_n11,
         npu_inst_pe_1_0_2_n10, npu_inst_pe_1_0_2_n9, npu_inst_pe_1_0_2_n8,
         npu_inst_pe_1_0_2_n7, npu_inst_pe_1_0_2_n6, npu_inst_pe_1_0_2_n5,
         npu_inst_pe_1_0_2_n4, npu_inst_pe_1_0_2_n3, npu_inst_pe_1_0_2_n2,
         npu_inst_pe_1_0_2_n1, npu_inst_pe_1_0_2_sub_77_carry_7_,
         npu_inst_pe_1_0_2_sub_77_carry_6_, npu_inst_pe_1_0_2_sub_77_carry_5_,
         npu_inst_pe_1_0_2_sub_77_carry_4_, npu_inst_pe_1_0_2_sub_77_carry_3_,
         npu_inst_pe_1_0_2_sub_77_carry_2_, npu_inst_pe_1_0_2_sub_77_carry_1_,
         npu_inst_pe_1_0_2_add_79_carry_7_, npu_inst_pe_1_0_2_add_79_carry_6_,
         npu_inst_pe_1_0_2_add_79_carry_5_, npu_inst_pe_1_0_2_add_79_carry_4_,
         npu_inst_pe_1_0_2_add_79_carry_3_, npu_inst_pe_1_0_2_add_79_carry_2_,
         npu_inst_pe_1_0_2_add_79_carry_1_, npu_inst_pe_1_0_2_n97,
         npu_inst_pe_1_0_2_n96, npu_inst_pe_1_0_2_n95, npu_inst_pe_1_0_2_n94,
         npu_inst_pe_1_0_2_n93, npu_inst_pe_1_0_2_n92, npu_inst_pe_1_0_2_n91,
         npu_inst_pe_1_0_2_n90, npu_inst_pe_1_0_2_n89, npu_inst_pe_1_0_2_n88,
         npu_inst_pe_1_0_2_n87, npu_inst_pe_1_0_2_n86, npu_inst_pe_1_0_2_n85,
         npu_inst_pe_1_0_2_n84, npu_inst_pe_1_0_2_n83, npu_inst_pe_1_0_2_n82,
         npu_inst_pe_1_0_2_n81, npu_inst_pe_1_0_2_n80, npu_inst_pe_1_0_2_n79,
         npu_inst_pe_1_0_2_n78, npu_inst_pe_1_0_2_n77, npu_inst_pe_1_0_2_n76,
         npu_inst_pe_1_0_2_n75, npu_inst_pe_1_0_2_n74, npu_inst_pe_1_0_2_n73,
         npu_inst_pe_1_0_2_n72, npu_inst_pe_1_0_2_n71, npu_inst_pe_1_0_2_n70,
         npu_inst_pe_1_0_2_n69, npu_inst_pe_1_0_2_n68, npu_inst_pe_1_0_2_n67,
         npu_inst_pe_1_0_2_n66, npu_inst_pe_1_0_2_n65, npu_inst_pe_1_0_2_n64,
         npu_inst_pe_1_0_2_n63, npu_inst_pe_1_0_2_n62, npu_inst_pe_1_0_2_n61,
         npu_inst_pe_1_0_2_n60, npu_inst_pe_1_0_2_n59, npu_inst_pe_1_0_2_n58,
         npu_inst_pe_1_0_2_n57, npu_inst_pe_1_0_2_n56, npu_inst_pe_1_0_2_n55,
         npu_inst_pe_1_0_2_n54, npu_inst_pe_1_0_2_n53, npu_inst_pe_1_0_2_n52,
         npu_inst_pe_1_0_2_n51, npu_inst_pe_1_0_2_n50, npu_inst_pe_1_0_2_n49,
         npu_inst_pe_1_0_2_n48, npu_inst_pe_1_0_2_n47, npu_inst_pe_1_0_2_n46,
         npu_inst_pe_1_0_2_n45, npu_inst_pe_1_0_2_n44, npu_inst_pe_1_0_2_n43,
         npu_inst_pe_1_0_2_n42, npu_inst_pe_1_0_2_n41, npu_inst_pe_1_0_2_n40,
         npu_inst_pe_1_0_2_n39, npu_inst_pe_1_0_2_n38, npu_inst_pe_1_0_2_n37,
         npu_inst_pe_1_0_2_n27, npu_inst_pe_1_0_2_n26,
         npu_inst_pe_1_0_2_net4438, npu_inst_pe_1_0_2_net4432,
         npu_inst_pe_1_0_2_N94, npu_inst_pe_1_0_2_N93, npu_inst_pe_1_0_2_N84,
         npu_inst_pe_1_0_2_N80, npu_inst_pe_1_0_2_N79, npu_inst_pe_1_0_2_N78,
         npu_inst_pe_1_0_2_N77, npu_inst_pe_1_0_2_N76, npu_inst_pe_1_0_2_N75,
         npu_inst_pe_1_0_2_N74, npu_inst_pe_1_0_2_N73, npu_inst_pe_1_0_2_N72,
         npu_inst_pe_1_0_2_N71, npu_inst_pe_1_0_2_N70, npu_inst_pe_1_0_2_N69,
         npu_inst_pe_1_0_2_N68, npu_inst_pe_1_0_2_N67, npu_inst_pe_1_0_2_N66,
         npu_inst_pe_1_0_2_N65, npu_inst_pe_1_0_2_int_data_0_,
         npu_inst_pe_1_0_2_int_data_1_, npu_inst_pe_1_0_2_int_q_weight_0_,
         npu_inst_pe_1_0_2_int_q_weight_1_,
         npu_inst_pe_1_0_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_2_int_q_reg_h_0__1_, npu_inst_pe_1_0_2_o_data_v_0_,
         npu_inst_pe_1_0_2_o_data_v_1_, npu_inst_pe_1_0_3_n118,
         npu_inst_pe_1_0_3_n117, npu_inst_pe_1_0_3_n116,
         npu_inst_pe_1_0_3_n115, npu_inst_pe_1_0_3_n114,
         npu_inst_pe_1_0_3_n113, npu_inst_pe_1_0_3_n112,
         npu_inst_pe_1_0_3_n111, npu_inst_pe_1_0_3_n110,
         npu_inst_pe_1_0_3_n109, npu_inst_pe_1_0_3_n108,
         npu_inst_pe_1_0_3_n107, npu_inst_pe_1_0_3_n106,
         npu_inst_pe_1_0_3_n105, npu_inst_pe_1_0_3_n104,
         npu_inst_pe_1_0_3_n103, npu_inst_pe_1_0_3_n102,
         npu_inst_pe_1_0_3_n101, npu_inst_pe_1_0_3_n100, npu_inst_pe_1_0_3_n99,
         npu_inst_pe_1_0_3_n98, npu_inst_pe_1_0_3_n36, npu_inst_pe_1_0_3_n35,
         npu_inst_pe_1_0_3_n34, npu_inst_pe_1_0_3_n33, npu_inst_pe_1_0_3_n32,
         npu_inst_pe_1_0_3_n31, npu_inst_pe_1_0_3_n30, npu_inst_pe_1_0_3_n29,
         npu_inst_pe_1_0_3_n28, npu_inst_pe_1_0_3_n25, npu_inst_pe_1_0_3_n24,
         npu_inst_pe_1_0_3_n23, npu_inst_pe_1_0_3_n22, npu_inst_pe_1_0_3_n21,
         npu_inst_pe_1_0_3_n20, npu_inst_pe_1_0_3_n19, npu_inst_pe_1_0_3_n18,
         npu_inst_pe_1_0_3_n17, npu_inst_pe_1_0_3_n16, npu_inst_pe_1_0_3_n15,
         npu_inst_pe_1_0_3_n14, npu_inst_pe_1_0_3_n13, npu_inst_pe_1_0_3_n12,
         npu_inst_pe_1_0_3_n11, npu_inst_pe_1_0_3_n10, npu_inst_pe_1_0_3_n9,
         npu_inst_pe_1_0_3_n8, npu_inst_pe_1_0_3_n7, npu_inst_pe_1_0_3_n6,
         npu_inst_pe_1_0_3_n5, npu_inst_pe_1_0_3_n4, npu_inst_pe_1_0_3_n3,
         npu_inst_pe_1_0_3_n2, npu_inst_pe_1_0_3_n1,
         npu_inst_pe_1_0_3_sub_77_carry_7_, npu_inst_pe_1_0_3_sub_77_carry_6_,
         npu_inst_pe_1_0_3_sub_77_carry_5_, npu_inst_pe_1_0_3_sub_77_carry_4_,
         npu_inst_pe_1_0_3_sub_77_carry_3_, npu_inst_pe_1_0_3_sub_77_carry_2_,
         npu_inst_pe_1_0_3_sub_77_carry_1_, npu_inst_pe_1_0_3_add_79_carry_7_,
         npu_inst_pe_1_0_3_add_79_carry_6_, npu_inst_pe_1_0_3_add_79_carry_5_,
         npu_inst_pe_1_0_3_add_79_carry_4_, npu_inst_pe_1_0_3_add_79_carry_3_,
         npu_inst_pe_1_0_3_add_79_carry_2_, npu_inst_pe_1_0_3_add_79_carry_1_,
         npu_inst_pe_1_0_3_n97, npu_inst_pe_1_0_3_n96, npu_inst_pe_1_0_3_n95,
         npu_inst_pe_1_0_3_n94, npu_inst_pe_1_0_3_n93, npu_inst_pe_1_0_3_n92,
         npu_inst_pe_1_0_3_n91, npu_inst_pe_1_0_3_n90, npu_inst_pe_1_0_3_n89,
         npu_inst_pe_1_0_3_n88, npu_inst_pe_1_0_3_n87, npu_inst_pe_1_0_3_n86,
         npu_inst_pe_1_0_3_n85, npu_inst_pe_1_0_3_n84, npu_inst_pe_1_0_3_n83,
         npu_inst_pe_1_0_3_n82, npu_inst_pe_1_0_3_n81, npu_inst_pe_1_0_3_n80,
         npu_inst_pe_1_0_3_n79, npu_inst_pe_1_0_3_n78, npu_inst_pe_1_0_3_n77,
         npu_inst_pe_1_0_3_n76, npu_inst_pe_1_0_3_n75, npu_inst_pe_1_0_3_n74,
         npu_inst_pe_1_0_3_n73, npu_inst_pe_1_0_3_n72, npu_inst_pe_1_0_3_n71,
         npu_inst_pe_1_0_3_n70, npu_inst_pe_1_0_3_n69, npu_inst_pe_1_0_3_n68,
         npu_inst_pe_1_0_3_n67, npu_inst_pe_1_0_3_n66, npu_inst_pe_1_0_3_n65,
         npu_inst_pe_1_0_3_n64, npu_inst_pe_1_0_3_n63, npu_inst_pe_1_0_3_n62,
         npu_inst_pe_1_0_3_n61, npu_inst_pe_1_0_3_n60, npu_inst_pe_1_0_3_n59,
         npu_inst_pe_1_0_3_n58, npu_inst_pe_1_0_3_n57, npu_inst_pe_1_0_3_n56,
         npu_inst_pe_1_0_3_n55, npu_inst_pe_1_0_3_n54, npu_inst_pe_1_0_3_n53,
         npu_inst_pe_1_0_3_n52, npu_inst_pe_1_0_3_n51, npu_inst_pe_1_0_3_n50,
         npu_inst_pe_1_0_3_n49, npu_inst_pe_1_0_3_n48, npu_inst_pe_1_0_3_n47,
         npu_inst_pe_1_0_3_n46, npu_inst_pe_1_0_3_n45, npu_inst_pe_1_0_3_n44,
         npu_inst_pe_1_0_3_n43, npu_inst_pe_1_0_3_n42, npu_inst_pe_1_0_3_n41,
         npu_inst_pe_1_0_3_n40, npu_inst_pe_1_0_3_n39, npu_inst_pe_1_0_3_n38,
         npu_inst_pe_1_0_3_n37, npu_inst_pe_1_0_3_n27, npu_inst_pe_1_0_3_n26,
         npu_inst_pe_1_0_3_net4415, npu_inst_pe_1_0_3_net4409,
         npu_inst_pe_1_0_3_N94, npu_inst_pe_1_0_3_N93, npu_inst_pe_1_0_3_N84,
         npu_inst_pe_1_0_3_N80, npu_inst_pe_1_0_3_N79, npu_inst_pe_1_0_3_N78,
         npu_inst_pe_1_0_3_N77, npu_inst_pe_1_0_3_N76, npu_inst_pe_1_0_3_N75,
         npu_inst_pe_1_0_3_N74, npu_inst_pe_1_0_3_N73, npu_inst_pe_1_0_3_N72,
         npu_inst_pe_1_0_3_N71, npu_inst_pe_1_0_3_N70, npu_inst_pe_1_0_3_N69,
         npu_inst_pe_1_0_3_N68, npu_inst_pe_1_0_3_N67, npu_inst_pe_1_0_3_N66,
         npu_inst_pe_1_0_3_N65, npu_inst_pe_1_0_3_int_data_0_,
         npu_inst_pe_1_0_3_int_data_1_, npu_inst_pe_1_0_3_int_q_weight_0_,
         npu_inst_pe_1_0_3_int_q_weight_1_,
         npu_inst_pe_1_0_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_3_int_q_reg_h_0__1_, npu_inst_pe_1_0_3_o_data_v_0_,
         npu_inst_pe_1_0_3_o_data_v_1_, npu_inst_pe_1_0_4_n117,
         npu_inst_pe_1_0_4_n116, npu_inst_pe_1_0_4_n115,
         npu_inst_pe_1_0_4_n114, npu_inst_pe_1_0_4_n113,
         npu_inst_pe_1_0_4_n112, npu_inst_pe_1_0_4_n111,
         npu_inst_pe_1_0_4_n110, npu_inst_pe_1_0_4_n109,
         npu_inst_pe_1_0_4_n108, npu_inst_pe_1_0_4_n107,
         npu_inst_pe_1_0_4_n106, npu_inst_pe_1_0_4_n105,
         npu_inst_pe_1_0_4_n104, npu_inst_pe_1_0_4_n103,
         npu_inst_pe_1_0_4_n102, npu_inst_pe_1_0_4_n101,
         npu_inst_pe_1_0_4_n100, npu_inst_pe_1_0_4_n99, npu_inst_pe_1_0_4_n98,
         npu_inst_pe_1_0_4_n36, npu_inst_pe_1_0_4_n35, npu_inst_pe_1_0_4_n34,
         npu_inst_pe_1_0_4_n33, npu_inst_pe_1_0_4_n32, npu_inst_pe_1_0_4_n31,
         npu_inst_pe_1_0_4_n30, npu_inst_pe_1_0_4_n29, npu_inst_pe_1_0_4_n28,
         npu_inst_pe_1_0_4_n25, npu_inst_pe_1_0_4_n24, npu_inst_pe_1_0_4_n23,
         npu_inst_pe_1_0_4_n22, npu_inst_pe_1_0_4_n21, npu_inst_pe_1_0_4_n20,
         npu_inst_pe_1_0_4_n19, npu_inst_pe_1_0_4_n18, npu_inst_pe_1_0_4_n17,
         npu_inst_pe_1_0_4_n16, npu_inst_pe_1_0_4_n15, npu_inst_pe_1_0_4_n14,
         npu_inst_pe_1_0_4_n13, npu_inst_pe_1_0_4_n12, npu_inst_pe_1_0_4_n11,
         npu_inst_pe_1_0_4_n10, npu_inst_pe_1_0_4_n9, npu_inst_pe_1_0_4_n8,
         npu_inst_pe_1_0_4_n7, npu_inst_pe_1_0_4_n6, npu_inst_pe_1_0_4_n5,
         npu_inst_pe_1_0_4_n4, npu_inst_pe_1_0_4_n3, npu_inst_pe_1_0_4_n2,
         npu_inst_pe_1_0_4_n1, npu_inst_pe_1_0_4_sub_77_carry_7_,
         npu_inst_pe_1_0_4_sub_77_carry_6_, npu_inst_pe_1_0_4_sub_77_carry_5_,
         npu_inst_pe_1_0_4_sub_77_carry_4_, npu_inst_pe_1_0_4_sub_77_carry_3_,
         npu_inst_pe_1_0_4_sub_77_carry_2_, npu_inst_pe_1_0_4_sub_77_carry_1_,
         npu_inst_pe_1_0_4_add_79_carry_7_, npu_inst_pe_1_0_4_add_79_carry_6_,
         npu_inst_pe_1_0_4_add_79_carry_5_, npu_inst_pe_1_0_4_add_79_carry_4_,
         npu_inst_pe_1_0_4_add_79_carry_3_, npu_inst_pe_1_0_4_add_79_carry_2_,
         npu_inst_pe_1_0_4_add_79_carry_1_, npu_inst_pe_1_0_4_n97,
         npu_inst_pe_1_0_4_n96, npu_inst_pe_1_0_4_n95, npu_inst_pe_1_0_4_n94,
         npu_inst_pe_1_0_4_n93, npu_inst_pe_1_0_4_n92, npu_inst_pe_1_0_4_n91,
         npu_inst_pe_1_0_4_n90, npu_inst_pe_1_0_4_n89, npu_inst_pe_1_0_4_n88,
         npu_inst_pe_1_0_4_n87, npu_inst_pe_1_0_4_n86, npu_inst_pe_1_0_4_n85,
         npu_inst_pe_1_0_4_n84, npu_inst_pe_1_0_4_n83, npu_inst_pe_1_0_4_n82,
         npu_inst_pe_1_0_4_n81, npu_inst_pe_1_0_4_n80, npu_inst_pe_1_0_4_n79,
         npu_inst_pe_1_0_4_n78, npu_inst_pe_1_0_4_n77, npu_inst_pe_1_0_4_n76,
         npu_inst_pe_1_0_4_n75, npu_inst_pe_1_0_4_n74, npu_inst_pe_1_0_4_n73,
         npu_inst_pe_1_0_4_n72, npu_inst_pe_1_0_4_n71, npu_inst_pe_1_0_4_n70,
         npu_inst_pe_1_0_4_n69, npu_inst_pe_1_0_4_n68, npu_inst_pe_1_0_4_n67,
         npu_inst_pe_1_0_4_n66, npu_inst_pe_1_0_4_n65, npu_inst_pe_1_0_4_n64,
         npu_inst_pe_1_0_4_n63, npu_inst_pe_1_0_4_n62, npu_inst_pe_1_0_4_n61,
         npu_inst_pe_1_0_4_n60, npu_inst_pe_1_0_4_n59, npu_inst_pe_1_0_4_n58,
         npu_inst_pe_1_0_4_n57, npu_inst_pe_1_0_4_n56, npu_inst_pe_1_0_4_n55,
         npu_inst_pe_1_0_4_n54, npu_inst_pe_1_0_4_n53, npu_inst_pe_1_0_4_n52,
         npu_inst_pe_1_0_4_n51, npu_inst_pe_1_0_4_n50, npu_inst_pe_1_0_4_n49,
         npu_inst_pe_1_0_4_n48, npu_inst_pe_1_0_4_n47, npu_inst_pe_1_0_4_n46,
         npu_inst_pe_1_0_4_n45, npu_inst_pe_1_0_4_n44, npu_inst_pe_1_0_4_n43,
         npu_inst_pe_1_0_4_n42, npu_inst_pe_1_0_4_n41, npu_inst_pe_1_0_4_n40,
         npu_inst_pe_1_0_4_n39, npu_inst_pe_1_0_4_n38, npu_inst_pe_1_0_4_n37,
         npu_inst_pe_1_0_4_n27, npu_inst_pe_1_0_4_n26,
         npu_inst_pe_1_0_4_net4392, npu_inst_pe_1_0_4_net4386,
         npu_inst_pe_1_0_4_N94, npu_inst_pe_1_0_4_N93, npu_inst_pe_1_0_4_N84,
         npu_inst_pe_1_0_4_N80, npu_inst_pe_1_0_4_N79, npu_inst_pe_1_0_4_N78,
         npu_inst_pe_1_0_4_N77, npu_inst_pe_1_0_4_N76, npu_inst_pe_1_0_4_N75,
         npu_inst_pe_1_0_4_N74, npu_inst_pe_1_0_4_N73, npu_inst_pe_1_0_4_N72,
         npu_inst_pe_1_0_4_N71, npu_inst_pe_1_0_4_N70, npu_inst_pe_1_0_4_N69,
         npu_inst_pe_1_0_4_N68, npu_inst_pe_1_0_4_N67, npu_inst_pe_1_0_4_N66,
         npu_inst_pe_1_0_4_N65, npu_inst_pe_1_0_4_int_data_0_,
         npu_inst_pe_1_0_4_int_data_1_, npu_inst_pe_1_0_4_int_q_weight_0_,
         npu_inst_pe_1_0_4_int_q_weight_1_,
         npu_inst_pe_1_0_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_4_int_q_reg_h_0__1_, npu_inst_pe_1_0_4_o_data_v_0_,
         npu_inst_pe_1_0_4_o_data_v_1_, npu_inst_pe_1_0_5_n118,
         npu_inst_pe_1_0_5_n117, npu_inst_pe_1_0_5_n116,
         npu_inst_pe_1_0_5_n115, npu_inst_pe_1_0_5_n114,
         npu_inst_pe_1_0_5_n113, npu_inst_pe_1_0_5_n112,
         npu_inst_pe_1_0_5_n111, npu_inst_pe_1_0_5_n110,
         npu_inst_pe_1_0_5_n109, npu_inst_pe_1_0_5_n108,
         npu_inst_pe_1_0_5_n107, npu_inst_pe_1_0_5_n106,
         npu_inst_pe_1_0_5_n105, npu_inst_pe_1_0_5_n104,
         npu_inst_pe_1_0_5_n103, npu_inst_pe_1_0_5_n102,
         npu_inst_pe_1_0_5_n101, npu_inst_pe_1_0_5_n100, npu_inst_pe_1_0_5_n99,
         npu_inst_pe_1_0_5_n98, npu_inst_pe_1_0_5_n36, npu_inst_pe_1_0_5_n35,
         npu_inst_pe_1_0_5_n34, npu_inst_pe_1_0_5_n33, npu_inst_pe_1_0_5_n32,
         npu_inst_pe_1_0_5_n31, npu_inst_pe_1_0_5_n30, npu_inst_pe_1_0_5_n29,
         npu_inst_pe_1_0_5_n28, npu_inst_pe_1_0_5_n25, npu_inst_pe_1_0_5_n24,
         npu_inst_pe_1_0_5_n23, npu_inst_pe_1_0_5_n22, npu_inst_pe_1_0_5_n21,
         npu_inst_pe_1_0_5_n20, npu_inst_pe_1_0_5_n19, npu_inst_pe_1_0_5_n18,
         npu_inst_pe_1_0_5_n17, npu_inst_pe_1_0_5_n16, npu_inst_pe_1_0_5_n15,
         npu_inst_pe_1_0_5_n14, npu_inst_pe_1_0_5_n13, npu_inst_pe_1_0_5_n12,
         npu_inst_pe_1_0_5_n11, npu_inst_pe_1_0_5_n10, npu_inst_pe_1_0_5_n9,
         npu_inst_pe_1_0_5_n8, npu_inst_pe_1_0_5_n7, npu_inst_pe_1_0_5_n6,
         npu_inst_pe_1_0_5_n5, npu_inst_pe_1_0_5_n4, npu_inst_pe_1_0_5_n3,
         npu_inst_pe_1_0_5_n2, npu_inst_pe_1_0_5_n1,
         npu_inst_pe_1_0_5_sub_77_carry_7_, npu_inst_pe_1_0_5_sub_77_carry_6_,
         npu_inst_pe_1_0_5_sub_77_carry_5_, npu_inst_pe_1_0_5_sub_77_carry_4_,
         npu_inst_pe_1_0_5_sub_77_carry_3_, npu_inst_pe_1_0_5_sub_77_carry_2_,
         npu_inst_pe_1_0_5_sub_77_carry_1_, npu_inst_pe_1_0_5_add_79_carry_7_,
         npu_inst_pe_1_0_5_add_79_carry_6_, npu_inst_pe_1_0_5_add_79_carry_5_,
         npu_inst_pe_1_0_5_add_79_carry_4_, npu_inst_pe_1_0_5_add_79_carry_3_,
         npu_inst_pe_1_0_5_add_79_carry_2_, npu_inst_pe_1_0_5_add_79_carry_1_,
         npu_inst_pe_1_0_5_n97, npu_inst_pe_1_0_5_n96, npu_inst_pe_1_0_5_n95,
         npu_inst_pe_1_0_5_n94, npu_inst_pe_1_0_5_n93, npu_inst_pe_1_0_5_n92,
         npu_inst_pe_1_0_5_n91, npu_inst_pe_1_0_5_n90, npu_inst_pe_1_0_5_n89,
         npu_inst_pe_1_0_5_n88, npu_inst_pe_1_0_5_n87, npu_inst_pe_1_0_5_n86,
         npu_inst_pe_1_0_5_n85, npu_inst_pe_1_0_5_n84, npu_inst_pe_1_0_5_n83,
         npu_inst_pe_1_0_5_n82, npu_inst_pe_1_0_5_n81, npu_inst_pe_1_0_5_n80,
         npu_inst_pe_1_0_5_n79, npu_inst_pe_1_0_5_n78, npu_inst_pe_1_0_5_n77,
         npu_inst_pe_1_0_5_n76, npu_inst_pe_1_0_5_n75, npu_inst_pe_1_0_5_n74,
         npu_inst_pe_1_0_5_n73, npu_inst_pe_1_0_5_n72, npu_inst_pe_1_0_5_n71,
         npu_inst_pe_1_0_5_n70, npu_inst_pe_1_0_5_n69, npu_inst_pe_1_0_5_n68,
         npu_inst_pe_1_0_5_n67, npu_inst_pe_1_0_5_n66, npu_inst_pe_1_0_5_n65,
         npu_inst_pe_1_0_5_n64, npu_inst_pe_1_0_5_n63, npu_inst_pe_1_0_5_n62,
         npu_inst_pe_1_0_5_n61, npu_inst_pe_1_0_5_n60, npu_inst_pe_1_0_5_n59,
         npu_inst_pe_1_0_5_n58, npu_inst_pe_1_0_5_n57, npu_inst_pe_1_0_5_n56,
         npu_inst_pe_1_0_5_n55, npu_inst_pe_1_0_5_n54, npu_inst_pe_1_0_5_n53,
         npu_inst_pe_1_0_5_n52, npu_inst_pe_1_0_5_n51, npu_inst_pe_1_0_5_n50,
         npu_inst_pe_1_0_5_n49, npu_inst_pe_1_0_5_n48, npu_inst_pe_1_0_5_n47,
         npu_inst_pe_1_0_5_n46, npu_inst_pe_1_0_5_n45, npu_inst_pe_1_0_5_n44,
         npu_inst_pe_1_0_5_n43, npu_inst_pe_1_0_5_n42, npu_inst_pe_1_0_5_n41,
         npu_inst_pe_1_0_5_n40, npu_inst_pe_1_0_5_n39, npu_inst_pe_1_0_5_n38,
         npu_inst_pe_1_0_5_n37, npu_inst_pe_1_0_5_n27, npu_inst_pe_1_0_5_n26,
         npu_inst_pe_1_0_5_net4369, npu_inst_pe_1_0_5_net4363,
         npu_inst_pe_1_0_5_N94, npu_inst_pe_1_0_5_N93, npu_inst_pe_1_0_5_N84,
         npu_inst_pe_1_0_5_N80, npu_inst_pe_1_0_5_N79, npu_inst_pe_1_0_5_N78,
         npu_inst_pe_1_0_5_N77, npu_inst_pe_1_0_5_N76, npu_inst_pe_1_0_5_N75,
         npu_inst_pe_1_0_5_N74, npu_inst_pe_1_0_5_N73, npu_inst_pe_1_0_5_N72,
         npu_inst_pe_1_0_5_N71, npu_inst_pe_1_0_5_N70, npu_inst_pe_1_0_5_N69,
         npu_inst_pe_1_0_5_N68, npu_inst_pe_1_0_5_N67, npu_inst_pe_1_0_5_N66,
         npu_inst_pe_1_0_5_N65, npu_inst_pe_1_0_5_int_data_0_,
         npu_inst_pe_1_0_5_int_data_1_, npu_inst_pe_1_0_5_int_q_weight_0_,
         npu_inst_pe_1_0_5_int_q_weight_1_,
         npu_inst_pe_1_0_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_5_int_q_reg_h_0__1_, npu_inst_pe_1_0_5_o_data_v_0_,
         npu_inst_pe_1_0_5_o_data_v_1_, npu_inst_pe_1_0_6_n118,
         npu_inst_pe_1_0_6_n117, npu_inst_pe_1_0_6_n116,
         npu_inst_pe_1_0_6_n115, npu_inst_pe_1_0_6_n114,
         npu_inst_pe_1_0_6_n113, npu_inst_pe_1_0_6_n112,
         npu_inst_pe_1_0_6_n111, npu_inst_pe_1_0_6_n110,
         npu_inst_pe_1_0_6_n109, npu_inst_pe_1_0_6_n108,
         npu_inst_pe_1_0_6_n107, npu_inst_pe_1_0_6_n106,
         npu_inst_pe_1_0_6_n105, npu_inst_pe_1_0_6_n104,
         npu_inst_pe_1_0_6_n103, npu_inst_pe_1_0_6_n102,
         npu_inst_pe_1_0_6_n101, npu_inst_pe_1_0_6_n100, npu_inst_pe_1_0_6_n99,
         npu_inst_pe_1_0_6_n98, npu_inst_pe_1_0_6_n36, npu_inst_pe_1_0_6_n35,
         npu_inst_pe_1_0_6_n34, npu_inst_pe_1_0_6_n33, npu_inst_pe_1_0_6_n32,
         npu_inst_pe_1_0_6_n31, npu_inst_pe_1_0_6_n30, npu_inst_pe_1_0_6_n29,
         npu_inst_pe_1_0_6_n28, npu_inst_pe_1_0_6_n25, npu_inst_pe_1_0_6_n24,
         npu_inst_pe_1_0_6_n23, npu_inst_pe_1_0_6_n22, npu_inst_pe_1_0_6_n21,
         npu_inst_pe_1_0_6_n20, npu_inst_pe_1_0_6_n19, npu_inst_pe_1_0_6_n18,
         npu_inst_pe_1_0_6_n17, npu_inst_pe_1_0_6_n16, npu_inst_pe_1_0_6_n15,
         npu_inst_pe_1_0_6_n14, npu_inst_pe_1_0_6_n13, npu_inst_pe_1_0_6_n12,
         npu_inst_pe_1_0_6_n11, npu_inst_pe_1_0_6_n10, npu_inst_pe_1_0_6_n9,
         npu_inst_pe_1_0_6_n8, npu_inst_pe_1_0_6_n7, npu_inst_pe_1_0_6_n6,
         npu_inst_pe_1_0_6_n5, npu_inst_pe_1_0_6_n4, npu_inst_pe_1_0_6_n3,
         npu_inst_pe_1_0_6_n2, npu_inst_pe_1_0_6_n1,
         npu_inst_pe_1_0_6_sub_77_carry_7_, npu_inst_pe_1_0_6_sub_77_carry_6_,
         npu_inst_pe_1_0_6_sub_77_carry_5_, npu_inst_pe_1_0_6_sub_77_carry_4_,
         npu_inst_pe_1_0_6_sub_77_carry_3_, npu_inst_pe_1_0_6_sub_77_carry_2_,
         npu_inst_pe_1_0_6_sub_77_carry_1_, npu_inst_pe_1_0_6_add_79_carry_7_,
         npu_inst_pe_1_0_6_add_79_carry_6_, npu_inst_pe_1_0_6_add_79_carry_5_,
         npu_inst_pe_1_0_6_add_79_carry_4_, npu_inst_pe_1_0_6_add_79_carry_3_,
         npu_inst_pe_1_0_6_add_79_carry_2_, npu_inst_pe_1_0_6_add_79_carry_1_,
         npu_inst_pe_1_0_6_n97, npu_inst_pe_1_0_6_n96, npu_inst_pe_1_0_6_n95,
         npu_inst_pe_1_0_6_n94, npu_inst_pe_1_0_6_n93, npu_inst_pe_1_0_6_n92,
         npu_inst_pe_1_0_6_n91, npu_inst_pe_1_0_6_n90, npu_inst_pe_1_0_6_n89,
         npu_inst_pe_1_0_6_n88, npu_inst_pe_1_0_6_n87, npu_inst_pe_1_0_6_n86,
         npu_inst_pe_1_0_6_n85, npu_inst_pe_1_0_6_n84, npu_inst_pe_1_0_6_n83,
         npu_inst_pe_1_0_6_n82, npu_inst_pe_1_0_6_n81, npu_inst_pe_1_0_6_n80,
         npu_inst_pe_1_0_6_n79, npu_inst_pe_1_0_6_n78, npu_inst_pe_1_0_6_n77,
         npu_inst_pe_1_0_6_n76, npu_inst_pe_1_0_6_n75, npu_inst_pe_1_0_6_n74,
         npu_inst_pe_1_0_6_n73, npu_inst_pe_1_0_6_n72, npu_inst_pe_1_0_6_n71,
         npu_inst_pe_1_0_6_n70, npu_inst_pe_1_0_6_n69, npu_inst_pe_1_0_6_n68,
         npu_inst_pe_1_0_6_n67, npu_inst_pe_1_0_6_n66, npu_inst_pe_1_0_6_n65,
         npu_inst_pe_1_0_6_n64, npu_inst_pe_1_0_6_n63, npu_inst_pe_1_0_6_n62,
         npu_inst_pe_1_0_6_n61, npu_inst_pe_1_0_6_n60, npu_inst_pe_1_0_6_n59,
         npu_inst_pe_1_0_6_n58, npu_inst_pe_1_0_6_n57, npu_inst_pe_1_0_6_n56,
         npu_inst_pe_1_0_6_n55, npu_inst_pe_1_0_6_n54, npu_inst_pe_1_0_6_n53,
         npu_inst_pe_1_0_6_n52, npu_inst_pe_1_0_6_n51, npu_inst_pe_1_0_6_n50,
         npu_inst_pe_1_0_6_n49, npu_inst_pe_1_0_6_n48, npu_inst_pe_1_0_6_n47,
         npu_inst_pe_1_0_6_n46, npu_inst_pe_1_0_6_n45, npu_inst_pe_1_0_6_n44,
         npu_inst_pe_1_0_6_n43, npu_inst_pe_1_0_6_n42, npu_inst_pe_1_0_6_n41,
         npu_inst_pe_1_0_6_n40, npu_inst_pe_1_0_6_n39, npu_inst_pe_1_0_6_n38,
         npu_inst_pe_1_0_6_n37, npu_inst_pe_1_0_6_n27, npu_inst_pe_1_0_6_n26,
         npu_inst_pe_1_0_6_net4346, npu_inst_pe_1_0_6_net4340,
         npu_inst_pe_1_0_6_N94, npu_inst_pe_1_0_6_N93, npu_inst_pe_1_0_6_N84,
         npu_inst_pe_1_0_6_N80, npu_inst_pe_1_0_6_N79, npu_inst_pe_1_0_6_N78,
         npu_inst_pe_1_0_6_N77, npu_inst_pe_1_0_6_N76, npu_inst_pe_1_0_6_N75,
         npu_inst_pe_1_0_6_N74, npu_inst_pe_1_0_6_N73, npu_inst_pe_1_0_6_N72,
         npu_inst_pe_1_0_6_N71, npu_inst_pe_1_0_6_N70, npu_inst_pe_1_0_6_N69,
         npu_inst_pe_1_0_6_N68, npu_inst_pe_1_0_6_N67, npu_inst_pe_1_0_6_N66,
         npu_inst_pe_1_0_6_N65, npu_inst_pe_1_0_6_int_data_0_,
         npu_inst_pe_1_0_6_int_data_1_, npu_inst_pe_1_0_6_int_q_weight_0_,
         npu_inst_pe_1_0_6_int_q_weight_1_,
         npu_inst_pe_1_0_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_6_int_q_reg_h_0__1_, npu_inst_pe_1_0_6_o_data_v_0_,
         npu_inst_pe_1_0_6_o_data_v_1_, npu_inst_pe_1_0_7_n118,
         npu_inst_pe_1_0_7_n117, npu_inst_pe_1_0_7_n116,
         npu_inst_pe_1_0_7_n115, npu_inst_pe_1_0_7_n114,
         npu_inst_pe_1_0_7_n113, npu_inst_pe_1_0_7_n112,
         npu_inst_pe_1_0_7_n111, npu_inst_pe_1_0_7_n110,
         npu_inst_pe_1_0_7_n109, npu_inst_pe_1_0_7_n108,
         npu_inst_pe_1_0_7_n107, npu_inst_pe_1_0_7_n106,
         npu_inst_pe_1_0_7_n105, npu_inst_pe_1_0_7_n104,
         npu_inst_pe_1_0_7_n103, npu_inst_pe_1_0_7_n102,
         npu_inst_pe_1_0_7_n101, npu_inst_pe_1_0_7_n100, npu_inst_pe_1_0_7_n99,
         npu_inst_pe_1_0_7_n98, npu_inst_pe_1_0_7_n36, npu_inst_pe_1_0_7_n35,
         npu_inst_pe_1_0_7_n34, npu_inst_pe_1_0_7_n33, npu_inst_pe_1_0_7_n32,
         npu_inst_pe_1_0_7_n31, npu_inst_pe_1_0_7_n30, npu_inst_pe_1_0_7_n29,
         npu_inst_pe_1_0_7_n28, npu_inst_pe_1_0_7_n25, npu_inst_pe_1_0_7_n24,
         npu_inst_pe_1_0_7_n23, npu_inst_pe_1_0_7_n22, npu_inst_pe_1_0_7_n21,
         npu_inst_pe_1_0_7_n20, npu_inst_pe_1_0_7_n19, npu_inst_pe_1_0_7_n18,
         npu_inst_pe_1_0_7_n17, npu_inst_pe_1_0_7_n16, npu_inst_pe_1_0_7_n15,
         npu_inst_pe_1_0_7_n14, npu_inst_pe_1_0_7_n13, npu_inst_pe_1_0_7_n12,
         npu_inst_pe_1_0_7_n11, npu_inst_pe_1_0_7_n10, npu_inst_pe_1_0_7_n9,
         npu_inst_pe_1_0_7_n8, npu_inst_pe_1_0_7_n7, npu_inst_pe_1_0_7_n6,
         npu_inst_pe_1_0_7_n5, npu_inst_pe_1_0_7_n4, npu_inst_pe_1_0_7_n3,
         npu_inst_pe_1_0_7_n2, npu_inst_pe_1_0_7_n1,
         npu_inst_pe_1_0_7_sub_77_carry_7_, npu_inst_pe_1_0_7_sub_77_carry_6_,
         npu_inst_pe_1_0_7_sub_77_carry_5_, npu_inst_pe_1_0_7_sub_77_carry_4_,
         npu_inst_pe_1_0_7_sub_77_carry_3_, npu_inst_pe_1_0_7_sub_77_carry_2_,
         npu_inst_pe_1_0_7_sub_77_carry_1_, npu_inst_pe_1_0_7_add_79_carry_7_,
         npu_inst_pe_1_0_7_add_79_carry_6_, npu_inst_pe_1_0_7_add_79_carry_5_,
         npu_inst_pe_1_0_7_add_79_carry_4_, npu_inst_pe_1_0_7_add_79_carry_3_,
         npu_inst_pe_1_0_7_add_79_carry_2_, npu_inst_pe_1_0_7_add_79_carry_1_,
         npu_inst_pe_1_0_7_n97, npu_inst_pe_1_0_7_n96, npu_inst_pe_1_0_7_n95,
         npu_inst_pe_1_0_7_n94, npu_inst_pe_1_0_7_n93, npu_inst_pe_1_0_7_n92,
         npu_inst_pe_1_0_7_n91, npu_inst_pe_1_0_7_n90, npu_inst_pe_1_0_7_n89,
         npu_inst_pe_1_0_7_n88, npu_inst_pe_1_0_7_n87, npu_inst_pe_1_0_7_n86,
         npu_inst_pe_1_0_7_n85, npu_inst_pe_1_0_7_n84, npu_inst_pe_1_0_7_n83,
         npu_inst_pe_1_0_7_n82, npu_inst_pe_1_0_7_n81, npu_inst_pe_1_0_7_n80,
         npu_inst_pe_1_0_7_n79, npu_inst_pe_1_0_7_n78, npu_inst_pe_1_0_7_n77,
         npu_inst_pe_1_0_7_n76, npu_inst_pe_1_0_7_n75, npu_inst_pe_1_0_7_n74,
         npu_inst_pe_1_0_7_n73, npu_inst_pe_1_0_7_n72, npu_inst_pe_1_0_7_n71,
         npu_inst_pe_1_0_7_n70, npu_inst_pe_1_0_7_n69, npu_inst_pe_1_0_7_n68,
         npu_inst_pe_1_0_7_n67, npu_inst_pe_1_0_7_n66, npu_inst_pe_1_0_7_n65,
         npu_inst_pe_1_0_7_n64, npu_inst_pe_1_0_7_n63, npu_inst_pe_1_0_7_n62,
         npu_inst_pe_1_0_7_n61, npu_inst_pe_1_0_7_n60, npu_inst_pe_1_0_7_n59,
         npu_inst_pe_1_0_7_n58, npu_inst_pe_1_0_7_n57, npu_inst_pe_1_0_7_n56,
         npu_inst_pe_1_0_7_n55, npu_inst_pe_1_0_7_n54, npu_inst_pe_1_0_7_n53,
         npu_inst_pe_1_0_7_n52, npu_inst_pe_1_0_7_n51, npu_inst_pe_1_0_7_n50,
         npu_inst_pe_1_0_7_n49, npu_inst_pe_1_0_7_n48, npu_inst_pe_1_0_7_n47,
         npu_inst_pe_1_0_7_n46, npu_inst_pe_1_0_7_n45, npu_inst_pe_1_0_7_n44,
         npu_inst_pe_1_0_7_n43, npu_inst_pe_1_0_7_n42, npu_inst_pe_1_0_7_n41,
         npu_inst_pe_1_0_7_n40, npu_inst_pe_1_0_7_n39, npu_inst_pe_1_0_7_n38,
         npu_inst_pe_1_0_7_n37, npu_inst_pe_1_0_7_n27, npu_inst_pe_1_0_7_n26,
         npu_inst_pe_1_0_7_net4323, npu_inst_pe_1_0_7_net4317,
         npu_inst_pe_1_0_7_N94, npu_inst_pe_1_0_7_N93, npu_inst_pe_1_0_7_N84,
         npu_inst_pe_1_0_7_N80, npu_inst_pe_1_0_7_N79, npu_inst_pe_1_0_7_N78,
         npu_inst_pe_1_0_7_N77, npu_inst_pe_1_0_7_N76, npu_inst_pe_1_0_7_N75,
         npu_inst_pe_1_0_7_N74, npu_inst_pe_1_0_7_N73, npu_inst_pe_1_0_7_N72,
         npu_inst_pe_1_0_7_N71, npu_inst_pe_1_0_7_N70, npu_inst_pe_1_0_7_N69,
         npu_inst_pe_1_0_7_N68, npu_inst_pe_1_0_7_N67, npu_inst_pe_1_0_7_N66,
         npu_inst_pe_1_0_7_N65, npu_inst_pe_1_0_7_int_data_0_,
         npu_inst_pe_1_0_7_int_data_1_, npu_inst_pe_1_0_7_int_q_weight_0_,
         npu_inst_pe_1_0_7_int_q_weight_1_,
         npu_inst_pe_1_0_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_0_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_0_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_0_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_0_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_0_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_0_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_0_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_0_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_0_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_0_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_0_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_0_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_0_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_0_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_0_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_0_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_0_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_0_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_0_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_0_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_0_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_0_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_0_7_int_q_reg_h_0__1_, npu_inst_pe_1_0_7_o_data_v_0_,
         npu_inst_pe_1_0_7_o_data_v_1_, npu_inst_pe_1_1_0_n118,
         npu_inst_pe_1_1_0_n117, npu_inst_pe_1_1_0_n116,
         npu_inst_pe_1_1_0_n115, npu_inst_pe_1_1_0_n114,
         npu_inst_pe_1_1_0_n113, npu_inst_pe_1_1_0_n112,
         npu_inst_pe_1_1_0_n111, npu_inst_pe_1_1_0_n110,
         npu_inst_pe_1_1_0_n109, npu_inst_pe_1_1_0_n108,
         npu_inst_pe_1_1_0_n107, npu_inst_pe_1_1_0_n106,
         npu_inst_pe_1_1_0_n105, npu_inst_pe_1_1_0_n104,
         npu_inst_pe_1_1_0_n103, npu_inst_pe_1_1_0_n102,
         npu_inst_pe_1_1_0_n101, npu_inst_pe_1_1_0_n100, npu_inst_pe_1_1_0_n99,
         npu_inst_pe_1_1_0_n98, npu_inst_pe_1_1_0_n36, npu_inst_pe_1_1_0_n35,
         npu_inst_pe_1_1_0_n34, npu_inst_pe_1_1_0_n33, npu_inst_pe_1_1_0_n32,
         npu_inst_pe_1_1_0_n31, npu_inst_pe_1_1_0_n30, npu_inst_pe_1_1_0_n29,
         npu_inst_pe_1_1_0_n28, npu_inst_pe_1_1_0_n25, npu_inst_pe_1_1_0_n24,
         npu_inst_pe_1_1_0_n23, npu_inst_pe_1_1_0_n22, npu_inst_pe_1_1_0_n21,
         npu_inst_pe_1_1_0_n20, npu_inst_pe_1_1_0_n19, npu_inst_pe_1_1_0_n18,
         npu_inst_pe_1_1_0_n17, npu_inst_pe_1_1_0_n16, npu_inst_pe_1_1_0_n15,
         npu_inst_pe_1_1_0_n14, npu_inst_pe_1_1_0_n13, npu_inst_pe_1_1_0_n12,
         npu_inst_pe_1_1_0_n11, npu_inst_pe_1_1_0_n10, npu_inst_pe_1_1_0_n9,
         npu_inst_pe_1_1_0_n8, npu_inst_pe_1_1_0_n7, npu_inst_pe_1_1_0_n6,
         npu_inst_pe_1_1_0_n5, npu_inst_pe_1_1_0_n4, npu_inst_pe_1_1_0_n3,
         npu_inst_pe_1_1_0_n2, npu_inst_pe_1_1_0_n1,
         npu_inst_pe_1_1_0_sub_77_carry_7_, npu_inst_pe_1_1_0_sub_77_carry_6_,
         npu_inst_pe_1_1_0_sub_77_carry_5_, npu_inst_pe_1_1_0_sub_77_carry_4_,
         npu_inst_pe_1_1_0_sub_77_carry_3_, npu_inst_pe_1_1_0_sub_77_carry_2_,
         npu_inst_pe_1_1_0_sub_77_carry_1_, npu_inst_pe_1_1_0_add_79_carry_7_,
         npu_inst_pe_1_1_0_add_79_carry_6_, npu_inst_pe_1_1_0_add_79_carry_5_,
         npu_inst_pe_1_1_0_add_79_carry_4_, npu_inst_pe_1_1_0_add_79_carry_3_,
         npu_inst_pe_1_1_0_add_79_carry_2_, npu_inst_pe_1_1_0_add_79_carry_1_,
         npu_inst_pe_1_1_0_n97, npu_inst_pe_1_1_0_n96, npu_inst_pe_1_1_0_n95,
         npu_inst_pe_1_1_0_n94, npu_inst_pe_1_1_0_n93, npu_inst_pe_1_1_0_n92,
         npu_inst_pe_1_1_0_n91, npu_inst_pe_1_1_0_n90, npu_inst_pe_1_1_0_n89,
         npu_inst_pe_1_1_0_n88, npu_inst_pe_1_1_0_n87, npu_inst_pe_1_1_0_n86,
         npu_inst_pe_1_1_0_n85, npu_inst_pe_1_1_0_n84, npu_inst_pe_1_1_0_n83,
         npu_inst_pe_1_1_0_n82, npu_inst_pe_1_1_0_n81, npu_inst_pe_1_1_0_n80,
         npu_inst_pe_1_1_0_n79, npu_inst_pe_1_1_0_n78, npu_inst_pe_1_1_0_n77,
         npu_inst_pe_1_1_0_n76, npu_inst_pe_1_1_0_n75, npu_inst_pe_1_1_0_n74,
         npu_inst_pe_1_1_0_n73, npu_inst_pe_1_1_0_n72, npu_inst_pe_1_1_0_n71,
         npu_inst_pe_1_1_0_n70, npu_inst_pe_1_1_0_n69, npu_inst_pe_1_1_0_n68,
         npu_inst_pe_1_1_0_n67, npu_inst_pe_1_1_0_n66, npu_inst_pe_1_1_0_n65,
         npu_inst_pe_1_1_0_n64, npu_inst_pe_1_1_0_n63, npu_inst_pe_1_1_0_n62,
         npu_inst_pe_1_1_0_n61, npu_inst_pe_1_1_0_n60, npu_inst_pe_1_1_0_n59,
         npu_inst_pe_1_1_0_n58, npu_inst_pe_1_1_0_n57, npu_inst_pe_1_1_0_n56,
         npu_inst_pe_1_1_0_n55, npu_inst_pe_1_1_0_n54, npu_inst_pe_1_1_0_n53,
         npu_inst_pe_1_1_0_n52, npu_inst_pe_1_1_0_n51, npu_inst_pe_1_1_0_n50,
         npu_inst_pe_1_1_0_n49, npu_inst_pe_1_1_0_n48, npu_inst_pe_1_1_0_n47,
         npu_inst_pe_1_1_0_n46, npu_inst_pe_1_1_0_n45, npu_inst_pe_1_1_0_n44,
         npu_inst_pe_1_1_0_n43, npu_inst_pe_1_1_0_n42, npu_inst_pe_1_1_0_n41,
         npu_inst_pe_1_1_0_n40, npu_inst_pe_1_1_0_n39, npu_inst_pe_1_1_0_n38,
         npu_inst_pe_1_1_0_n37, npu_inst_pe_1_1_0_n27, npu_inst_pe_1_1_0_n26,
         npu_inst_pe_1_1_0_net4300, npu_inst_pe_1_1_0_net4294,
         npu_inst_pe_1_1_0_N94, npu_inst_pe_1_1_0_N93, npu_inst_pe_1_1_0_N84,
         npu_inst_pe_1_1_0_N80, npu_inst_pe_1_1_0_N79, npu_inst_pe_1_1_0_N78,
         npu_inst_pe_1_1_0_N77, npu_inst_pe_1_1_0_N76, npu_inst_pe_1_1_0_N75,
         npu_inst_pe_1_1_0_N74, npu_inst_pe_1_1_0_N73, npu_inst_pe_1_1_0_N72,
         npu_inst_pe_1_1_0_N71, npu_inst_pe_1_1_0_N70, npu_inst_pe_1_1_0_N69,
         npu_inst_pe_1_1_0_N68, npu_inst_pe_1_1_0_N67, npu_inst_pe_1_1_0_N66,
         npu_inst_pe_1_1_0_N65, npu_inst_pe_1_1_0_int_data_0_,
         npu_inst_pe_1_1_0_int_data_1_, npu_inst_pe_1_1_0_int_q_weight_0_,
         npu_inst_pe_1_1_0_int_q_weight_1_,
         npu_inst_pe_1_1_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_0_int_q_reg_h_0__1_, npu_inst_pe_1_1_0_o_data_h_0_,
         npu_inst_pe_1_1_0_o_data_h_1_, npu_inst_pe_1_1_1_n118,
         npu_inst_pe_1_1_1_n117, npu_inst_pe_1_1_1_n116,
         npu_inst_pe_1_1_1_n115, npu_inst_pe_1_1_1_n114,
         npu_inst_pe_1_1_1_n113, npu_inst_pe_1_1_1_n112,
         npu_inst_pe_1_1_1_n111, npu_inst_pe_1_1_1_n110,
         npu_inst_pe_1_1_1_n109, npu_inst_pe_1_1_1_n108,
         npu_inst_pe_1_1_1_n107, npu_inst_pe_1_1_1_n106,
         npu_inst_pe_1_1_1_n105, npu_inst_pe_1_1_1_n104,
         npu_inst_pe_1_1_1_n103, npu_inst_pe_1_1_1_n102,
         npu_inst_pe_1_1_1_n101, npu_inst_pe_1_1_1_n100, npu_inst_pe_1_1_1_n99,
         npu_inst_pe_1_1_1_n98, npu_inst_pe_1_1_1_n36, npu_inst_pe_1_1_1_n35,
         npu_inst_pe_1_1_1_n34, npu_inst_pe_1_1_1_n33, npu_inst_pe_1_1_1_n32,
         npu_inst_pe_1_1_1_n31, npu_inst_pe_1_1_1_n30, npu_inst_pe_1_1_1_n29,
         npu_inst_pe_1_1_1_n28, npu_inst_pe_1_1_1_n25, npu_inst_pe_1_1_1_n24,
         npu_inst_pe_1_1_1_n23, npu_inst_pe_1_1_1_n22, npu_inst_pe_1_1_1_n21,
         npu_inst_pe_1_1_1_n20, npu_inst_pe_1_1_1_n19, npu_inst_pe_1_1_1_n18,
         npu_inst_pe_1_1_1_n17, npu_inst_pe_1_1_1_n16, npu_inst_pe_1_1_1_n15,
         npu_inst_pe_1_1_1_n14, npu_inst_pe_1_1_1_n13, npu_inst_pe_1_1_1_n12,
         npu_inst_pe_1_1_1_n11, npu_inst_pe_1_1_1_n10, npu_inst_pe_1_1_1_n9,
         npu_inst_pe_1_1_1_n8, npu_inst_pe_1_1_1_n7, npu_inst_pe_1_1_1_n6,
         npu_inst_pe_1_1_1_n5, npu_inst_pe_1_1_1_n4, npu_inst_pe_1_1_1_n3,
         npu_inst_pe_1_1_1_n2, npu_inst_pe_1_1_1_n1,
         npu_inst_pe_1_1_1_sub_77_carry_7_, npu_inst_pe_1_1_1_sub_77_carry_6_,
         npu_inst_pe_1_1_1_sub_77_carry_5_, npu_inst_pe_1_1_1_sub_77_carry_4_,
         npu_inst_pe_1_1_1_sub_77_carry_3_, npu_inst_pe_1_1_1_sub_77_carry_2_,
         npu_inst_pe_1_1_1_sub_77_carry_1_, npu_inst_pe_1_1_1_add_79_carry_7_,
         npu_inst_pe_1_1_1_add_79_carry_6_, npu_inst_pe_1_1_1_add_79_carry_5_,
         npu_inst_pe_1_1_1_add_79_carry_4_, npu_inst_pe_1_1_1_add_79_carry_3_,
         npu_inst_pe_1_1_1_add_79_carry_2_, npu_inst_pe_1_1_1_add_79_carry_1_,
         npu_inst_pe_1_1_1_n97, npu_inst_pe_1_1_1_n96, npu_inst_pe_1_1_1_n95,
         npu_inst_pe_1_1_1_n94, npu_inst_pe_1_1_1_n93, npu_inst_pe_1_1_1_n92,
         npu_inst_pe_1_1_1_n91, npu_inst_pe_1_1_1_n90, npu_inst_pe_1_1_1_n89,
         npu_inst_pe_1_1_1_n88, npu_inst_pe_1_1_1_n87, npu_inst_pe_1_1_1_n86,
         npu_inst_pe_1_1_1_n85, npu_inst_pe_1_1_1_n84, npu_inst_pe_1_1_1_n83,
         npu_inst_pe_1_1_1_n82, npu_inst_pe_1_1_1_n81, npu_inst_pe_1_1_1_n80,
         npu_inst_pe_1_1_1_n79, npu_inst_pe_1_1_1_n78, npu_inst_pe_1_1_1_n77,
         npu_inst_pe_1_1_1_n76, npu_inst_pe_1_1_1_n75, npu_inst_pe_1_1_1_n74,
         npu_inst_pe_1_1_1_n73, npu_inst_pe_1_1_1_n72, npu_inst_pe_1_1_1_n71,
         npu_inst_pe_1_1_1_n70, npu_inst_pe_1_1_1_n69, npu_inst_pe_1_1_1_n68,
         npu_inst_pe_1_1_1_n67, npu_inst_pe_1_1_1_n66, npu_inst_pe_1_1_1_n65,
         npu_inst_pe_1_1_1_n64, npu_inst_pe_1_1_1_n63, npu_inst_pe_1_1_1_n62,
         npu_inst_pe_1_1_1_n61, npu_inst_pe_1_1_1_n60, npu_inst_pe_1_1_1_n59,
         npu_inst_pe_1_1_1_n58, npu_inst_pe_1_1_1_n57, npu_inst_pe_1_1_1_n56,
         npu_inst_pe_1_1_1_n55, npu_inst_pe_1_1_1_n54, npu_inst_pe_1_1_1_n53,
         npu_inst_pe_1_1_1_n52, npu_inst_pe_1_1_1_n51, npu_inst_pe_1_1_1_n50,
         npu_inst_pe_1_1_1_n49, npu_inst_pe_1_1_1_n48, npu_inst_pe_1_1_1_n47,
         npu_inst_pe_1_1_1_n46, npu_inst_pe_1_1_1_n45, npu_inst_pe_1_1_1_n44,
         npu_inst_pe_1_1_1_n43, npu_inst_pe_1_1_1_n42, npu_inst_pe_1_1_1_n41,
         npu_inst_pe_1_1_1_n40, npu_inst_pe_1_1_1_n39, npu_inst_pe_1_1_1_n38,
         npu_inst_pe_1_1_1_n37, npu_inst_pe_1_1_1_n27, npu_inst_pe_1_1_1_n26,
         npu_inst_pe_1_1_1_net4277, npu_inst_pe_1_1_1_net4271,
         npu_inst_pe_1_1_1_N94, npu_inst_pe_1_1_1_N93, npu_inst_pe_1_1_1_N84,
         npu_inst_pe_1_1_1_N80, npu_inst_pe_1_1_1_N79, npu_inst_pe_1_1_1_N78,
         npu_inst_pe_1_1_1_N77, npu_inst_pe_1_1_1_N76, npu_inst_pe_1_1_1_N75,
         npu_inst_pe_1_1_1_N74, npu_inst_pe_1_1_1_N73, npu_inst_pe_1_1_1_N72,
         npu_inst_pe_1_1_1_N71, npu_inst_pe_1_1_1_N70, npu_inst_pe_1_1_1_N69,
         npu_inst_pe_1_1_1_N68, npu_inst_pe_1_1_1_N67, npu_inst_pe_1_1_1_N66,
         npu_inst_pe_1_1_1_N65, npu_inst_pe_1_1_1_int_data_0_,
         npu_inst_pe_1_1_1_int_data_1_, npu_inst_pe_1_1_1_int_q_weight_0_,
         npu_inst_pe_1_1_1_int_q_weight_1_,
         npu_inst_pe_1_1_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_1_int_q_reg_h_0__1_, npu_inst_pe_1_1_2_n118,
         npu_inst_pe_1_1_2_n117, npu_inst_pe_1_1_2_n116,
         npu_inst_pe_1_1_2_n115, npu_inst_pe_1_1_2_n114,
         npu_inst_pe_1_1_2_n113, npu_inst_pe_1_1_2_n112,
         npu_inst_pe_1_1_2_n111, npu_inst_pe_1_1_2_n110,
         npu_inst_pe_1_1_2_n109, npu_inst_pe_1_1_2_n108,
         npu_inst_pe_1_1_2_n107, npu_inst_pe_1_1_2_n106,
         npu_inst_pe_1_1_2_n105, npu_inst_pe_1_1_2_n104,
         npu_inst_pe_1_1_2_n103, npu_inst_pe_1_1_2_n102,
         npu_inst_pe_1_1_2_n101, npu_inst_pe_1_1_2_n100, npu_inst_pe_1_1_2_n99,
         npu_inst_pe_1_1_2_n98, npu_inst_pe_1_1_2_n36, npu_inst_pe_1_1_2_n35,
         npu_inst_pe_1_1_2_n34, npu_inst_pe_1_1_2_n33, npu_inst_pe_1_1_2_n32,
         npu_inst_pe_1_1_2_n31, npu_inst_pe_1_1_2_n30, npu_inst_pe_1_1_2_n29,
         npu_inst_pe_1_1_2_n28, npu_inst_pe_1_1_2_n25, npu_inst_pe_1_1_2_n24,
         npu_inst_pe_1_1_2_n23, npu_inst_pe_1_1_2_n22, npu_inst_pe_1_1_2_n21,
         npu_inst_pe_1_1_2_n20, npu_inst_pe_1_1_2_n19, npu_inst_pe_1_1_2_n18,
         npu_inst_pe_1_1_2_n17, npu_inst_pe_1_1_2_n16, npu_inst_pe_1_1_2_n15,
         npu_inst_pe_1_1_2_n14, npu_inst_pe_1_1_2_n13, npu_inst_pe_1_1_2_n12,
         npu_inst_pe_1_1_2_n11, npu_inst_pe_1_1_2_n10, npu_inst_pe_1_1_2_n9,
         npu_inst_pe_1_1_2_n8, npu_inst_pe_1_1_2_n7, npu_inst_pe_1_1_2_n6,
         npu_inst_pe_1_1_2_n5, npu_inst_pe_1_1_2_n4, npu_inst_pe_1_1_2_n3,
         npu_inst_pe_1_1_2_n2, npu_inst_pe_1_1_2_n1,
         npu_inst_pe_1_1_2_sub_77_carry_7_, npu_inst_pe_1_1_2_sub_77_carry_6_,
         npu_inst_pe_1_1_2_sub_77_carry_5_, npu_inst_pe_1_1_2_sub_77_carry_4_,
         npu_inst_pe_1_1_2_sub_77_carry_3_, npu_inst_pe_1_1_2_sub_77_carry_2_,
         npu_inst_pe_1_1_2_sub_77_carry_1_, npu_inst_pe_1_1_2_add_79_carry_7_,
         npu_inst_pe_1_1_2_add_79_carry_6_, npu_inst_pe_1_1_2_add_79_carry_5_,
         npu_inst_pe_1_1_2_add_79_carry_4_, npu_inst_pe_1_1_2_add_79_carry_3_,
         npu_inst_pe_1_1_2_add_79_carry_2_, npu_inst_pe_1_1_2_add_79_carry_1_,
         npu_inst_pe_1_1_2_n97, npu_inst_pe_1_1_2_n96, npu_inst_pe_1_1_2_n95,
         npu_inst_pe_1_1_2_n94, npu_inst_pe_1_1_2_n93, npu_inst_pe_1_1_2_n92,
         npu_inst_pe_1_1_2_n91, npu_inst_pe_1_1_2_n90, npu_inst_pe_1_1_2_n89,
         npu_inst_pe_1_1_2_n88, npu_inst_pe_1_1_2_n87, npu_inst_pe_1_1_2_n86,
         npu_inst_pe_1_1_2_n85, npu_inst_pe_1_1_2_n84, npu_inst_pe_1_1_2_n83,
         npu_inst_pe_1_1_2_n82, npu_inst_pe_1_1_2_n81, npu_inst_pe_1_1_2_n80,
         npu_inst_pe_1_1_2_n79, npu_inst_pe_1_1_2_n78, npu_inst_pe_1_1_2_n77,
         npu_inst_pe_1_1_2_n76, npu_inst_pe_1_1_2_n75, npu_inst_pe_1_1_2_n74,
         npu_inst_pe_1_1_2_n73, npu_inst_pe_1_1_2_n72, npu_inst_pe_1_1_2_n71,
         npu_inst_pe_1_1_2_n70, npu_inst_pe_1_1_2_n69, npu_inst_pe_1_1_2_n68,
         npu_inst_pe_1_1_2_n67, npu_inst_pe_1_1_2_n66, npu_inst_pe_1_1_2_n65,
         npu_inst_pe_1_1_2_n64, npu_inst_pe_1_1_2_n63, npu_inst_pe_1_1_2_n62,
         npu_inst_pe_1_1_2_n61, npu_inst_pe_1_1_2_n60, npu_inst_pe_1_1_2_n59,
         npu_inst_pe_1_1_2_n58, npu_inst_pe_1_1_2_n57, npu_inst_pe_1_1_2_n56,
         npu_inst_pe_1_1_2_n55, npu_inst_pe_1_1_2_n54, npu_inst_pe_1_1_2_n53,
         npu_inst_pe_1_1_2_n52, npu_inst_pe_1_1_2_n51, npu_inst_pe_1_1_2_n50,
         npu_inst_pe_1_1_2_n49, npu_inst_pe_1_1_2_n48, npu_inst_pe_1_1_2_n47,
         npu_inst_pe_1_1_2_n46, npu_inst_pe_1_1_2_n45, npu_inst_pe_1_1_2_n44,
         npu_inst_pe_1_1_2_n43, npu_inst_pe_1_1_2_n42, npu_inst_pe_1_1_2_n41,
         npu_inst_pe_1_1_2_n40, npu_inst_pe_1_1_2_n39, npu_inst_pe_1_1_2_n38,
         npu_inst_pe_1_1_2_n37, npu_inst_pe_1_1_2_n27, npu_inst_pe_1_1_2_n26,
         npu_inst_pe_1_1_2_net4254, npu_inst_pe_1_1_2_net4248,
         npu_inst_pe_1_1_2_N94, npu_inst_pe_1_1_2_N93, npu_inst_pe_1_1_2_N84,
         npu_inst_pe_1_1_2_N80, npu_inst_pe_1_1_2_N79, npu_inst_pe_1_1_2_N78,
         npu_inst_pe_1_1_2_N77, npu_inst_pe_1_1_2_N76, npu_inst_pe_1_1_2_N75,
         npu_inst_pe_1_1_2_N74, npu_inst_pe_1_1_2_N73, npu_inst_pe_1_1_2_N72,
         npu_inst_pe_1_1_2_N71, npu_inst_pe_1_1_2_N70, npu_inst_pe_1_1_2_N69,
         npu_inst_pe_1_1_2_N68, npu_inst_pe_1_1_2_N67, npu_inst_pe_1_1_2_N66,
         npu_inst_pe_1_1_2_N65, npu_inst_pe_1_1_2_int_data_0_,
         npu_inst_pe_1_1_2_int_data_1_, npu_inst_pe_1_1_2_int_q_weight_0_,
         npu_inst_pe_1_1_2_int_q_weight_1_,
         npu_inst_pe_1_1_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_2_int_q_reg_h_0__1_, npu_inst_pe_1_1_3_n118,
         npu_inst_pe_1_1_3_n117, npu_inst_pe_1_1_3_n116,
         npu_inst_pe_1_1_3_n115, npu_inst_pe_1_1_3_n114,
         npu_inst_pe_1_1_3_n113, npu_inst_pe_1_1_3_n112,
         npu_inst_pe_1_1_3_n111, npu_inst_pe_1_1_3_n110,
         npu_inst_pe_1_1_3_n109, npu_inst_pe_1_1_3_n108,
         npu_inst_pe_1_1_3_n107, npu_inst_pe_1_1_3_n106,
         npu_inst_pe_1_1_3_n105, npu_inst_pe_1_1_3_n104,
         npu_inst_pe_1_1_3_n103, npu_inst_pe_1_1_3_n102,
         npu_inst_pe_1_1_3_n101, npu_inst_pe_1_1_3_n100, npu_inst_pe_1_1_3_n99,
         npu_inst_pe_1_1_3_n98, npu_inst_pe_1_1_3_n36, npu_inst_pe_1_1_3_n35,
         npu_inst_pe_1_1_3_n34, npu_inst_pe_1_1_3_n33, npu_inst_pe_1_1_3_n32,
         npu_inst_pe_1_1_3_n31, npu_inst_pe_1_1_3_n30, npu_inst_pe_1_1_3_n29,
         npu_inst_pe_1_1_3_n28, npu_inst_pe_1_1_3_n25, npu_inst_pe_1_1_3_n24,
         npu_inst_pe_1_1_3_n23, npu_inst_pe_1_1_3_n22, npu_inst_pe_1_1_3_n21,
         npu_inst_pe_1_1_3_n20, npu_inst_pe_1_1_3_n19, npu_inst_pe_1_1_3_n18,
         npu_inst_pe_1_1_3_n17, npu_inst_pe_1_1_3_n16, npu_inst_pe_1_1_3_n15,
         npu_inst_pe_1_1_3_n14, npu_inst_pe_1_1_3_n13, npu_inst_pe_1_1_3_n12,
         npu_inst_pe_1_1_3_n11, npu_inst_pe_1_1_3_n10, npu_inst_pe_1_1_3_n9,
         npu_inst_pe_1_1_3_n8, npu_inst_pe_1_1_3_n7, npu_inst_pe_1_1_3_n6,
         npu_inst_pe_1_1_3_n5, npu_inst_pe_1_1_3_n4, npu_inst_pe_1_1_3_n3,
         npu_inst_pe_1_1_3_n2, npu_inst_pe_1_1_3_n1,
         npu_inst_pe_1_1_3_sub_77_carry_7_, npu_inst_pe_1_1_3_sub_77_carry_6_,
         npu_inst_pe_1_1_3_sub_77_carry_5_, npu_inst_pe_1_1_3_sub_77_carry_4_,
         npu_inst_pe_1_1_3_sub_77_carry_3_, npu_inst_pe_1_1_3_sub_77_carry_2_,
         npu_inst_pe_1_1_3_sub_77_carry_1_, npu_inst_pe_1_1_3_add_79_carry_7_,
         npu_inst_pe_1_1_3_add_79_carry_6_, npu_inst_pe_1_1_3_add_79_carry_5_,
         npu_inst_pe_1_1_3_add_79_carry_4_, npu_inst_pe_1_1_3_add_79_carry_3_,
         npu_inst_pe_1_1_3_add_79_carry_2_, npu_inst_pe_1_1_3_add_79_carry_1_,
         npu_inst_pe_1_1_3_n97, npu_inst_pe_1_1_3_n96, npu_inst_pe_1_1_3_n95,
         npu_inst_pe_1_1_3_n94, npu_inst_pe_1_1_3_n93, npu_inst_pe_1_1_3_n92,
         npu_inst_pe_1_1_3_n91, npu_inst_pe_1_1_3_n90, npu_inst_pe_1_1_3_n89,
         npu_inst_pe_1_1_3_n88, npu_inst_pe_1_1_3_n87, npu_inst_pe_1_1_3_n86,
         npu_inst_pe_1_1_3_n85, npu_inst_pe_1_1_3_n84, npu_inst_pe_1_1_3_n83,
         npu_inst_pe_1_1_3_n82, npu_inst_pe_1_1_3_n81, npu_inst_pe_1_1_3_n80,
         npu_inst_pe_1_1_3_n79, npu_inst_pe_1_1_3_n78, npu_inst_pe_1_1_3_n77,
         npu_inst_pe_1_1_3_n76, npu_inst_pe_1_1_3_n75, npu_inst_pe_1_1_3_n74,
         npu_inst_pe_1_1_3_n73, npu_inst_pe_1_1_3_n72, npu_inst_pe_1_1_3_n71,
         npu_inst_pe_1_1_3_n70, npu_inst_pe_1_1_3_n69, npu_inst_pe_1_1_3_n68,
         npu_inst_pe_1_1_3_n67, npu_inst_pe_1_1_3_n66, npu_inst_pe_1_1_3_n65,
         npu_inst_pe_1_1_3_n64, npu_inst_pe_1_1_3_n63, npu_inst_pe_1_1_3_n62,
         npu_inst_pe_1_1_3_n61, npu_inst_pe_1_1_3_n60, npu_inst_pe_1_1_3_n59,
         npu_inst_pe_1_1_3_n58, npu_inst_pe_1_1_3_n57, npu_inst_pe_1_1_3_n56,
         npu_inst_pe_1_1_3_n55, npu_inst_pe_1_1_3_n54, npu_inst_pe_1_1_3_n53,
         npu_inst_pe_1_1_3_n52, npu_inst_pe_1_1_3_n51, npu_inst_pe_1_1_3_n50,
         npu_inst_pe_1_1_3_n49, npu_inst_pe_1_1_3_n48, npu_inst_pe_1_1_3_n47,
         npu_inst_pe_1_1_3_n46, npu_inst_pe_1_1_3_n45, npu_inst_pe_1_1_3_n44,
         npu_inst_pe_1_1_3_n43, npu_inst_pe_1_1_3_n42, npu_inst_pe_1_1_3_n41,
         npu_inst_pe_1_1_3_n40, npu_inst_pe_1_1_3_n39, npu_inst_pe_1_1_3_n38,
         npu_inst_pe_1_1_3_n37, npu_inst_pe_1_1_3_n27, npu_inst_pe_1_1_3_n26,
         npu_inst_pe_1_1_3_net4231, npu_inst_pe_1_1_3_net4225,
         npu_inst_pe_1_1_3_N94, npu_inst_pe_1_1_3_N93, npu_inst_pe_1_1_3_N84,
         npu_inst_pe_1_1_3_N80, npu_inst_pe_1_1_3_N79, npu_inst_pe_1_1_3_N78,
         npu_inst_pe_1_1_3_N77, npu_inst_pe_1_1_3_N76, npu_inst_pe_1_1_3_N75,
         npu_inst_pe_1_1_3_N74, npu_inst_pe_1_1_3_N73, npu_inst_pe_1_1_3_N72,
         npu_inst_pe_1_1_3_N71, npu_inst_pe_1_1_3_N70, npu_inst_pe_1_1_3_N69,
         npu_inst_pe_1_1_3_N68, npu_inst_pe_1_1_3_N67, npu_inst_pe_1_1_3_N66,
         npu_inst_pe_1_1_3_N65, npu_inst_pe_1_1_3_int_data_0_,
         npu_inst_pe_1_1_3_int_data_1_, npu_inst_pe_1_1_3_int_q_weight_0_,
         npu_inst_pe_1_1_3_int_q_weight_1_,
         npu_inst_pe_1_1_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_3_int_q_reg_h_0__1_, npu_inst_pe_1_1_4_n118,
         npu_inst_pe_1_1_4_n117, npu_inst_pe_1_1_4_n116,
         npu_inst_pe_1_1_4_n115, npu_inst_pe_1_1_4_n114,
         npu_inst_pe_1_1_4_n113, npu_inst_pe_1_1_4_n112,
         npu_inst_pe_1_1_4_n111, npu_inst_pe_1_1_4_n110,
         npu_inst_pe_1_1_4_n109, npu_inst_pe_1_1_4_n108,
         npu_inst_pe_1_1_4_n107, npu_inst_pe_1_1_4_n106,
         npu_inst_pe_1_1_4_n105, npu_inst_pe_1_1_4_n104,
         npu_inst_pe_1_1_4_n103, npu_inst_pe_1_1_4_n102,
         npu_inst_pe_1_1_4_n101, npu_inst_pe_1_1_4_n100, npu_inst_pe_1_1_4_n99,
         npu_inst_pe_1_1_4_n98, npu_inst_pe_1_1_4_n36, npu_inst_pe_1_1_4_n35,
         npu_inst_pe_1_1_4_n34, npu_inst_pe_1_1_4_n33, npu_inst_pe_1_1_4_n32,
         npu_inst_pe_1_1_4_n31, npu_inst_pe_1_1_4_n30, npu_inst_pe_1_1_4_n29,
         npu_inst_pe_1_1_4_n28, npu_inst_pe_1_1_4_n25, npu_inst_pe_1_1_4_n24,
         npu_inst_pe_1_1_4_n23, npu_inst_pe_1_1_4_n22, npu_inst_pe_1_1_4_n21,
         npu_inst_pe_1_1_4_n20, npu_inst_pe_1_1_4_n19, npu_inst_pe_1_1_4_n18,
         npu_inst_pe_1_1_4_n17, npu_inst_pe_1_1_4_n16, npu_inst_pe_1_1_4_n15,
         npu_inst_pe_1_1_4_n14, npu_inst_pe_1_1_4_n13, npu_inst_pe_1_1_4_n12,
         npu_inst_pe_1_1_4_n11, npu_inst_pe_1_1_4_n10, npu_inst_pe_1_1_4_n9,
         npu_inst_pe_1_1_4_n8, npu_inst_pe_1_1_4_n7, npu_inst_pe_1_1_4_n6,
         npu_inst_pe_1_1_4_n5, npu_inst_pe_1_1_4_n4, npu_inst_pe_1_1_4_n3,
         npu_inst_pe_1_1_4_n2, npu_inst_pe_1_1_4_n1,
         npu_inst_pe_1_1_4_sub_77_carry_7_, npu_inst_pe_1_1_4_sub_77_carry_6_,
         npu_inst_pe_1_1_4_sub_77_carry_5_, npu_inst_pe_1_1_4_sub_77_carry_4_,
         npu_inst_pe_1_1_4_sub_77_carry_3_, npu_inst_pe_1_1_4_sub_77_carry_2_,
         npu_inst_pe_1_1_4_sub_77_carry_1_, npu_inst_pe_1_1_4_add_79_carry_7_,
         npu_inst_pe_1_1_4_add_79_carry_6_, npu_inst_pe_1_1_4_add_79_carry_5_,
         npu_inst_pe_1_1_4_add_79_carry_4_, npu_inst_pe_1_1_4_add_79_carry_3_,
         npu_inst_pe_1_1_4_add_79_carry_2_, npu_inst_pe_1_1_4_add_79_carry_1_,
         npu_inst_pe_1_1_4_n97, npu_inst_pe_1_1_4_n96, npu_inst_pe_1_1_4_n95,
         npu_inst_pe_1_1_4_n94, npu_inst_pe_1_1_4_n93, npu_inst_pe_1_1_4_n92,
         npu_inst_pe_1_1_4_n91, npu_inst_pe_1_1_4_n90, npu_inst_pe_1_1_4_n89,
         npu_inst_pe_1_1_4_n88, npu_inst_pe_1_1_4_n87, npu_inst_pe_1_1_4_n86,
         npu_inst_pe_1_1_4_n85, npu_inst_pe_1_1_4_n84, npu_inst_pe_1_1_4_n83,
         npu_inst_pe_1_1_4_n82, npu_inst_pe_1_1_4_n81, npu_inst_pe_1_1_4_n80,
         npu_inst_pe_1_1_4_n79, npu_inst_pe_1_1_4_n78, npu_inst_pe_1_1_4_n77,
         npu_inst_pe_1_1_4_n76, npu_inst_pe_1_1_4_n75, npu_inst_pe_1_1_4_n74,
         npu_inst_pe_1_1_4_n73, npu_inst_pe_1_1_4_n72, npu_inst_pe_1_1_4_n71,
         npu_inst_pe_1_1_4_n70, npu_inst_pe_1_1_4_n69, npu_inst_pe_1_1_4_n68,
         npu_inst_pe_1_1_4_n67, npu_inst_pe_1_1_4_n66, npu_inst_pe_1_1_4_n65,
         npu_inst_pe_1_1_4_n64, npu_inst_pe_1_1_4_n63, npu_inst_pe_1_1_4_n62,
         npu_inst_pe_1_1_4_n61, npu_inst_pe_1_1_4_n60, npu_inst_pe_1_1_4_n59,
         npu_inst_pe_1_1_4_n58, npu_inst_pe_1_1_4_n57, npu_inst_pe_1_1_4_n56,
         npu_inst_pe_1_1_4_n55, npu_inst_pe_1_1_4_n54, npu_inst_pe_1_1_4_n53,
         npu_inst_pe_1_1_4_n52, npu_inst_pe_1_1_4_n51, npu_inst_pe_1_1_4_n50,
         npu_inst_pe_1_1_4_n49, npu_inst_pe_1_1_4_n48, npu_inst_pe_1_1_4_n47,
         npu_inst_pe_1_1_4_n46, npu_inst_pe_1_1_4_n45, npu_inst_pe_1_1_4_n44,
         npu_inst_pe_1_1_4_n43, npu_inst_pe_1_1_4_n42, npu_inst_pe_1_1_4_n41,
         npu_inst_pe_1_1_4_n40, npu_inst_pe_1_1_4_n39, npu_inst_pe_1_1_4_n38,
         npu_inst_pe_1_1_4_n37, npu_inst_pe_1_1_4_n27, npu_inst_pe_1_1_4_n26,
         npu_inst_pe_1_1_4_net4208, npu_inst_pe_1_1_4_net4202,
         npu_inst_pe_1_1_4_N94, npu_inst_pe_1_1_4_N93, npu_inst_pe_1_1_4_N84,
         npu_inst_pe_1_1_4_N80, npu_inst_pe_1_1_4_N79, npu_inst_pe_1_1_4_N78,
         npu_inst_pe_1_1_4_N77, npu_inst_pe_1_1_4_N76, npu_inst_pe_1_1_4_N75,
         npu_inst_pe_1_1_4_N74, npu_inst_pe_1_1_4_N73, npu_inst_pe_1_1_4_N72,
         npu_inst_pe_1_1_4_N71, npu_inst_pe_1_1_4_N70, npu_inst_pe_1_1_4_N69,
         npu_inst_pe_1_1_4_N68, npu_inst_pe_1_1_4_N67, npu_inst_pe_1_1_4_N66,
         npu_inst_pe_1_1_4_N65, npu_inst_pe_1_1_4_int_data_0_,
         npu_inst_pe_1_1_4_int_data_1_, npu_inst_pe_1_1_4_int_q_weight_0_,
         npu_inst_pe_1_1_4_int_q_weight_1_,
         npu_inst_pe_1_1_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_4_int_q_reg_h_0__1_, npu_inst_pe_1_1_5_n118,
         npu_inst_pe_1_1_5_n117, npu_inst_pe_1_1_5_n116,
         npu_inst_pe_1_1_5_n115, npu_inst_pe_1_1_5_n114,
         npu_inst_pe_1_1_5_n113, npu_inst_pe_1_1_5_n112,
         npu_inst_pe_1_1_5_n111, npu_inst_pe_1_1_5_n110,
         npu_inst_pe_1_1_5_n109, npu_inst_pe_1_1_5_n108,
         npu_inst_pe_1_1_5_n107, npu_inst_pe_1_1_5_n106,
         npu_inst_pe_1_1_5_n105, npu_inst_pe_1_1_5_n104,
         npu_inst_pe_1_1_5_n103, npu_inst_pe_1_1_5_n102,
         npu_inst_pe_1_1_5_n101, npu_inst_pe_1_1_5_n100, npu_inst_pe_1_1_5_n99,
         npu_inst_pe_1_1_5_n98, npu_inst_pe_1_1_5_n36, npu_inst_pe_1_1_5_n35,
         npu_inst_pe_1_1_5_n34, npu_inst_pe_1_1_5_n33, npu_inst_pe_1_1_5_n32,
         npu_inst_pe_1_1_5_n31, npu_inst_pe_1_1_5_n30, npu_inst_pe_1_1_5_n29,
         npu_inst_pe_1_1_5_n28, npu_inst_pe_1_1_5_n25, npu_inst_pe_1_1_5_n24,
         npu_inst_pe_1_1_5_n23, npu_inst_pe_1_1_5_n22, npu_inst_pe_1_1_5_n21,
         npu_inst_pe_1_1_5_n20, npu_inst_pe_1_1_5_n19, npu_inst_pe_1_1_5_n18,
         npu_inst_pe_1_1_5_n17, npu_inst_pe_1_1_5_n16, npu_inst_pe_1_1_5_n15,
         npu_inst_pe_1_1_5_n14, npu_inst_pe_1_1_5_n13, npu_inst_pe_1_1_5_n12,
         npu_inst_pe_1_1_5_n11, npu_inst_pe_1_1_5_n10, npu_inst_pe_1_1_5_n9,
         npu_inst_pe_1_1_5_n8, npu_inst_pe_1_1_5_n7, npu_inst_pe_1_1_5_n6,
         npu_inst_pe_1_1_5_n5, npu_inst_pe_1_1_5_n4, npu_inst_pe_1_1_5_n3,
         npu_inst_pe_1_1_5_n2, npu_inst_pe_1_1_5_n1,
         npu_inst_pe_1_1_5_sub_77_carry_7_, npu_inst_pe_1_1_5_sub_77_carry_6_,
         npu_inst_pe_1_1_5_sub_77_carry_5_, npu_inst_pe_1_1_5_sub_77_carry_4_,
         npu_inst_pe_1_1_5_sub_77_carry_3_, npu_inst_pe_1_1_5_sub_77_carry_2_,
         npu_inst_pe_1_1_5_sub_77_carry_1_, npu_inst_pe_1_1_5_add_79_carry_7_,
         npu_inst_pe_1_1_5_add_79_carry_6_, npu_inst_pe_1_1_5_add_79_carry_5_,
         npu_inst_pe_1_1_5_add_79_carry_4_, npu_inst_pe_1_1_5_add_79_carry_3_,
         npu_inst_pe_1_1_5_add_79_carry_2_, npu_inst_pe_1_1_5_add_79_carry_1_,
         npu_inst_pe_1_1_5_n97, npu_inst_pe_1_1_5_n96, npu_inst_pe_1_1_5_n95,
         npu_inst_pe_1_1_5_n94, npu_inst_pe_1_1_5_n93, npu_inst_pe_1_1_5_n92,
         npu_inst_pe_1_1_5_n91, npu_inst_pe_1_1_5_n90, npu_inst_pe_1_1_5_n89,
         npu_inst_pe_1_1_5_n88, npu_inst_pe_1_1_5_n87, npu_inst_pe_1_1_5_n86,
         npu_inst_pe_1_1_5_n85, npu_inst_pe_1_1_5_n84, npu_inst_pe_1_1_5_n83,
         npu_inst_pe_1_1_5_n82, npu_inst_pe_1_1_5_n81, npu_inst_pe_1_1_5_n80,
         npu_inst_pe_1_1_5_n79, npu_inst_pe_1_1_5_n78, npu_inst_pe_1_1_5_n77,
         npu_inst_pe_1_1_5_n76, npu_inst_pe_1_1_5_n75, npu_inst_pe_1_1_5_n74,
         npu_inst_pe_1_1_5_n73, npu_inst_pe_1_1_5_n72, npu_inst_pe_1_1_5_n71,
         npu_inst_pe_1_1_5_n70, npu_inst_pe_1_1_5_n69, npu_inst_pe_1_1_5_n68,
         npu_inst_pe_1_1_5_n67, npu_inst_pe_1_1_5_n66, npu_inst_pe_1_1_5_n65,
         npu_inst_pe_1_1_5_n64, npu_inst_pe_1_1_5_n63, npu_inst_pe_1_1_5_n62,
         npu_inst_pe_1_1_5_n61, npu_inst_pe_1_1_5_n60, npu_inst_pe_1_1_5_n59,
         npu_inst_pe_1_1_5_n58, npu_inst_pe_1_1_5_n57, npu_inst_pe_1_1_5_n56,
         npu_inst_pe_1_1_5_n55, npu_inst_pe_1_1_5_n54, npu_inst_pe_1_1_5_n53,
         npu_inst_pe_1_1_5_n52, npu_inst_pe_1_1_5_n51, npu_inst_pe_1_1_5_n50,
         npu_inst_pe_1_1_5_n49, npu_inst_pe_1_1_5_n48, npu_inst_pe_1_1_5_n47,
         npu_inst_pe_1_1_5_n46, npu_inst_pe_1_1_5_n45, npu_inst_pe_1_1_5_n44,
         npu_inst_pe_1_1_5_n43, npu_inst_pe_1_1_5_n42, npu_inst_pe_1_1_5_n41,
         npu_inst_pe_1_1_5_n40, npu_inst_pe_1_1_5_n39, npu_inst_pe_1_1_5_n38,
         npu_inst_pe_1_1_5_n37, npu_inst_pe_1_1_5_n27, npu_inst_pe_1_1_5_n26,
         npu_inst_pe_1_1_5_net4185, npu_inst_pe_1_1_5_net4179,
         npu_inst_pe_1_1_5_N94, npu_inst_pe_1_1_5_N93, npu_inst_pe_1_1_5_N84,
         npu_inst_pe_1_1_5_N80, npu_inst_pe_1_1_5_N79, npu_inst_pe_1_1_5_N78,
         npu_inst_pe_1_1_5_N77, npu_inst_pe_1_1_5_N76, npu_inst_pe_1_1_5_N75,
         npu_inst_pe_1_1_5_N74, npu_inst_pe_1_1_5_N73, npu_inst_pe_1_1_5_N72,
         npu_inst_pe_1_1_5_N71, npu_inst_pe_1_1_5_N70, npu_inst_pe_1_1_5_N69,
         npu_inst_pe_1_1_5_N68, npu_inst_pe_1_1_5_N67, npu_inst_pe_1_1_5_N66,
         npu_inst_pe_1_1_5_N65, npu_inst_pe_1_1_5_int_data_0_,
         npu_inst_pe_1_1_5_int_data_1_, npu_inst_pe_1_1_5_int_q_weight_0_,
         npu_inst_pe_1_1_5_int_q_weight_1_,
         npu_inst_pe_1_1_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_5_int_q_reg_h_0__1_, npu_inst_pe_1_1_6_n118,
         npu_inst_pe_1_1_6_n117, npu_inst_pe_1_1_6_n116,
         npu_inst_pe_1_1_6_n115, npu_inst_pe_1_1_6_n114,
         npu_inst_pe_1_1_6_n113, npu_inst_pe_1_1_6_n112,
         npu_inst_pe_1_1_6_n111, npu_inst_pe_1_1_6_n110,
         npu_inst_pe_1_1_6_n109, npu_inst_pe_1_1_6_n108,
         npu_inst_pe_1_1_6_n107, npu_inst_pe_1_1_6_n106,
         npu_inst_pe_1_1_6_n105, npu_inst_pe_1_1_6_n104,
         npu_inst_pe_1_1_6_n103, npu_inst_pe_1_1_6_n102,
         npu_inst_pe_1_1_6_n101, npu_inst_pe_1_1_6_n100, npu_inst_pe_1_1_6_n99,
         npu_inst_pe_1_1_6_n98, npu_inst_pe_1_1_6_n36, npu_inst_pe_1_1_6_n35,
         npu_inst_pe_1_1_6_n34, npu_inst_pe_1_1_6_n33, npu_inst_pe_1_1_6_n32,
         npu_inst_pe_1_1_6_n31, npu_inst_pe_1_1_6_n30, npu_inst_pe_1_1_6_n29,
         npu_inst_pe_1_1_6_n28, npu_inst_pe_1_1_6_n25, npu_inst_pe_1_1_6_n24,
         npu_inst_pe_1_1_6_n23, npu_inst_pe_1_1_6_n22, npu_inst_pe_1_1_6_n21,
         npu_inst_pe_1_1_6_n20, npu_inst_pe_1_1_6_n19, npu_inst_pe_1_1_6_n18,
         npu_inst_pe_1_1_6_n17, npu_inst_pe_1_1_6_n16, npu_inst_pe_1_1_6_n15,
         npu_inst_pe_1_1_6_n14, npu_inst_pe_1_1_6_n13, npu_inst_pe_1_1_6_n12,
         npu_inst_pe_1_1_6_n11, npu_inst_pe_1_1_6_n10, npu_inst_pe_1_1_6_n9,
         npu_inst_pe_1_1_6_n8, npu_inst_pe_1_1_6_n7, npu_inst_pe_1_1_6_n6,
         npu_inst_pe_1_1_6_n5, npu_inst_pe_1_1_6_n4, npu_inst_pe_1_1_6_n3,
         npu_inst_pe_1_1_6_n2, npu_inst_pe_1_1_6_n1,
         npu_inst_pe_1_1_6_sub_77_carry_7_, npu_inst_pe_1_1_6_sub_77_carry_6_,
         npu_inst_pe_1_1_6_sub_77_carry_5_, npu_inst_pe_1_1_6_sub_77_carry_4_,
         npu_inst_pe_1_1_6_sub_77_carry_3_, npu_inst_pe_1_1_6_sub_77_carry_2_,
         npu_inst_pe_1_1_6_sub_77_carry_1_, npu_inst_pe_1_1_6_add_79_carry_7_,
         npu_inst_pe_1_1_6_add_79_carry_6_, npu_inst_pe_1_1_6_add_79_carry_5_,
         npu_inst_pe_1_1_6_add_79_carry_4_, npu_inst_pe_1_1_6_add_79_carry_3_,
         npu_inst_pe_1_1_6_add_79_carry_2_, npu_inst_pe_1_1_6_add_79_carry_1_,
         npu_inst_pe_1_1_6_n97, npu_inst_pe_1_1_6_n96, npu_inst_pe_1_1_6_n95,
         npu_inst_pe_1_1_6_n94, npu_inst_pe_1_1_6_n93, npu_inst_pe_1_1_6_n92,
         npu_inst_pe_1_1_6_n91, npu_inst_pe_1_1_6_n90, npu_inst_pe_1_1_6_n89,
         npu_inst_pe_1_1_6_n88, npu_inst_pe_1_1_6_n87, npu_inst_pe_1_1_6_n86,
         npu_inst_pe_1_1_6_n85, npu_inst_pe_1_1_6_n84, npu_inst_pe_1_1_6_n83,
         npu_inst_pe_1_1_6_n82, npu_inst_pe_1_1_6_n81, npu_inst_pe_1_1_6_n80,
         npu_inst_pe_1_1_6_n79, npu_inst_pe_1_1_6_n78, npu_inst_pe_1_1_6_n77,
         npu_inst_pe_1_1_6_n76, npu_inst_pe_1_1_6_n75, npu_inst_pe_1_1_6_n74,
         npu_inst_pe_1_1_6_n73, npu_inst_pe_1_1_6_n72, npu_inst_pe_1_1_6_n71,
         npu_inst_pe_1_1_6_n70, npu_inst_pe_1_1_6_n69, npu_inst_pe_1_1_6_n68,
         npu_inst_pe_1_1_6_n67, npu_inst_pe_1_1_6_n66, npu_inst_pe_1_1_6_n65,
         npu_inst_pe_1_1_6_n64, npu_inst_pe_1_1_6_n63, npu_inst_pe_1_1_6_n62,
         npu_inst_pe_1_1_6_n61, npu_inst_pe_1_1_6_n60, npu_inst_pe_1_1_6_n59,
         npu_inst_pe_1_1_6_n58, npu_inst_pe_1_1_6_n57, npu_inst_pe_1_1_6_n56,
         npu_inst_pe_1_1_6_n55, npu_inst_pe_1_1_6_n54, npu_inst_pe_1_1_6_n53,
         npu_inst_pe_1_1_6_n52, npu_inst_pe_1_1_6_n51, npu_inst_pe_1_1_6_n50,
         npu_inst_pe_1_1_6_n49, npu_inst_pe_1_1_6_n48, npu_inst_pe_1_1_6_n47,
         npu_inst_pe_1_1_6_n46, npu_inst_pe_1_1_6_n45, npu_inst_pe_1_1_6_n44,
         npu_inst_pe_1_1_6_n43, npu_inst_pe_1_1_6_n42, npu_inst_pe_1_1_6_n41,
         npu_inst_pe_1_1_6_n40, npu_inst_pe_1_1_6_n39, npu_inst_pe_1_1_6_n38,
         npu_inst_pe_1_1_6_n37, npu_inst_pe_1_1_6_n27, npu_inst_pe_1_1_6_n26,
         npu_inst_pe_1_1_6_net4162, npu_inst_pe_1_1_6_net4156,
         npu_inst_pe_1_1_6_N94, npu_inst_pe_1_1_6_N93, npu_inst_pe_1_1_6_N84,
         npu_inst_pe_1_1_6_N80, npu_inst_pe_1_1_6_N79, npu_inst_pe_1_1_6_N78,
         npu_inst_pe_1_1_6_N77, npu_inst_pe_1_1_6_N76, npu_inst_pe_1_1_6_N75,
         npu_inst_pe_1_1_6_N74, npu_inst_pe_1_1_6_N73, npu_inst_pe_1_1_6_N72,
         npu_inst_pe_1_1_6_N71, npu_inst_pe_1_1_6_N70, npu_inst_pe_1_1_6_N69,
         npu_inst_pe_1_1_6_N68, npu_inst_pe_1_1_6_N67, npu_inst_pe_1_1_6_N66,
         npu_inst_pe_1_1_6_N65, npu_inst_pe_1_1_6_int_data_0_,
         npu_inst_pe_1_1_6_int_data_1_, npu_inst_pe_1_1_6_int_q_weight_0_,
         npu_inst_pe_1_1_6_int_q_weight_1_,
         npu_inst_pe_1_1_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_6_int_q_reg_h_0__1_, npu_inst_pe_1_1_7_n118,
         npu_inst_pe_1_1_7_n117, npu_inst_pe_1_1_7_n116,
         npu_inst_pe_1_1_7_n115, npu_inst_pe_1_1_7_n114,
         npu_inst_pe_1_1_7_n113, npu_inst_pe_1_1_7_n112,
         npu_inst_pe_1_1_7_n111, npu_inst_pe_1_1_7_n110,
         npu_inst_pe_1_1_7_n109, npu_inst_pe_1_1_7_n108,
         npu_inst_pe_1_1_7_n107, npu_inst_pe_1_1_7_n106,
         npu_inst_pe_1_1_7_n105, npu_inst_pe_1_1_7_n104,
         npu_inst_pe_1_1_7_n103, npu_inst_pe_1_1_7_n102,
         npu_inst_pe_1_1_7_n101, npu_inst_pe_1_1_7_n100, npu_inst_pe_1_1_7_n99,
         npu_inst_pe_1_1_7_n98, npu_inst_pe_1_1_7_n36, npu_inst_pe_1_1_7_n35,
         npu_inst_pe_1_1_7_n34, npu_inst_pe_1_1_7_n33, npu_inst_pe_1_1_7_n32,
         npu_inst_pe_1_1_7_n31, npu_inst_pe_1_1_7_n30, npu_inst_pe_1_1_7_n29,
         npu_inst_pe_1_1_7_n28, npu_inst_pe_1_1_7_n25, npu_inst_pe_1_1_7_n24,
         npu_inst_pe_1_1_7_n23, npu_inst_pe_1_1_7_n22, npu_inst_pe_1_1_7_n21,
         npu_inst_pe_1_1_7_n20, npu_inst_pe_1_1_7_n19, npu_inst_pe_1_1_7_n18,
         npu_inst_pe_1_1_7_n17, npu_inst_pe_1_1_7_n16, npu_inst_pe_1_1_7_n15,
         npu_inst_pe_1_1_7_n14, npu_inst_pe_1_1_7_n13, npu_inst_pe_1_1_7_n12,
         npu_inst_pe_1_1_7_n11, npu_inst_pe_1_1_7_n10, npu_inst_pe_1_1_7_n9,
         npu_inst_pe_1_1_7_n8, npu_inst_pe_1_1_7_n7, npu_inst_pe_1_1_7_n6,
         npu_inst_pe_1_1_7_n5, npu_inst_pe_1_1_7_n4, npu_inst_pe_1_1_7_n3,
         npu_inst_pe_1_1_7_n2, npu_inst_pe_1_1_7_n1,
         npu_inst_pe_1_1_7_sub_77_carry_7_, npu_inst_pe_1_1_7_sub_77_carry_6_,
         npu_inst_pe_1_1_7_sub_77_carry_5_, npu_inst_pe_1_1_7_sub_77_carry_4_,
         npu_inst_pe_1_1_7_sub_77_carry_3_, npu_inst_pe_1_1_7_sub_77_carry_2_,
         npu_inst_pe_1_1_7_sub_77_carry_1_, npu_inst_pe_1_1_7_add_79_carry_7_,
         npu_inst_pe_1_1_7_add_79_carry_6_, npu_inst_pe_1_1_7_add_79_carry_5_,
         npu_inst_pe_1_1_7_add_79_carry_4_, npu_inst_pe_1_1_7_add_79_carry_3_,
         npu_inst_pe_1_1_7_add_79_carry_2_, npu_inst_pe_1_1_7_add_79_carry_1_,
         npu_inst_pe_1_1_7_n97, npu_inst_pe_1_1_7_n96, npu_inst_pe_1_1_7_n95,
         npu_inst_pe_1_1_7_n94, npu_inst_pe_1_1_7_n93, npu_inst_pe_1_1_7_n92,
         npu_inst_pe_1_1_7_n91, npu_inst_pe_1_1_7_n90, npu_inst_pe_1_1_7_n89,
         npu_inst_pe_1_1_7_n88, npu_inst_pe_1_1_7_n87, npu_inst_pe_1_1_7_n86,
         npu_inst_pe_1_1_7_n85, npu_inst_pe_1_1_7_n84, npu_inst_pe_1_1_7_n83,
         npu_inst_pe_1_1_7_n82, npu_inst_pe_1_1_7_n81, npu_inst_pe_1_1_7_n80,
         npu_inst_pe_1_1_7_n79, npu_inst_pe_1_1_7_n78, npu_inst_pe_1_1_7_n77,
         npu_inst_pe_1_1_7_n76, npu_inst_pe_1_1_7_n75, npu_inst_pe_1_1_7_n74,
         npu_inst_pe_1_1_7_n73, npu_inst_pe_1_1_7_n72, npu_inst_pe_1_1_7_n71,
         npu_inst_pe_1_1_7_n70, npu_inst_pe_1_1_7_n69, npu_inst_pe_1_1_7_n68,
         npu_inst_pe_1_1_7_n67, npu_inst_pe_1_1_7_n66, npu_inst_pe_1_1_7_n65,
         npu_inst_pe_1_1_7_n64, npu_inst_pe_1_1_7_n63, npu_inst_pe_1_1_7_n62,
         npu_inst_pe_1_1_7_n61, npu_inst_pe_1_1_7_n60, npu_inst_pe_1_1_7_n59,
         npu_inst_pe_1_1_7_n58, npu_inst_pe_1_1_7_n57, npu_inst_pe_1_1_7_n56,
         npu_inst_pe_1_1_7_n55, npu_inst_pe_1_1_7_n54, npu_inst_pe_1_1_7_n53,
         npu_inst_pe_1_1_7_n52, npu_inst_pe_1_1_7_n51, npu_inst_pe_1_1_7_n50,
         npu_inst_pe_1_1_7_n49, npu_inst_pe_1_1_7_n48, npu_inst_pe_1_1_7_n47,
         npu_inst_pe_1_1_7_n46, npu_inst_pe_1_1_7_n45, npu_inst_pe_1_1_7_n44,
         npu_inst_pe_1_1_7_n43, npu_inst_pe_1_1_7_n42, npu_inst_pe_1_1_7_n41,
         npu_inst_pe_1_1_7_n40, npu_inst_pe_1_1_7_n39, npu_inst_pe_1_1_7_n38,
         npu_inst_pe_1_1_7_n37, npu_inst_pe_1_1_7_n27, npu_inst_pe_1_1_7_n26,
         npu_inst_pe_1_1_7_net4139, npu_inst_pe_1_1_7_net4133,
         npu_inst_pe_1_1_7_N94, npu_inst_pe_1_1_7_N93, npu_inst_pe_1_1_7_N84,
         npu_inst_pe_1_1_7_N80, npu_inst_pe_1_1_7_N79, npu_inst_pe_1_1_7_N78,
         npu_inst_pe_1_1_7_N77, npu_inst_pe_1_1_7_N76, npu_inst_pe_1_1_7_N75,
         npu_inst_pe_1_1_7_N74, npu_inst_pe_1_1_7_N73, npu_inst_pe_1_1_7_N72,
         npu_inst_pe_1_1_7_N71, npu_inst_pe_1_1_7_N70, npu_inst_pe_1_1_7_N69,
         npu_inst_pe_1_1_7_N68, npu_inst_pe_1_1_7_N67, npu_inst_pe_1_1_7_N66,
         npu_inst_pe_1_1_7_N65, npu_inst_pe_1_1_7_int_data_0_,
         npu_inst_pe_1_1_7_int_data_1_, npu_inst_pe_1_1_7_int_q_weight_0_,
         npu_inst_pe_1_1_7_int_q_weight_1_,
         npu_inst_pe_1_1_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_1_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_1_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_1_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_1_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_1_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_1_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_1_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_1_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_1_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_1_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_1_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_1_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_1_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_1_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_1_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_1_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_1_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_1_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_1_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_1_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_1_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_1_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_1_7_int_q_reg_h_0__1_, npu_inst_pe_1_2_0_n117,
         npu_inst_pe_1_2_0_n116, npu_inst_pe_1_2_0_n115,
         npu_inst_pe_1_2_0_n114, npu_inst_pe_1_2_0_n113,
         npu_inst_pe_1_2_0_n112, npu_inst_pe_1_2_0_n111,
         npu_inst_pe_1_2_0_n110, npu_inst_pe_1_2_0_n109,
         npu_inst_pe_1_2_0_n108, npu_inst_pe_1_2_0_n107,
         npu_inst_pe_1_2_0_n106, npu_inst_pe_1_2_0_n105,
         npu_inst_pe_1_2_0_n104, npu_inst_pe_1_2_0_n103,
         npu_inst_pe_1_2_0_n102, npu_inst_pe_1_2_0_n101,
         npu_inst_pe_1_2_0_n100, npu_inst_pe_1_2_0_n99, npu_inst_pe_1_2_0_n98,
         npu_inst_pe_1_2_0_n36, npu_inst_pe_1_2_0_n35, npu_inst_pe_1_2_0_n34,
         npu_inst_pe_1_2_0_n33, npu_inst_pe_1_2_0_n32, npu_inst_pe_1_2_0_n31,
         npu_inst_pe_1_2_0_n30, npu_inst_pe_1_2_0_n29, npu_inst_pe_1_2_0_n28,
         npu_inst_pe_1_2_0_n25, npu_inst_pe_1_2_0_n24, npu_inst_pe_1_2_0_n23,
         npu_inst_pe_1_2_0_n22, npu_inst_pe_1_2_0_n21, npu_inst_pe_1_2_0_n20,
         npu_inst_pe_1_2_0_n19, npu_inst_pe_1_2_0_n18, npu_inst_pe_1_2_0_n17,
         npu_inst_pe_1_2_0_n16, npu_inst_pe_1_2_0_n15, npu_inst_pe_1_2_0_n14,
         npu_inst_pe_1_2_0_n13, npu_inst_pe_1_2_0_n12, npu_inst_pe_1_2_0_n11,
         npu_inst_pe_1_2_0_n10, npu_inst_pe_1_2_0_n9, npu_inst_pe_1_2_0_n8,
         npu_inst_pe_1_2_0_n7, npu_inst_pe_1_2_0_n6, npu_inst_pe_1_2_0_n5,
         npu_inst_pe_1_2_0_n4, npu_inst_pe_1_2_0_n3, npu_inst_pe_1_2_0_n2,
         npu_inst_pe_1_2_0_n1, npu_inst_pe_1_2_0_sub_77_carry_7_,
         npu_inst_pe_1_2_0_sub_77_carry_6_, npu_inst_pe_1_2_0_sub_77_carry_5_,
         npu_inst_pe_1_2_0_sub_77_carry_4_, npu_inst_pe_1_2_0_sub_77_carry_3_,
         npu_inst_pe_1_2_0_sub_77_carry_2_, npu_inst_pe_1_2_0_sub_77_carry_1_,
         npu_inst_pe_1_2_0_add_79_carry_7_, npu_inst_pe_1_2_0_add_79_carry_6_,
         npu_inst_pe_1_2_0_add_79_carry_5_, npu_inst_pe_1_2_0_add_79_carry_4_,
         npu_inst_pe_1_2_0_add_79_carry_3_, npu_inst_pe_1_2_0_add_79_carry_2_,
         npu_inst_pe_1_2_0_add_79_carry_1_, npu_inst_pe_1_2_0_n97,
         npu_inst_pe_1_2_0_n96, npu_inst_pe_1_2_0_n95, npu_inst_pe_1_2_0_n94,
         npu_inst_pe_1_2_0_n93, npu_inst_pe_1_2_0_n92, npu_inst_pe_1_2_0_n91,
         npu_inst_pe_1_2_0_n90, npu_inst_pe_1_2_0_n89, npu_inst_pe_1_2_0_n88,
         npu_inst_pe_1_2_0_n87, npu_inst_pe_1_2_0_n86, npu_inst_pe_1_2_0_n85,
         npu_inst_pe_1_2_0_n84, npu_inst_pe_1_2_0_n83, npu_inst_pe_1_2_0_n82,
         npu_inst_pe_1_2_0_n81, npu_inst_pe_1_2_0_n80, npu_inst_pe_1_2_0_n79,
         npu_inst_pe_1_2_0_n78, npu_inst_pe_1_2_0_n77, npu_inst_pe_1_2_0_n76,
         npu_inst_pe_1_2_0_n75, npu_inst_pe_1_2_0_n74, npu_inst_pe_1_2_0_n73,
         npu_inst_pe_1_2_0_n72, npu_inst_pe_1_2_0_n71, npu_inst_pe_1_2_0_n70,
         npu_inst_pe_1_2_0_n69, npu_inst_pe_1_2_0_n68, npu_inst_pe_1_2_0_n67,
         npu_inst_pe_1_2_0_n66, npu_inst_pe_1_2_0_n65, npu_inst_pe_1_2_0_n64,
         npu_inst_pe_1_2_0_n63, npu_inst_pe_1_2_0_n62, npu_inst_pe_1_2_0_n61,
         npu_inst_pe_1_2_0_n60, npu_inst_pe_1_2_0_n59, npu_inst_pe_1_2_0_n58,
         npu_inst_pe_1_2_0_n57, npu_inst_pe_1_2_0_n56, npu_inst_pe_1_2_0_n55,
         npu_inst_pe_1_2_0_n54, npu_inst_pe_1_2_0_n53, npu_inst_pe_1_2_0_n52,
         npu_inst_pe_1_2_0_n51, npu_inst_pe_1_2_0_n50, npu_inst_pe_1_2_0_n49,
         npu_inst_pe_1_2_0_n48, npu_inst_pe_1_2_0_n47, npu_inst_pe_1_2_0_n46,
         npu_inst_pe_1_2_0_n45, npu_inst_pe_1_2_0_n44, npu_inst_pe_1_2_0_n43,
         npu_inst_pe_1_2_0_n42, npu_inst_pe_1_2_0_n41, npu_inst_pe_1_2_0_n40,
         npu_inst_pe_1_2_0_n39, npu_inst_pe_1_2_0_n38, npu_inst_pe_1_2_0_n37,
         npu_inst_pe_1_2_0_n27, npu_inst_pe_1_2_0_n26,
         npu_inst_pe_1_2_0_net4116, npu_inst_pe_1_2_0_net4110,
         npu_inst_pe_1_2_0_N94, npu_inst_pe_1_2_0_N93, npu_inst_pe_1_2_0_N84,
         npu_inst_pe_1_2_0_N80, npu_inst_pe_1_2_0_N79, npu_inst_pe_1_2_0_N78,
         npu_inst_pe_1_2_0_N77, npu_inst_pe_1_2_0_N76, npu_inst_pe_1_2_0_N75,
         npu_inst_pe_1_2_0_N74, npu_inst_pe_1_2_0_N73, npu_inst_pe_1_2_0_N72,
         npu_inst_pe_1_2_0_N71, npu_inst_pe_1_2_0_N70, npu_inst_pe_1_2_0_N69,
         npu_inst_pe_1_2_0_N68, npu_inst_pe_1_2_0_N67, npu_inst_pe_1_2_0_N66,
         npu_inst_pe_1_2_0_N65, npu_inst_pe_1_2_0_int_data_0_,
         npu_inst_pe_1_2_0_int_data_1_, npu_inst_pe_1_2_0_int_q_weight_0_,
         npu_inst_pe_1_2_0_int_q_weight_1_,
         npu_inst_pe_1_2_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_0_int_q_reg_h_0__1_, npu_inst_pe_1_2_0_o_data_h_0_,
         npu_inst_pe_1_2_0_o_data_h_1_, npu_inst_pe_1_2_1_n118,
         npu_inst_pe_1_2_1_n117, npu_inst_pe_1_2_1_n116,
         npu_inst_pe_1_2_1_n115, npu_inst_pe_1_2_1_n114,
         npu_inst_pe_1_2_1_n113, npu_inst_pe_1_2_1_n112,
         npu_inst_pe_1_2_1_n111, npu_inst_pe_1_2_1_n110,
         npu_inst_pe_1_2_1_n109, npu_inst_pe_1_2_1_n108,
         npu_inst_pe_1_2_1_n107, npu_inst_pe_1_2_1_n106,
         npu_inst_pe_1_2_1_n105, npu_inst_pe_1_2_1_n104,
         npu_inst_pe_1_2_1_n103, npu_inst_pe_1_2_1_n102,
         npu_inst_pe_1_2_1_n101, npu_inst_pe_1_2_1_n100, npu_inst_pe_1_2_1_n99,
         npu_inst_pe_1_2_1_n98, npu_inst_pe_1_2_1_n36, npu_inst_pe_1_2_1_n35,
         npu_inst_pe_1_2_1_n34, npu_inst_pe_1_2_1_n33, npu_inst_pe_1_2_1_n32,
         npu_inst_pe_1_2_1_n31, npu_inst_pe_1_2_1_n30, npu_inst_pe_1_2_1_n29,
         npu_inst_pe_1_2_1_n28, npu_inst_pe_1_2_1_n25, npu_inst_pe_1_2_1_n24,
         npu_inst_pe_1_2_1_n23, npu_inst_pe_1_2_1_n22, npu_inst_pe_1_2_1_n21,
         npu_inst_pe_1_2_1_n20, npu_inst_pe_1_2_1_n19, npu_inst_pe_1_2_1_n18,
         npu_inst_pe_1_2_1_n17, npu_inst_pe_1_2_1_n16, npu_inst_pe_1_2_1_n15,
         npu_inst_pe_1_2_1_n14, npu_inst_pe_1_2_1_n13, npu_inst_pe_1_2_1_n12,
         npu_inst_pe_1_2_1_n11, npu_inst_pe_1_2_1_n10, npu_inst_pe_1_2_1_n9,
         npu_inst_pe_1_2_1_n8, npu_inst_pe_1_2_1_n7, npu_inst_pe_1_2_1_n6,
         npu_inst_pe_1_2_1_n5, npu_inst_pe_1_2_1_n4, npu_inst_pe_1_2_1_n3,
         npu_inst_pe_1_2_1_n2, npu_inst_pe_1_2_1_n1,
         npu_inst_pe_1_2_1_sub_77_carry_7_, npu_inst_pe_1_2_1_sub_77_carry_6_,
         npu_inst_pe_1_2_1_sub_77_carry_5_, npu_inst_pe_1_2_1_sub_77_carry_4_,
         npu_inst_pe_1_2_1_sub_77_carry_3_, npu_inst_pe_1_2_1_sub_77_carry_2_,
         npu_inst_pe_1_2_1_sub_77_carry_1_, npu_inst_pe_1_2_1_add_79_carry_7_,
         npu_inst_pe_1_2_1_add_79_carry_6_, npu_inst_pe_1_2_1_add_79_carry_5_,
         npu_inst_pe_1_2_1_add_79_carry_4_, npu_inst_pe_1_2_1_add_79_carry_3_,
         npu_inst_pe_1_2_1_add_79_carry_2_, npu_inst_pe_1_2_1_add_79_carry_1_,
         npu_inst_pe_1_2_1_n97, npu_inst_pe_1_2_1_n96, npu_inst_pe_1_2_1_n95,
         npu_inst_pe_1_2_1_n94, npu_inst_pe_1_2_1_n93, npu_inst_pe_1_2_1_n92,
         npu_inst_pe_1_2_1_n91, npu_inst_pe_1_2_1_n90, npu_inst_pe_1_2_1_n89,
         npu_inst_pe_1_2_1_n88, npu_inst_pe_1_2_1_n87, npu_inst_pe_1_2_1_n86,
         npu_inst_pe_1_2_1_n85, npu_inst_pe_1_2_1_n84, npu_inst_pe_1_2_1_n83,
         npu_inst_pe_1_2_1_n82, npu_inst_pe_1_2_1_n81, npu_inst_pe_1_2_1_n80,
         npu_inst_pe_1_2_1_n79, npu_inst_pe_1_2_1_n78, npu_inst_pe_1_2_1_n77,
         npu_inst_pe_1_2_1_n76, npu_inst_pe_1_2_1_n75, npu_inst_pe_1_2_1_n74,
         npu_inst_pe_1_2_1_n73, npu_inst_pe_1_2_1_n72, npu_inst_pe_1_2_1_n71,
         npu_inst_pe_1_2_1_n70, npu_inst_pe_1_2_1_n69, npu_inst_pe_1_2_1_n68,
         npu_inst_pe_1_2_1_n67, npu_inst_pe_1_2_1_n66, npu_inst_pe_1_2_1_n65,
         npu_inst_pe_1_2_1_n64, npu_inst_pe_1_2_1_n63, npu_inst_pe_1_2_1_n62,
         npu_inst_pe_1_2_1_n61, npu_inst_pe_1_2_1_n60, npu_inst_pe_1_2_1_n59,
         npu_inst_pe_1_2_1_n58, npu_inst_pe_1_2_1_n57, npu_inst_pe_1_2_1_n56,
         npu_inst_pe_1_2_1_n55, npu_inst_pe_1_2_1_n54, npu_inst_pe_1_2_1_n53,
         npu_inst_pe_1_2_1_n52, npu_inst_pe_1_2_1_n51, npu_inst_pe_1_2_1_n50,
         npu_inst_pe_1_2_1_n49, npu_inst_pe_1_2_1_n48, npu_inst_pe_1_2_1_n47,
         npu_inst_pe_1_2_1_n46, npu_inst_pe_1_2_1_n45, npu_inst_pe_1_2_1_n44,
         npu_inst_pe_1_2_1_n43, npu_inst_pe_1_2_1_n42, npu_inst_pe_1_2_1_n41,
         npu_inst_pe_1_2_1_n40, npu_inst_pe_1_2_1_n39, npu_inst_pe_1_2_1_n38,
         npu_inst_pe_1_2_1_n37, npu_inst_pe_1_2_1_n27, npu_inst_pe_1_2_1_n26,
         npu_inst_pe_1_2_1_net4093, npu_inst_pe_1_2_1_net4087,
         npu_inst_pe_1_2_1_N94, npu_inst_pe_1_2_1_N93, npu_inst_pe_1_2_1_N84,
         npu_inst_pe_1_2_1_N80, npu_inst_pe_1_2_1_N79, npu_inst_pe_1_2_1_N78,
         npu_inst_pe_1_2_1_N77, npu_inst_pe_1_2_1_N76, npu_inst_pe_1_2_1_N75,
         npu_inst_pe_1_2_1_N74, npu_inst_pe_1_2_1_N73, npu_inst_pe_1_2_1_N72,
         npu_inst_pe_1_2_1_N71, npu_inst_pe_1_2_1_N70, npu_inst_pe_1_2_1_N69,
         npu_inst_pe_1_2_1_N68, npu_inst_pe_1_2_1_N67, npu_inst_pe_1_2_1_N66,
         npu_inst_pe_1_2_1_N65, npu_inst_pe_1_2_1_int_data_0_,
         npu_inst_pe_1_2_1_int_data_1_, npu_inst_pe_1_2_1_int_q_weight_0_,
         npu_inst_pe_1_2_1_int_q_weight_1_,
         npu_inst_pe_1_2_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_1_int_q_reg_h_0__1_, npu_inst_pe_1_2_2_n118,
         npu_inst_pe_1_2_2_n117, npu_inst_pe_1_2_2_n116,
         npu_inst_pe_1_2_2_n115, npu_inst_pe_1_2_2_n114,
         npu_inst_pe_1_2_2_n113, npu_inst_pe_1_2_2_n112,
         npu_inst_pe_1_2_2_n111, npu_inst_pe_1_2_2_n110,
         npu_inst_pe_1_2_2_n109, npu_inst_pe_1_2_2_n108,
         npu_inst_pe_1_2_2_n107, npu_inst_pe_1_2_2_n106,
         npu_inst_pe_1_2_2_n105, npu_inst_pe_1_2_2_n104,
         npu_inst_pe_1_2_2_n103, npu_inst_pe_1_2_2_n102,
         npu_inst_pe_1_2_2_n101, npu_inst_pe_1_2_2_n100, npu_inst_pe_1_2_2_n99,
         npu_inst_pe_1_2_2_n98, npu_inst_pe_1_2_2_n36, npu_inst_pe_1_2_2_n35,
         npu_inst_pe_1_2_2_n34, npu_inst_pe_1_2_2_n33, npu_inst_pe_1_2_2_n32,
         npu_inst_pe_1_2_2_n31, npu_inst_pe_1_2_2_n30, npu_inst_pe_1_2_2_n29,
         npu_inst_pe_1_2_2_n28, npu_inst_pe_1_2_2_n25, npu_inst_pe_1_2_2_n24,
         npu_inst_pe_1_2_2_n23, npu_inst_pe_1_2_2_n22, npu_inst_pe_1_2_2_n21,
         npu_inst_pe_1_2_2_n20, npu_inst_pe_1_2_2_n19, npu_inst_pe_1_2_2_n18,
         npu_inst_pe_1_2_2_n17, npu_inst_pe_1_2_2_n16, npu_inst_pe_1_2_2_n15,
         npu_inst_pe_1_2_2_n14, npu_inst_pe_1_2_2_n13, npu_inst_pe_1_2_2_n12,
         npu_inst_pe_1_2_2_n11, npu_inst_pe_1_2_2_n10, npu_inst_pe_1_2_2_n9,
         npu_inst_pe_1_2_2_n8, npu_inst_pe_1_2_2_n7, npu_inst_pe_1_2_2_n6,
         npu_inst_pe_1_2_2_n5, npu_inst_pe_1_2_2_n4, npu_inst_pe_1_2_2_n3,
         npu_inst_pe_1_2_2_n2, npu_inst_pe_1_2_2_n1,
         npu_inst_pe_1_2_2_sub_77_carry_7_, npu_inst_pe_1_2_2_sub_77_carry_6_,
         npu_inst_pe_1_2_2_sub_77_carry_5_, npu_inst_pe_1_2_2_sub_77_carry_4_,
         npu_inst_pe_1_2_2_sub_77_carry_3_, npu_inst_pe_1_2_2_sub_77_carry_2_,
         npu_inst_pe_1_2_2_sub_77_carry_1_, npu_inst_pe_1_2_2_add_79_carry_7_,
         npu_inst_pe_1_2_2_add_79_carry_6_, npu_inst_pe_1_2_2_add_79_carry_5_,
         npu_inst_pe_1_2_2_add_79_carry_4_, npu_inst_pe_1_2_2_add_79_carry_3_,
         npu_inst_pe_1_2_2_add_79_carry_2_, npu_inst_pe_1_2_2_add_79_carry_1_,
         npu_inst_pe_1_2_2_n97, npu_inst_pe_1_2_2_n96, npu_inst_pe_1_2_2_n95,
         npu_inst_pe_1_2_2_n94, npu_inst_pe_1_2_2_n93, npu_inst_pe_1_2_2_n92,
         npu_inst_pe_1_2_2_n91, npu_inst_pe_1_2_2_n90, npu_inst_pe_1_2_2_n89,
         npu_inst_pe_1_2_2_n88, npu_inst_pe_1_2_2_n87, npu_inst_pe_1_2_2_n86,
         npu_inst_pe_1_2_2_n85, npu_inst_pe_1_2_2_n84, npu_inst_pe_1_2_2_n83,
         npu_inst_pe_1_2_2_n82, npu_inst_pe_1_2_2_n81, npu_inst_pe_1_2_2_n80,
         npu_inst_pe_1_2_2_n79, npu_inst_pe_1_2_2_n78, npu_inst_pe_1_2_2_n77,
         npu_inst_pe_1_2_2_n76, npu_inst_pe_1_2_2_n75, npu_inst_pe_1_2_2_n74,
         npu_inst_pe_1_2_2_n73, npu_inst_pe_1_2_2_n72, npu_inst_pe_1_2_2_n71,
         npu_inst_pe_1_2_2_n70, npu_inst_pe_1_2_2_n69, npu_inst_pe_1_2_2_n68,
         npu_inst_pe_1_2_2_n67, npu_inst_pe_1_2_2_n66, npu_inst_pe_1_2_2_n65,
         npu_inst_pe_1_2_2_n64, npu_inst_pe_1_2_2_n63, npu_inst_pe_1_2_2_n62,
         npu_inst_pe_1_2_2_n61, npu_inst_pe_1_2_2_n60, npu_inst_pe_1_2_2_n59,
         npu_inst_pe_1_2_2_n58, npu_inst_pe_1_2_2_n57, npu_inst_pe_1_2_2_n56,
         npu_inst_pe_1_2_2_n55, npu_inst_pe_1_2_2_n54, npu_inst_pe_1_2_2_n53,
         npu_inst_pe_1_2_2_n52, npu_inst_pe_1_2_2_n51, npu_inst_pe_1_2_2_n50,
         npu_inst_pe_1_2_2_n49, npu_inst_pe_1_2_2_n48, npu_inst_pe_1_2_2_n47,
         npu_inst_pe_1_2_2_n46, npu_inst_pe_1_2_2_n45, npu_inst_pe_1_2_2_n44,
         npu_inst_pe_1_2_2_n43, npu_inst_pe_1_2_2_n42, npu_inst_pe_1_2_2_n41,
         npu_inst_pe_1_2_2_n40, npu_inst_pe_1_2_2_n39, npu_inst_pe_1_2_2_n38,
         npu_inst_pe_1_2_2_n37, npu_inst_pe_1_2_2_n27, npu_inst_pe_1_2_2_n26,
         npu_inst_pe_1_2_2_net4070, npu_inst_pe_1_2_2_net4064,
         npu_inst_pe_1_2_2_N94, npu_inst_pe_1_2_2_N93, npu_inst_pe_1_2_2_N84,
         npu_inst_pe_1_2_2_N80, npu_inst_pe_1_2_2_N79, npu_inst_pe_1_2_2_N78,
         npu_inst_pe_1_2_2_N77, npu_inst_pe_1_2_2_N76, npu_inst_pe_1_2_2_N75,
         npu_inst_pe_1_2_2_N74, npu_inst_pe_1_2_2_N73, npu_inst_pe_1_2_2_N72,
         npu_inst_pe_1_2_2_N71, npu_inst_pe_1_2_2_N70, npu_inst_pe_1_2_2_N69,
         npu_inst_pe_1_2_2_N68, npu_inst_pe_1_2_2_N67, npu_inst_pe_1_2_2_N66,
         npu_inst_pe_1_2_2_N65, npu_inst_pe_1_2_2_int_data_0_,
         npu_inst_pe_1_2_2_int_data_1_, npu_inst_pe_1_2_2_int_q_weight_0_,
         npu_inst_pe_1_2_2_int_q_weight_1_,
         npu_inst_pe_1_2_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_2_int_q_reg_h_0__1_, npu_inst_pe_1_2_3_n118,
         npu_inst_pe_1_2_3_n117, npu_inst_pe_1_2_3_n116,
         npu_inst_pe_1_2_3_n115, npu_inst_pe_1_2_3_n114,
         npu_inst_pe_1_2_3_n113, npu_inst_pe_1_2_3_n112,
         npu_inst_pe_1_2_3_n111, npu_inst_pe_1_2_3_n110,
         npu_inst_pe_1_2_3_n109, npu_inst_pe_1_2_3_n108,
         npu_inst_pe_1_2_3_n107, npu_inst_pe_1_2_3_n106,
         npu_inst_pe_1_2_3_n105, npu_inst_pe_1_2_3_n104,
         npu_inst_pe_1_2_3_n103, npu_inst_pe_1_2_3_n102,
         npu_inst_pe_1_2_3_n101, npu_inst_pe_1_2_3_n100, npu_inst_pe_1_2_3_n99,
         npu_inst_pe_1_2_3_n98, npu_inst_pe_1_2_3_n36, npu_inst_pe_1_2_3_n35,
         npu_inst_pe_1_2_3_n34, npu_inst_pe_1_2_3_n33, npu_inst_pe_1_2_3_n32,
         npu_inst_pe_1_2_3_n31, npu_inst_pe_1_2_3_n30, npu_inst_pe_1_2_3_n29,
         npu_inst_pe_1_2_3_n28, npu_inst_pe_1_2_3_n25, npu_inst_pe_1_2_3_n24,
         npu_inst_pe_1_2_3_n23, npu_inst_pe_1_2_3_n22, npu_inst_pe_1_2_3_n21,
         npu_inst_pe_1_2_3_n20, npu_inst_pe_1_2_3_n19, npu_inst_pe_1_2_3_n18,
         npu_inst_pe_1_2_3_n17, npu_inst_pe_1_2_3_n16, npu_inst_pe_1_2_3_n15,
         npu_inst_pe_1_2_3_n14, npu_inst_pe_1_2_3_n13, npu_inst_pe_1_2_3_n12,
         npu_inst_pe_1_2_3_n11, npu_inst_pe_1_2_3_n10, npu_inst_pe_1_2_3_n9,
         npu_inst_pe_1_2_3_n8, npu_inst_pe_1_2_3_n7, npu_inst_pe_1_2_3_n6,
         npu_inst_pe_1_2_3_n5, npu_inst_pe_1_2_3_n4, npu_inst_pe_1_2_3_n3,
         npu_inst_pe_1_2_3_n2, npu_inst_pe_1_2_3_n1,
         npu_inst_pe_1_2_3_sub_77_carry_7_, npu_inst_pe_1_2_3_sub_77_carry_6_,
         npu_inst_pe_1_2_3_sub_77_carry_5_, npu_inst_pe_1_2_3_sub_77_carry_4_,
         npu_inst_pe_1_2_3_sub_77_carry_3_, npu_inst_pe_1_2_3_sub_77_carry_2_,
         npu_inst_pe_1_2_3_sub_77_carry_1_, npu_inst_pe_1_2_3_add_79_carry_7_,
         npu_inst_pe_1_2_3_add_79_carry_6_, npu_inst_pe_1_2_3_add_79_carry_5_,
         npu_inst_pe_1_2_3_add_79_carry_4_, npu_inst_pe_1_2_3_add_79_carry_3_,
         npu_inst_pe_1_2_3_add_79_carry_2_, npu_inst_pe_1_2_3_add_79_carry_1_,
         npu_inst_pe_1_2_3_n97, npu_inst_pe_1_2_3_n96, npu_inst_pe_1_2_3_n95,
         npu_inst_pe_1_2_3_n94, npu_inst_pe_1_2_3_n93, npu_inst_pe_1_2_3_n92,
         npu_inst_pe_1_2_3_n91, npu_inst_pe_1_2_3_n90, npu_inst_pe_1_2_3_n89,
         npu_inst_pe_1_2_3_n88, npu_inst_pe_1_2_3_n87, npu_inst_pe_1_2_3_n86,
         npu_inst_pe_1_2_3_n85, npu_inst_pe_1_2_3_n84, npu_inst_pe_1_2_3_n83,
         npu_inst_pe_1_2_3_n82, npu_inst_pe_1_2_3_n81, npu_inst_pe_1_2_3_n80,
         npu_inst_pe_1_2_3_n79, npu_inst_pe_1_2_3_n78, npu_inst_pe_1_2_3_n77,
         npu_inst_pe_1_2_3_n76, npu_inst_pe_1_2_3_n75, npu_inst_pe_1_2_3_n74,
         npu_inst_pe_1_2_3_n73, npu_inst_pe_1_2_3_n72, npu_inst_pe_1_2_3_n71,
         npu_inst_pe_1_2_3_n70, npu_inst_pe_1_2_3_n69, npu_inst_pe_1_2_3_n68,
         npu_inst_pe_1_2_3_n67, npu_inst_pe_1_2_3_n66, npu_inst_pe_1_2_3_n65,
         npu_inst_pe_1_2_3_n64, npu_inst_pe_1_2_3_n63, npu_inst_pe_1_2_3_n62,
         npu_inst_pe_1_2_3_n61, npu_inst_pe_1_2_3_n60, npu_inst_pe_1_2_3_n59,
         npu_inst_pe_1_2_3_n58, npu_inst_pe_1_2_3_n57, npu_inst_pe_1_2_3_n56,
         npu_inst_pe_1_2_3_n55, npu_inst_pe_1_2_3_n54, npu_inst_pe_1_2_3_n53,
         npu_inst_pe_1_2_3_n52, npu_inst_pe_1_2_3_n51, npu_inst_pe_1_2_3_n50,
         npu_inst_pe_1_2_3_n49, npu_inst_pe_1_2_3_n48, npu_inst_pe_1_2_3_n47,
         npu_inst_pe_1_2_3_n46, npu_inst_pe_1_2_3_n45, npu_inst_pe_1_2_3_n44,
         npu_inst_pe_1_2_3_n43, npu_inst_pe_1_2_3_n42, npu_inst_pe_1_2_3_n41,
         npu_inst_pe_1_2_3_n40, npu_inst_pe_1_2_3_n39, npu_inst_pe_1_2_3_n38,
         npu_inst_pe_1_2_3_n37, npu_inst_pe_1_2_3_n27, npu_inst_pe_1_2_3_n26,
         npu_inst_pe_1_2_3_net4047, npu_inst_pe_1_2_3_net4041,
         npu_inst_pe_1_2_3_N94, npu_inst_pe_1_2_3_N93, npu_inst_pe_1_2_3_N84,
         npu_inst_pe_1_2_3_N80, npu_inst_pe_1_2_3_N79, npu_inst_pe_1_2_3_N78,
         npu_inst_pe_1_2_3_N77, npu_inst_pe_1_2_3_N76, npu_inst_pe_1_2_3_N75,
         npu_inst_pe_1_2_3_N74, npu_inst_pe_1_2_3_N73, npu_inst_pe_1_2_3_N72,
         npu_inst_pe_1_2_3_N71, npu_inst_pe_1_2_3_N70, npu_inst_pe_1_2_3_N69,
         npu_inst_pe_1_2_3_N68, npu_inst_pe_1_2_3_N67, npu_inst_pe_1_2_3_N66,
         npu_inst_pe_1_2_3_N65, npu_inst_pe_1_2_3_int_data_0_,
         npu_inst_pe_1_2_3_int_data_1_, npu_inst_pe_1_2_3_int_q_weight_0_,
         npu_inst_pe_1_2_3_int_q_weight_1_,
         npu_inst_pe_1_2_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_3_int_q_reg_h_0__1_, npu_inst_pe_1_2_4_n118,
         npu_inst_pe_1_2_4_n117, npu_inst_pe_1_2_4_n116,
         npu_inst_pe_1_2_4_n115, npu_inst_pe_1_2_4_n114,
         npu_inst_pe_1_2_4_n113, npu_inst_pe_1_2_4_n112,
         npu_inst_pe_1_2_4_n111, npu_inst_pe_1_2_4_n110,
         npu_inst_pe_1_2_4_n109, npu_inst_pe_1_2_4_n108,
         npu_inst_pe_1_2_4_n107, npu_inst_pe_1_2_4_n106,
         npu_inst_pe_1_2_4_n105, npu_inst_pe_1_2_4_n104,
         npu_inst_pe_1_2_4_n103, npu_inst_pe_1_2_4_n102,
         npu_inst_pe_1_2_4_n101, npu_inst_pe_1_2_4_n100, npu_inst_pe_1_2_4_n99,
         npu_inst_pe_1_2_4_n98, npu_inst_pe_1_2_4_n36, npu_inst_pe_1_2_4_n35,
         npu_inst_pe_1_2_4_n34, npu_inst_pe_1_2_4_n33, npu_inst_pe_1_2_4_n32,
         npu_inst_pe_1_2_4_n31, npu_inst_pe_1_2_4_n30, npu_inst_pe_1_2_4_n29,
         npu_inst_pe_1_2_4_n28, npu_inst_pe_1_2_4_n25, npu_inst_pe_1_2_4_n24,
         npu_inst_pe_1_2_4_n23, npu_inst_pe_1_2_4_n22, npu_inst_pe_1_2_4_n21,
         npu_inst_pe_1_2_4_n20, npu_inst_pe_1_2_4_n19, npu_inst_pe_1_2_4_n18,
         npu_inst_pe_1_2_4_n17, npu_inst_pe_1_2_4_n16, npu_inst_pe_1_2_4_n15,
         npu_inst_pe_1_2_4_n14, npu_inst_pe_1_2_4_n13, npu_inst_pe_1_2_4_n12,
         npu_inst_pe_1_2_4_n11, npu_inst_pe_1_2_4_n10, npu_inst_pe_1_2_4_n9,
         npu_inst_pe_1_2_4_n8, npu_inst_pe_1_2_4_n7, npu_inst_pe_1_2_4_n6,
         npu_inst_pe_1_2_4_n5, npu_inst_pe_1_2_4_n4, npu_inst_pe_1_2_4_n3,
         npu_inst_pe_1_2_4_n2, npu_inst_pe_1_2_4_n1,
         npu_inst_pe_1_2_4_sub_77_carry_7_, npu_inst_pe_1_2_4_sub_77_carry_6_,
         npu_inst_pe_1_2_4_sub_77_carry_5_, npu_inst_pe_1_2_4_sub_77_carry_4_,
         npu_inst_pe_1_2_4_sub_77_carry_3_, npu_inst_pe_1_2_4_sub_77_carry_2_,
         npu_inst_pe_1_2_4_sub_77_carry_1_, npu_inst_pe_1_2_4_add_79_carry_7_,
         npu_inst_pe_1_2_4_add_79_carry_6_, npu_inst_pe_1_2_4_add_79_carry_5_,
         npu_inst_pe_1_2_4_add_79_carry_4_, npu_inst_pe_1_2_4_add_79_carry_3_,
         npu_inst_pe_1_2_4_add_79_carry_2_, npu_inst_pe_1_2_4_add_79_carry_1_,
         npu_inst_pe_1_2_4_n97, npu_inst_pe_1_2_4_n96, npu_inst_pe_1_2_4_n95,
         npu_inst_pe_1_2_4_n94, npu_inst_pe_1_2_4_n93, npu_inst_pe_1_2_4_n92,
         npu_inst_pe_1_2_4_n91, npu_inst_pe_1_2_4_n90, npu_inst_pe_1_2_4_n89,
         npu_inst_pe_1_2_4_n88, npu_inst_pe_1_2_4_n87, npu_inst_pe_1_2_4_n86,
         npu_inst_pe_1_2_4_n85, npu_inst_pe_1_2_4_n84, npu_inst_pe_1_2_4_n83,
         npu_inst_pe_1_2_4_n82, npu_inst_pe_1_2_4_n81, npu_inst_pe_1_2_4_n80,
         npu_inst_pe_1_2_4_n79, npu_inst_pe_1_2_4_n78, npu_inst_pe_1_2_4_n77,
         npu_inst_pe_1_2_4_n76, npu_inst_pe_1_2_4_n75, npu_inst_pe_1_2_4_n74,
         npu_inst_pe_1_2_4_n73, npu_inst_pe_1_2_4_n72, npu_inst_pe_1_2_4_n71,
         npu_inst_pe_1_2_4_n70, npu_inst_pe_1_2_4_n69, npu_inst_pe_1_2_4_n68,
         npu_inst_pe_1_2_4_n67, npu_inst_pe_1_2_4_n66, npu_inst_pe_1_2_4_n65,
         npu_inst_pe_1_2_4_n64, npu_inst_pe_1_2_4_n63, npu_inst_pe_1_2_4_n62,
         npu_inst_pe_1_2_4_n61, npu_inst_pe_1_2_4_n60, npu_inst_pe_1_2_4_n59,
         npu_inst_pe_1_2_4_n58, npu_inst_pe_1_2_4_n57, npu_inst_pe_1_2_4_n56,
         npu_inst_pe_1_2_4_n55, npu_inst_pe_1_2_4_n54, npu_inst_pe_1_2_4_n53,
         npu_inst_pe_1_2_4_n52, npu_inst_pe_1_2_4_n51, npu_inst_pe_1_2_4_n50,
         npu_inst_pe_1_2_4_n49, npu_inst_pe_1_2_4_n48, npu_inst_pe_1_2_4_n47,
         npu_inst_pe_1_2_4_n46, npu_inst_pe_1_2_4_n45, npu_inst_pe_1_2_4_n44,
         npu_inst_pe_1_2_4_n43, npu_inst_pe_1_2_4_n42, npu_inst_pe_1_2_4_n41,
         npu_inst_pe_1_2_4_n40, npu_inst_pe_1_2_4_n39, npu_inst_pe_1_2_4_n38,
         npu_inst_pe_1_2_4_n37, npu_inst_pe_1_2_4_n27, npu_inst_pe_1_2_4_n26,
         npu_inst_pe_1_2_4_net4024, npu_inst_pe_1_2_4_net4018,
         npu_inst_pe_1_2_4_N94, npu_inst_pe_1_2_4_N93, npu_inst_pe_1_2_4_N84,
         npu_inst_pe_1_2_4_N80, npu_inst_pe_1_2_4_N79, npu_inst_pe_1_2_4_N78,
         npu_inst_pe_1_2_4_N77, npu_inst_pe_1_2_4_N76, npu_inst_pe_1_2_4_N75,
         npu_inst_pe_1_2_4_N74, npu_inst_pe_1_2_4_N73, npu_inst_pe_1_2_4_N72,
         npu_inst_pe_1_2_4_N71, npu_inst_pe_1_2_4_N70, npu_inst_pe_1_2_4_N69,
         npu_inst_pe_1_2_4_N68, npu_inst_pe_1_2_4_N67, npu_inst_pe_1_2_4_N66,
         npu_inst_pe_1_2_4_N65, npu_inst_pe_1_2_4_int_data_0_,
         npu_inst_pe_1_2_4_int_data_1_, npu_inst_pe_1_2_4_int_q_weight_0_,
         npu_inst_pe_1_2_4_int_q_weight_1_,
         npu_inst_pe_1_2_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_4_int_q_reg_h_0__1_, npu_inst_pe_1_2_5_n118,
         npu_inst_pe_1_2_5_n117, npu_inst_pe_1_2_5_n116,
         npu_inst_pe_1_2_5_n115, npu_inst_pe_1_2_5_n114,
         npu_inst_pe_1_2_5_n113, npu_inst_pe_1_2_5_n112,
         npu_inst_pe_1_2_5_n111, npu_inst_pe_1_2_5_n110,
         npu_inst_pe_1_2_5_n109, npu_inst_pe_1_2_5_n108,
         npu_inst_pe_1_2_5_n107, npu_inst_pe_1_2_5_n106,
         npu_inst_pe_1_2_5_n105, npu_inst_pe_1_2_5_n104,
         npu_inst_pe_1_2_5_n103, npu_inst_pe_1_2_5_n102,
         npu_inst_pe_1_2_5_n101, npu_inst_pe_1_2_5_n100, npu_inst_pe_1_2_5_n99,
         npu_inst_pe_1_2_5_n98, npu_inst_pe_1_2_5_n36, npu_inst_pe_1_2_5_n35,
         npu_inst_pe_1_2_5_n34, npu_inst_pe_1_2_5_n33, npu_inst_pe_1_2_5_n32,
         npu_inst_pe_1_2_5_n31, npu_inst_pe_1_2_5_n30, npu_inst_pe_1_2_5_n29,
         npu_inst_pe_1_2_5_n28, npu_inst_pe_1_2_5_n25, npu_inst_pe_1_2_5_n24,
         npu_inst_pe_1_2_5_n23, npu_inst_pe_1_2_5_n22, npu_inst_pe_1_2_5_n21,
         npu_inst_pe_1_2_5_n20, npu_inst_pe_1_2_5_n19, npu_inst_pe_1_2_5_n18,
         npu_inst_pe_1_2_5_n17, npu_inst_pe_1_2_5_n16, npu_inst_pe_1_2_5_n15,
         npu_inst_pe_1_2_5_n14, npu_inst_pe_1_2_5_n13, npu_inst_pe_1_2_5_n12,
         npu_inst_pe_1_2_5_n11, npu_inst_pe_1_2_5_n10, npu_inst_pe_1_2_5_n9,
         npu_inst_pe_1_2_5_n8, npu_inst_pe_1_2_5_n7, npu_inst_pe_1_2_5_n6,
         npu_inst_pe_1_2_5_n5, npu_inst_pe_1_2_5_n4, npu_inst_pe_1_2_5_n3,
         npu_inst_pe_1_2_5_n2, npu_inst_pe_1_2_5_n1,
         npu_inst_pe_1_2_5_sub_77_carry_7_, npu_inst_pe_1_2_5_sub_77_carry_6_,
         npu_inst_pe_1_2_5_sub_77_carry_5_, npu_inst_pe_1_2_5_sub_77_carry_4_,
         npu_inst_pe_1_2_5_sub_77_carry_3_, npu_inst_pe_1_2_5_sub_77_carry_2_,
         npu_inst_pe_1_2_5_sub_77_carry_1_, npu_inst_pe_1_2_5_add_79_carry_7_,
         npu_inst_pe_1_2_5_add_79_carry_6_, npu_inst_pe_1_2_5_add_79_carry_5_,
         npu_inst_pe_1_2_5_add_79_carry_4_, npu_inst_pe_1_2_5_add_79_carry_3_,
         npu_inst_pe_1_2_5_add_79_carry_2_, npu_inst_pe_1_2_5_add_79_carry_1_,
         npu_inst_pe_1_2_5_n97, npu_inst_pe_1_2_5_n96, npu_inst_pe_1_2_5_n95,
         npu_inst_pe_1_2_5_n94, npu_inst_pe_1_2_5_n93, npu_inst_pe_1_2_5_n92,
         npu_inst_pe_1_2_5_n91, npu_inst_pe_1_2_5_n90, npu_inst_pe_1_2_5_n89,
         npu_inst_pe_1_2_5_n88, npu_inst_pe_1_2_5_n87, npu_inst_pe_1_2_5_n86,
         npu_inst_pe_1_2_5_n85, npu_inst_pe_1_2_5_n84, npu_inst_pe_1_2_5_n83,
         npu_inst_pe_1_2_5_n82, npu_inst_pe_1_2_5_n81, npu_inst_pe_1_2_5_n80,
         npu_inst_pe_1_2_5_n79, npu_inst_pe_1_2_5_n78, npu_inst_pe_1_2_5_n77,
         npu_inst_pe_1_2_5_n76, npu_inst_pe_1_2_5_n75, npu_inst_pe_1_2_5_n74,
         npu_inst_pe_1_2_5_n73, npu_inst_pe_1_2_5_n72, npu_inst_pe_1_2_5_n71,
         npu_inst_pe_1_2_5_n70, npu_inst_pe_1_2_5_n69, npu_inst_pe_1_2_5_n68,
         npu_inst_pe_1_2_5_n67, npu_inst_pe_1_2_5_n66, npu_inst_pe_1_2_5_n65,
         npu_inst_pe_1_2_5_n64, npu_inst_pe_1_2_5_n63, npu_inst_pe_1_2_5_n62,
         npu_inst_pe_1_2_5_n61, npu_inst_pe_1_2_5_n60, npu_inst_pe_1_2_5_n59,
         npu_inst_pe_1_2_5_n58, npu_inst_pe_1_2_5_n57, npu_inst_pe_1_2_5_n56,
         npu_inst_pe_1_2_5_n55, npu_inst_pe_1_2_5_n54, npu_inst_pe_1_2_5_n53,
         npu_inst_pe_1_2_5_n52, npu_inst_pe_1_2_5_n51, npu_inst_pe_1_2_5_n50,
         npu_inst_pe_1_2_5_n49, npu_inst_pe_1_2_5_n48, npu_inst_pe_1_2_5_n47,
         npu_inst_pe_1_2_5_n46, npu_inst_pe_1_2_5_n45, npu_inst_pe_1_2_5_n44,
         npu_inst_pe_1_2_5_n43, npu_inst_pe_1_2_5_n42, npu_inst_pe_1_2_5_n41,
         npu_inst_pe_1_2_5_n40, npu_inst_pe_1_2_5_n39, npu_inst_pe_1_2_5_n38,
         npu_inst_pe_1_2_5_n37, npu_inst_pe_1_2_5_n27, npu_inst_pe_1_2_5_n26,
         npu_inst_pe_1_2_5_net4001, npu_inst_pe_1_2_5_net3995,
         npu_inst_pe_1_2_5_N94, npu_inst_pe_1_2_5_N93, npu_inst_pe_1_2_5_N84,
         npu_inst_pe_1_2_5_N80, npu_inst_pe_1_2_5_N79, npu_inst_pe_1_2_5_N78,
         npu_inst_pe_1_2_5_N77, npu_inst_pe_1_2_5_N76, npu_inst_pe_1_2_5_N75,
         npu_inst_pe_1_2_5_N74, npu_inst_pe_1_2_5_N73, npu_inst_pe_1_2_5_N72,
         npu_inst_pe_1_2_5_N71, npu_inst_pe_1_2_5_N70, npu_inst_pe_1_2_5_N69,
         npu_inst_pe_1_2_5_N68, npu_inst_pe_1_2_5_N67, npu_inst_pe_1_2_5_N66,
         npu_inst_pe_1_2_5_N65, npu_inst_pe_1_2_5_int_data_0_,
         npu_inst_pe_1_2_5_int_data_1_, npu_inst_pe_1_2_5_int_q_weight_0_,
         npu_inst_pe_1_2_5_int_q_weight_1_,
         npu_inst_pe_1_2_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_5_int_q_reg_h_0__1_, npu_inst_pe_1_2_6_n118,
         npu_inst_pe_1_2_6_n117, npu_inst_pe_1_2_6_n116,
         npu_inst_pe_1_2_6_n115, npu_inst_pe_1_2_6_n114,
         npu_inst_pe_1_2_6_n113, npu_inst_pe_1_2_6_n112,
         npu_inst_pe_1_2_6_n111, npu_inst_pe_1_2_6_n110,
         npu_inst_pe_1_2_6_n109, npu_inst_pe_1_2_6_n108,
         npu_inst_pe_1_2_6_n107, npu_inst_pe_1_2_6_n106,
         npu_inst_pe_1_2_6_n105, npu_inst_pe_1_2_6_n104,
         npu_inst_pe_1_2_6_n103, npu_inst_pe_1_2_6_n102,
         npu_inst_pe_1_2_6_n101, npu_inst_pe_1_2_6_n100, npu_inst_pe_1_2_6_n99,
         npu_inst_pe_1_2_6_n98, npu_inst_pe_1_2_6_n36, npu_inst_pe_1_2_6_n35,
         npu_inst_pe_1_2_6_n34, npu_inst_pe_1_2_6_n33, npu_inst_pe_1_2_6_n32,
         npu_inst_pe_1_2_6_n31, npu_inst_pe_1_2_6_n30, npu_inst_pe_1_2_6_n29,
         npu_inst_pe_1_2_6_n28, npu_inst_pe_1_2_6_n25, npu_inst_pe_1_2_6_n24,
         npu_inst_pe_1_2_6_n23, npu_inst_pe_1_2_6_n22, npu_inst_pe_1_2_6_n21,
         npu_inst_pe_1_2_6_n20, npu_inst_pe_1_2_6_n19, npu_inst_pe_1_2_6_n18,
         npu_inst_pe_1_2_6_n17, npu_inst_pe_1_2_6_n16, npu_inst_pe_1_2_6_n15,
         npu_inst_pe_1_2_6_n14, npu_inst_pe_1_2_6_n13, npu_inst_pe_1_2_6_n12,
         npu_inst_pe_1_2_6_n11, npu_inst_pe_1_2_6_n10, npu_inst_pe_1_2_6_n9,
         npu_inst_pe_1_2_6_n8, npu_inst_pe_1_2_6_n7, npu_inst_pe_1_2_6_n6,
         npu_inst_pe_1_2_6_n5, npu_inst_pe_1_2_6_n4, npu_inst_pe_1_2_6_n3,
         npu_inst_pe_1_2_6_n2, npu_inst_pe_1_2_6_n1,
         npu_inst_pe_1_2_6_sub_77_carry_7_, npu_inst_pe_1_2_6_sub_77_carry_6_,
         npu_inst_pe_1_2_6_sub_77_carry_5_, npu_inst_pe_1_2_6_sub_77_carry_4_,
         npu_inst_pe_1_2_6_sub_77_carry_3_, npu_inst_pe_1_2_6_sub_77_carry_2_,
         npu_inst_pe_1_2_6_sub_77_carry_1_, npu_inst_pe_1_2_6_add_79_carry_7_,
         npu_inst_pe_1_2_6_add_79_carry_6_, npu_inst_pe_1_2_6_add_79_carry_5_,
         npu_inst_pe_1_2_6_add_79_carry_4_, npu_inst_pe_1_2_6_add_79_carry_3_,
         npu_inst_pe_1_2_6_add_79_carry_2_, npu_inst_pe_1_2_6_add_79_carry_1_,
         npu_inst_pe_1_2_6_n97, npu_inst_pe_1_2_6_n96, npu_inst_pe_1_2_6_n95,
         npu_inst_pe_1_2_6_n94, npu_inst_pe_1_2_6_n93, npu_inst_pe_1_2_6_n92,
         npu_inst_pe_1_2_6_n91, npu_inst_pe_1_2_6_n90, npu_inst_pe_1_2_6_n89,
         npu_inst_pe_1_2_6_n88, npu_inst_pe_1_2_6_n87, npu_inst_pe_1_2_6_n86,
         npu_inst_pe_1_2_6_n85, npu_inst_pe_1_2_6_n84, npu_inst_pe_1_2_6_n83,
         npu_inst_pe_1_2_6_n82, npu_inst_pe_1_2_6_n81, npu_inst_pe_1_2_6_n80,
         npu_inst_pe_1_2_6_n79, npu_inst_pe_1_2_6_n78, npu_inst_pe_1_2_6_n77,
         npu_inst_pe_1_2_6_n76, npu_inst_pe_1_2_6_n75, npu_inst_pe_1_2_6_n74,
         npu_inst_pe_1_2_6_n73, npu_inst_pe_1_2_6_n72, npu_inst_pe_1_2_6_n71,
         npu_inst_pe_1_2_6_n70, npu_inst_pe_1_2_6_n69, npu_inst_pe_1_2_6_n68,
         npu_inst_pe_1_2_6_n67, npu_inst_pe_1_2_6_n66, npu_inst_pe_1_2_6_n65,
         npu_inst_pe_1_2_6_n64, npu_inst_pe_1_2_6_n63, npu_inst_pe_1_2_6_n62,
         npu_inst_pe_1_2_6_n61, npu_inst_pe_1_2_6_n60, npu_inst_pe_1_2_6_n59,
         npu_inst_pe_1_2_6_n58, npu_inst_pe_1_2_6_n57, npu_inst_pe_1_2_6_n56,
         npu_inst_pe_1_2_6_n55, npu_inst_pe_1_2_6_n54, npu_inst_pe_1_2_6_n53,
         npu_inst_pe_1_2_6_n52, npu_inst_pe_1_2_6_n51, npu_inst_pe_1_2_6_n50,
         npu_inst_pe_1_2_6_n49, npu_inst_pe_1_2_6_n48, npu_inst_pe_1_2_6_n47,
         npu_inst_pe_1_2_6_n46, npu_inst_pe_1_2_6_n45, npu_inst_pe_1_2_6_n44,
         npu_inst_pe_1_2_6_n43, npu_inst_pe_1_2_6_n42, npu_inst_pe_1_2_6_n41,
         npu_inst_pe_1_2_6_n40, npu_inst_pe_1_2_6_n39, npu_inst_pe_1_2_6_n38,
         npu_inst_pe_1_2_6_n37, npu_inst_pe_1_2_6_n27, npu_inst_pe_1_2_6_n26,
         npu_inst_pe_1_2_6_net3978, npu_inst_pe_1_2_6_net3972,
         npu_inst_pe_1_2_6_N94, npu_inst_pe_1_2_6_N93, npu_inst_pe_1_2_6_N84,
         npu_inst_pe_1_2_6_N80, npu_inst_pe_1_2_6_N79, npu_inst_pe_1_2_6_N78,
         npu_inst_pe_1_2_6_N77, npu_inst_pe_1_2_6_N76, npu_inst_pe_1_2_6_N75,
         npu_inst_pe_1_2_6_N74, npu_inst_pe_1_2_6_N73, npu_inst_pe_1_2_6_N72,
         npu_inst_pe_1_2_6_N71, npu_inst_pe_1_2_6_N70, npu_inst_pe_1_2_6_N69,
         npu_inst_pe_1_2_6_N68, npu_inst_pe_1_2_6_N67, npu_inst_pe_1_2_6_N66,
         npu_inst_pe_1_2_6_N65, npu_inst_pe_1_2_6_int_data_0_,
         npu_inst_pe_1_2_6_int_data_1_, npu_inst_pe_1_2_6_int_q_weight_0_,
         npu_inst_pe_1_2_6_int_q_weight_1_,
         npu_inst_pe_1_2_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_6_int_q_reg_h_0__1_, npu_inst_pe_1_2_7_n118,
         npu_inst_pe_1_2_7_n117, npu_inst_pe_1_2_7_n116,
         npu_inst_pe_1_2_7_n115, npu_inst_pe_1_2_7_n114,
         npu_inst_pe_1_2_7_n113, npu_inst_pe_1_2_7_n112,
         npu_inst_pe_1_2_7_n111, npu_inst_pe_1_2_7_n110,
         npu_inst_pe_1_2_7_n109, npu_inst_pe_1_2_7_n108,
         npu_inst_pe_1_2_7_n107, npu_inst_pe_1_2_7_n106,
         npu_inst_pe_1_2_7_n105, npu_inst_pe_1_2_7_n104,
         npu_inst_pe_1_2_7_n103, npu_inst_pe_1_2_7_n102,
         npu_inst_pe_1_2_7_n101, npu_inst_pe_1_2_7_n100, npu_inst_pe_1_2_7_n99,
         npu_inst_pe_1_2_7_n98, npu_inst_pe_1_2_7_n36, npu_inst_pe_1_2_7_n35,
         npu_inst_pe_1_2_7_n34, npu_inst_pe_1_2_7_n33, npu_inst_pe_1_2_7_n32,
         npu_inst_pe_1_2_7_n31, npu_inst_pe_1_2_7_n30, npu_inst_pe_1_2_7_n29,
         npu_inst_pe_1_2_7_n28, npu_inst_pe_1_2_7_n25, npu_inst_pe_1_2_7_n24,
         npu_inst_pe_1_2_7_n23, npu_inst_pe_1_2_7_n22, npu_inst_pe_1_2_7_n21,
         npu_inst_pe_1_2_7_n20, npu_inst_pe_1_2_7_n19, npu_inst_pe_1_2_7_n18,
         npu_inst_pe_1_2_7_n17, npu_inst_pe_1_2_7_n16, npu_inst_pe_1_2_7_n15,
         npu_inst_pe_1_2_7_n14, npu_inst_pe_1_2_7_n13, npu_inst_pe_1_2_7_n12,
         npu_inst_pe_1_2_7_n11, npu_inst_pe_1_2_7_n10, npu_inst_pe_1_2_7_n9,
         npu_inst_pe_1_2_7_n8, npu_inst_pe_1_2_7_n7, npu_inst_pe_1_2_7_n6,
         npu_inst_pe_1_2_7_n5, npu_inst_pe_1_2_7_n4, npu_inst_pe_1_2_7_n3,
         npu_inst_pe_1_2_7_n2, npu_inst_pe_1_2_7_n1,
         npu_inst_pe_1_2_7_sub_77_carry_7_, npu_inst_pe_1_2_7_sub_77_carry_6_,
         npu_inst_pe_1_2_7_sub_77_carry_5_, npu_inst_pe_1_2_7_sub_77_carry_4_,
         npu_inst_pe_1_2_7_sub_77_carry_3_, npu_inst_pe_1_2_7_sub_77_carry_2_,
         npu_inst_pe_1_2_7_sub_77_carry_1_, npu_inst_pe_1_2_7_add_79_carry_7_,
         npu_inst_pe_1_2_7_add_79_carry_6_, npu_inst_pe_1_2_7_add_79_carry_5_,
         npu_inst_pe_1_2_7_add_79_carry_4_, npu_inst_pe_1_2_7_add_79_carry_3_,
         npu_inst_pe_1_2_7_add_79_carry_2_, npu_inst_pe_1_2_7_add_79_carry_1_,
         npu_inst_pe_1_2_7_n97, npu_inst_pe_1_2_7_n96, npu_inst_pe_1_2_7_n95,
         npu_inst_pe_1_2_7_n94, npu_inst_pe_1_2_7_n93, npu_inst_pe_1_2_7_n92,
         npu_inst_pe_1_2_7_n91, npu_inst_pe_1_2_7_n90, npu_inst_pe_1_2_7_n89,
         npu_inst_pe_1_2_7_n88, npu_inst_pe_1_2_7_n87, npu_inst_pe_1_2_7_n86,
         npu_inst_pe_1_2_7_n85, npu_inst_pe_1_2_7_n84, npu_inst_pe_1_2_7_n83,
         npu_inst_pe_1_2_7_n82, npu_inst_pe_1_2_7_n81, npu_inst_pe_1_2_7_n80,
         npu_inst_pe_1_2_7_n79, npu_inst_pe_1_2_7_n78, npu_inst_pe_1_2_7_n77,
         npu_inst_pe_1_2_7_n76, npu_inst_pe_1_2_7_n75, npu_inst_pe_1_2_7_n74,
         npu_inst_pe_1_2_7_n73, npu_inst_pe_1_2_7_n72, npu_inst_pe_1_2_7_n71,
         npu_inst_pe_1_2_7_n70, npu_inst_pe_1_2_7_n69, npu_inst_pe_1_2_7_n68,
         npu_inst_pe_1_2_7_n67, npu_inst_pe_1_2_7_n66, npu_inst_pe_1_2_7_n65,
         npu_inst_pe_1_2_7_n64, npu_inst_pe_1_2_7_n63, npu_inst_pe_1_2_7_n62,
         npu_inst_pe_1_2_7_n61, npu_inst_pe_1_2_7_n60, npu_inst_pe_1_2_7_n59,
         npu_inst_pe_1_2_7_n58, npu_inst_pe_1_2_7_n57, npu_inst_pe_1_2_7_n56,
         npu_inst_pe_1_2_7_n55, npu_inst_pe_1_2_7_n54, npu_inst_pe_1_2_7_n53,
         npu_inst_pe_1_2_7_n52, npu_inst_pe_1_2_7_n51, npu_inst_pe_1_2_7_n50,
         npu_inst_pe_1_2_7_n49, npu_inst_pe_1_2_7_n48, npu_inst_pe_1_2_7_n47,
         npu_inst_pe_1_2_7_n46, npu_inst_pe_1_2_7_n45, npu_inst_pe_1_2_7_n44,
         npu_inst_pe_1_2_7_n43, npu_inst_pe_1_2_7_n42, npu_inst_pe_1_2_7_n41,
         npu_inst_pe_1_2_7_n40, npu_inst_pe_1_2_7_n39, npu_inst_pe_1_2_7_n38,
         npu_inst_pe_1_2_7_n37, npu_inst_pe_1_2_7_n27, npu_inst_pe_1_2_7_n26,
         npu_inst_pe_1_2_7_net3955, npu_inst_pe_1_2_7_net3949,
         npu_inst_pe_1_2_7_N94, npu_inst_pe_1_2_7_N93, npu_inst_pe_1_2_7_N84,
         npu_inst_pe_1_2_7_N80, npu_inst_pe_1_2_7_N79, npu_inst_pe_1_2_7_N78,
         npu_inst_pe_1_2_7_N77, npu_inst_pe_1_2_7_N76, npu_inst_pe_1_2_7_N75,
         npu_inst_pe_1_2_7_N74, npu_inst_pe_1_2_7_N73, npu_inst_pe_1_2_7_N72,
         npu_inst_pe_1_2_7_N71, npu_inst_pe_1_2_7_N70, npu_inst_pe_1_2_7_N69,
         npu_inst_pe_1_2_7_N68, npu_inst_pe_1_2_7_N67, npu_inst_pe_1_2_7_N66,
         npu_inst_pe_1_2_7_N65, npu_inst_pe_1_2_7_int_data_0_,
         npu_inst_pe_1_2_7_int_data_1_, npu_inst_pe_1_2_7_int_q_weight_0_,
         npu_inst_pe_1_2_7_int_q_weight_1_,
         npu_inst_pe_1_2_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_2_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_2_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_2_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_2_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_2_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_2_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_2_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_2_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_2_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_2_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_2_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_2_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_2_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_2_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_2_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_2_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_2_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_2_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_2_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_2_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_2_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_2_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_2_7_int_q_reg_h_0__1_, npu_inst_pe_1_3_0_n118,
         npu_inst_pe_1_3_0_n117, npu_inst_pe_1_3_0_n116,
         npu_inst_pe_1_3_0_n115, npu_inst_pe_1_3_0_n114,
         npu_inst_pe_1_3_0_n113, npu_inst_pe_1_3_0_n112,
         npu_inst_pe_1_3_0_n111, npu_inst_pe_1_3_0_n110,
         npu_inst_pe_1_3_0_n109, npu_inst_pe_1_3_0_n108,
         npu_inst_pe_1_3_0_n107, npu_inst_pe_1_3_0_n106,
         npu_inst_pe_1_3_0_n105, npu_inst_pe_1_3_0_n104,
         npu_inst_pe_1_3_0_n103, npu_inst_pe_1_3_0_n102,
         npu_inst_pe_1_3_0_n101, npu_inst_pe_1_3_0_n100, npu_inst_pe_1_3_0_n99,
         npu_inst_pe_1_3_0_n98, npu_inst_pe_1_3_0_n36, npu_inst_pe_1_3_0_n35,
         npu_inst_pe_1_3_0_n34, npu_inst_pe_1_3_0_n33, npu_inst_pe_1_3_0_n32,
         npu_inst_pe_1_3_0_n31, npu_inst_pe_1_3_0_n30, npu_inst_pe_1_3_0_n29,
         npu_inst_pe_1_3_0_n28, npu_inst_pe_1_3_0_n25, npu_inst_pe_1_3_0_n24,
         npu_inst_pe_1_3_0_n23, npu_inst_pe_1_3_0_n22, npu_inst_pe_1_3_0_n21,
         npu_inst_pe_1_3_0_n20, npu_inst_pe_1_3_0_n19, npu_inst_pe_1_3_0_n18,
         npu_inst_pe_1_3_0_n17, npu_inst_pe_1_3_0_n16, npu_inst_pe_1_3_0_n15,
         npu_inst_pe_1_3_0_n14, npu_inst_pe_1_3_0_n13, npu_inst_pe_1_3_0_n12,
         npu_inst_pe_1_3_0_n11, npu_inst_pe_1_3_0_n10, npu_inst_pe_1_3_0_n9,
         npu_inst_pe_1_3_0_n8, npu_inst_pe_1_3_0_n7, npu_inst_pe_1_3_0_n6,
         npu_inst_pe_1_3_0_n5, npu_inst_pe_1_3_0_n4, npu_inst_pe_1_3_0_n3,
         npu_inst_pe_1_3_0_n2, npu_inst_pe_1_3_0_n1,
         npu_inst_pe_1_3_0_sub_77_carry_7_, npu_inst_pe_1_3_0_sub_77_carry_6_,
         npu_inst_pe_1_3_0_sub_77_carry_5_, npu_inst_pe_1_3_0_sub_77_carry_4_,
         npu_inst_pe_1_3_0_sub_77_carry_3_, npu_inst_pe_1_3_0_sub_77_carry_2_,
         npu_inst_pe_1_3_0_sub_77_carry_1_, npu_inst_pe_1_3_0_add_79_carry_7_,
         npu_inst_pe_1_3_0_add_79_carry_6_, npu_inst_pe_1_3_0_add_79_carry_5_,
         npu_inst_pe_1_3_0_add_79_carry_4_, npu_inst_pe_1_3_0_add_79_carry_3_,
         npu_inst_pe_1_3_0_add_79_carry_2_, npu_inst_pe_1_3_0_add_79_carry_1_,
         npu_inst_pe_1_3_0_n97, npu_inst_pe_1_3_0_n96, npu_inst_pe_1_3_0_n95,
         npu_inst_pe_1_3_0_n94, npu_inst_pe_1_3_0_n93, npu_inst_pe_1_3_0_n92,
         npu_inst_pe_1_3_0_n91, npu_inst_pe_1_3_0_n90, npu_inst_pe_1_3_0_n89,
         npu_inst_pe_1_3_0_n88, npu_inst_pe_1_3_0_n87, npu_inst_pe_1_3_0_n86,
         npu_inst_pe_1_3_0_n85, npu_inst_pe_1_3_0_n84, npu_inst_pe_1_3_0_n83,
         npu_inst_pe_1_3_0_n82, npu_inst_pe_1_3_0_n81, npu_inst_pe_1_3_0_n80,
         npu_inst_pe_1_3_0_n79, npu_inst_pe_1_3_0_n78, npu_inst_pe_1_3_0_n77,
         npu_inst_pe_1_3_0_n76, npu_inst_pe_1_3_0_n75, npu_inst_pe_1_3_0_n74,
         npu_inst_pe_1_3_0_n73, npu_inst_pe_1_3_0_n72, npu_inst_pe_1_3_0_n71,
         npu_inst_pe_1_3_0_n70, npu_inst_pe_1_3_0_n69, npu_inst_pe_1_3_0_n68,
         npu_inst_pe_1_3_0_n67, npu_inst_pe_1_3_0_n66, npu_inst_pe_1_3_0_n65,
         npu_inst_pe_1_3_0_n64, npu_inst_pe_1_3_0_n63, npu_inst_pe_1_3_0_n62,
         npu_inst_pe_1_3_0_n61, npu_inst_pe_1_3_0_n60, npu_inst_pe_1_3_0_n59,
         npu_inst_pe_1_3_0_n58, npu_inst_pe_1_3_0_n57, npu_inst_pe_1_3_0_n56,
         npu_inst_pe_1_3_0_n55, npu_inst_pe_1_3_0_n54, npu_inst_pe_1_3_0_n53,
         npu_inst_pe_1_3_0_n52, npu_inst_pe_1_3_0_n51, npu_inst_pe_1_3_0_n50,
         npu_inst_pe_1_3_0_n49, npu_inst_pe_1_3_0_n48, npu_inst_pe_1_3_0_n47,
         npu_inst_pe_1_3_0_n46, npu_inst_pe_1_3_0_n45, npu_inst_pe_1_3_0_n44,
         npu_inst_pe_1_3_0_n43, npu_inst_pe_1_3_0_n42, npu_inst_pe_1_3_0_n41,
         npu_inst_pe_1_3_0_n40, npu_inst_pe_1_3_0_n39, npu_inst_pe_1_3_0_n38,
         npu_inst_pe_1_3_0_n37, npu_inst_pe_1_3_0_n27, npu_inst_pe_1_3_0_n26,
         npu_inst_pe_1_3_0_net3932, npu_inst_pe_1_3_0_net3926,
         npu_inst_pe_1_3_0_N94, npu_inst_pe_1_3_0_N93, npu_inst_pe_1_3_0_N84,
         npu_inst_pe_1_3_0_N80, npu_inst_pe_1_3_0_N79, npu_inst_pe_1_3_0_N78,
         npu_inst_pe_1_3_0_N77, npu_inst_pe_1_3_0_N76, npu_inst_pe_1_3_0_N75,
         npu_inst_pe_1_3_0_N74, npu_inst_pe_1_3_0_N73, npu_inst_pe_1_3_0_N72,
         npu_inst_pe_1_3_0_N71, npu_inst_pe_1_3_0_N70, npu_inst_pe_1_3_0_N69,
         npu_inst_pe_1_3_0_N68, npu_inst_pe_1_3_0_N67, npu_inst_pe_1_3_0_N66,
         npu_inst_pe_1_3_0_N65, npu_inst_pe_1_3_0_int_data_0_,
         npu_inst_pe_1_3_0_int_data_1_, npu_inst_pe_1_3_0_int_q_weight_0_,
         npu_inst_pe_1_3_0_int_q_weight_1_,
         npu_inst_pe_1_3_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_0_int_q_reg_h_0__1_, npu_inst_pe_1_3_0_o_data_h_0_,
         npu_inst_pe_1_3_0_o_data_h_1_, npu_inst_pe_1_3_1_n118,
         npu_inst_pe_1_3_1_n117, npu_inst_pe_1_3_1_n116,
         npu_inst_pe_1_3_1_n115, npu_inst_pe_1_3_1_n114,
         npu_inst_pe_1_3_1_n113, npu_inst_pe_1_3_1_n112,
         npu_inst_pe_1_3_1_n111, npu_inst_pe_1_3_1_n110,
         npu_inst_pe_1_3_1_n109, npu_inst_pe_1_3_1_n108,
         npu_inst_pe_1_3_1_n107, npu_inst_pe_1_3_1_n106,
         npu_inst_pe_1_3_1_n105, npu_inst_pe_1_3_1_n104,
         npu_inst_pe_1_3_1_n103, npu_inst_pe_1_3_1_n102,
         npu_inst_pe_1_3_1_n101, npu_inst_pe_1_3_1_n100, npu_inst_pe_1_3_1_n99,
         npu_inst_pe_1_3_1_n98, npu_inst_pe_1_3_1_n36, npu_inst_pe_1_3_1_n35,
         npu_inst_pe_1_3_1_n34, npu_inst_pe_1_3_1_n33, npu_inst_pe_1_3_1_n32,
         npu_inst_pe_1_3_1_n31, npu_inst_pe_1_3_1_n30, npu_inst_pe_1_3_1_n29,
         npu_inst_pe_1_3_1_n28, npu_inst_pe_1_3_1_n25, npu_inst_pe_1_3_1_n24,
         npu_inst_pe_1_3_1_n23, npu_inst_pe_1_3_1_n22, npu_inst_pe_1_3_1_n21,
         npu_inst_pe_1_3_1_n20, npu_inst_pe_1_3_1_n19, npu_inst_pe_1_3_1_n18,
         npu_inst_pe_1_3_1_n17, npu_inst_pe_1_3_1_n16, npu_inst_pe_1_3_1_n15,
         npu_inst_pe_1_3_1_n14, npu_inst_pe_1_3_1_n13, npu_inst_pe_1_3_1_n12,
         npu_inst_pe_1_3_1_n11, npu_inst_pe_1_3_1_n10, npu_inst_pe_1_3_1_n9,
         npu_inst_pe_1_3_1_n8, npu_inst_pe_1_3_1_n7, npu_inst_pe_1_3_1_n6,
         npu_inst_pe_1_3_1_n5, npu_inst_pe_1_3_1_n4, npu_inst_pe_1_3_1_n3,
         npu_inst_pe_1_3_1_n2, npu_inst_pe_1_3_1_n1,
         npu_inst_pe_1_3_1_sub_77_carry_7_, npu_inst_pe_1_3_1_sub_77_carry_6_,
         npu_inst_pe_1_3_1_sub_77_carry_5_, npu_inst_pe_1_3_1_sub_77_carry_4_,
         npu_inst_pe_1_3_1_sub_77_carry_3_, npu_inst_pe_1_3_1_sub_77_carry_2_,
         npu_inst_pe_1_3_1_sub_77_carry_1_, npu_inst_pe_1_3_1_add_79_carry_7_,
         npu_inst_pe_1_3_1_add_79_carry_6_, npu_inst_pe_1_3_1_add_79_carry_5_,
         npu_inst_pe_1_3_1_add_79_carry_4_, npu_inst_pe_1_3_1_add_79_carry_3_,
         npu_inst_pe_1_3_1_add_79_carry_2_, npu_inst_pe_1_3_1_add_79_carry_1_,
         npu_inst_pe_1_3_1_n97, npu_inst_pe_1_3_1_n96, npu_inst_pe_1_3_1_n95,
         npu_inst_pe_1_3_1_n94, npu_inst_pe_1_3_1_n93, npu_inst_pe_1_3_1_n92,
         npu_inst_pe_1_3_1_n91, npu_inst_pe_1_3_1_n90, npu_inst_pe_1_3_1_n89,
         npu_inst_pe_1_3_1_n88, npu_inst_pe_1_3_1_n87, npu_inst_pe_1_3_1_n86,
         npu_inst_pe_1_3_1_n85, npu_inst_pe_1_3_1_n84, npu_inst_pe_1_3_1_n83,
         npu_inst_pe_1_3_1_n82, npu_inst_pe_1_3_1_n81, npu_inst_pe_1_3_1_n80,
         npu_inst_pe_1_3_1_n79, npu_inst_pe_1_3_1_n78, npu_inst_pe_1_3_1_n77,
         npu_inst_pe_1_3_1_n76, npu_inst_pe_1_3_1_n75, npu_inst_pe_1_3_1_n74,
         npu_inst_pe_1_3_1_n73, npu_inst_pe_1_3_1_n72, npu_inst_pe_1_3_1_n71,
         npu_inst_pe_1_3_1_n70, npu_inst_pe_1_3_1_n69, npu_inst_pe_1_3_1_n68,
         npu_inst_pe_1_3_1_n67, npu_inst_pe_1_3_1_n66, npu_inst_pe_1_3_1_n65,
         npu_inst_pe_1_3_1_n64, npu_inst_pe_1_3_1_n63, npu_inst_pe_1_3_1_n62,
         npu_inst_pe_1_3_1_n61, npu_inst_pe_1_3_1_n60, npu_inst_pe_1_3_1_n59,
         npu_inst_pe_1_3_1_n58, npu_inst_pe_1_3_1_n57, npu_inst_pe_1_3_1_n56,
         npu_inst_pe_1_3_1_n55, npu_inst_pe_1_3_1_n54, npu_inst_pe_1_3_1_n53,
         npu_inst_pe_1_3_1_n52, npu_inst_pe_1_3_1_n51, npu_inst_pe_1_3_1_n50,
         npu_inst_pe_1_3_1_n49, npu_inst_pe_1_3_1_n48, npu_inst_pe_1_3_1_n47,
         npu_inst_pe_1_3_1_n46, npu_inst_pe_1_3_1_n45, npu_inst_pe_1_3_1_n44,
         npu_inst_pe_1_3_1_n43, npu_inst_pe_1_3_1_n42, npu_inst_pe_1_3_1_n41,
         npu_inst_pe_1_3_1_n40, npu_inst_pe_1_3_1_n39, npu_inst_pe_1_3_1_n38,
         npu_inst_pe_1_3_1_n37, npu_inst_pe_1_3_1_n27, npu_inst_pe_1_3_1_n26,
         npu_inst_pe_1_3_1_net3909, npu_inst_pe_1_3_1_net3903,
         npu_inst_pe_1_3_1_N94, npu_inst_pe_1_3_1_N93, npu_inst_pe_1_3_1_N84,
         npu_inst_pe_1_3_1_N80, npu_inst_pe_1_3_1_N79, npu_inst_pe_1_3_1_N78,
         npu_inst_pe_1_3_1_N77, npu_inst_pe_1_3_1_N76, npu_inst_pe_1_3_1_N75,
         npu_inst_pe_1_3_1_N74, npu_inst_pe_1_3_1_N73, npu_inst_pe_1_3_1_N72,
         npu_inst_pe_1_3_1_N71, npu_inst_pe_1_3_1_N70, npu_inst_pe_1_3_1_N69,
         npu_inst_pe_1_3_1_N68, npu_inst_pe_1_3_1_N67, npu_inst_pe_1_3_1_N66,
         npu_inst_pe_1_3_1_N65, npu_inst_pe_1_3_1_int_data_0_,
         npu_inst_pe_1_3_1_int_data_1_, npu_inst_pe_1_3_1_int_q_weight_0_,
         npu_inst_pe_1_3_1_int_q_weight_1_,
         npu_inst_pe_1_3_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_1_int_q_reg_h_0__1_, npu_inst_pe_1_3_2_n118,
         npu_inst_pe_1_3_2_n117, npu_inst_pe_1_3_2_n116,
         npu_inst_pe_1_3_2_n115, npu_inst_pe_1_3_2_n114,
         npu_inst_pe_1_3_2_n113, npu_inst_pe_1_3_2_n112,
         npu_inst_pe_1_3_2_n111, npu_inst_pe_1_3_2_n110,
         npu_inst_pe_1_3_2_n109, npu_inst_pe_1_3_2_n108,
         npu_inst_pe_1_3_2_n107, npu_inst_pe_1_3_2_n106,
         npu_inst_pe_1_3_2_n105, npu_inst_pe_1_3_2_n104,
         npu_inst_pe_1_3_2_n103, npu_inst_pe_1_3_2_n102,
         npu_inst_pe_1_3_2_n101, npu_inst_pe_1_3_2_n100, npu_inst_pe_1_3_2_n99,
         npu_inst_pe_1_3_2_n98, npu_inst_pe_1_3_2_n36, npu_inst_pe_1_3_2_n35,
         npu_inst_pe_1_3_2_n34, npu_inst_pe_1_3_2_n33, npu_inst_pe_1_3_2_n32,
         npu_inst_pe_1_3_2_n31, npu_inst_pe_1_3_2_n30, npu_inst_pe_1_3_2_n29,
         npu_inst_pe_1_3_2_n28, npu_inst_pe_1_3_2_n25, npu_inst_pe_1_3_2_n24,
         npu_inst_pe_1_3_2_n23, npu_inst_pe_1_3_2_n22, npu_inst_pe_1_3_2_n21,
         npu_inst_pe_1_3_2_n20, npu_inst_pe_1_3_2_n19, npu_inst_pe_1_3_2_n18,
         npu_inst_pe_1_3_2_n17, npu_inst_pe_1_3_2_n16, npu_inst_pe_1_3_2_n15,
         npu_inst_pe_1_3_2_n14, npu_inst_pe_1_3_2_n13, npu_inst_pe_1_3_2_n12,
         npu_inst_pe_1_3_2_n11, npu_inst_pe_1_3_2_n10, npu_inst_pe_1_3_2_n9,
         npu_inst_pe_1_3_2_n8, npu_inst_pe_1_3_2_n7, npu_inst_pe_1_3_2_n6,
         npu_inst_pe_1_3_2_n5, npu_inst_pe_1_3_2_n4, npu_inst_pe_1_3_2_n3,
         npu_inst_pe_1_3_2_n2, npu_inst_pe_1_3_2_n1,
         npu_inst_pe_1_3_2_sub_77_carry_7_, npu_inst_pe_1_3_2_sub_77_carry_6_,
         npu_inst_pe_1_3_2_sub_77_carry_5_, npu_inst_pe_1_3_2_sub_77_carry_4_,
         npu_inst_pe_1_3_2_sub_77_carry_3_, npu_inst_pe_1_3_2_sub_77_carry_2_,
         npu_inst_pe_1_3_2_sub_77_carry_1_, npu_inst_pe_1_3_2_add_79_carry_7_,
         npu_inst_pe_1_3_2_add_79_carry_6_, npu_inst_pe_1_3_2_add_79_carry_5_,
         npu_inst_pe_1_3_2_add_79_carry_4_, npu_inst_pe_1_3_2_add_79_carry_3_,
         npu_inst_pe_1_3_2_add_79_carry_2_, npu_inst_pe_1_3_2_add_79_carry_1_,
         npu_inst_pe_1_3_2_n97, npu_inst_pe_1_3_2_n96, npu_inst_pe_1_3_2_n95,
         npu_inst_pe_1_3_2_n94, npu_inst_pe_1_3_2_n93, npu_inst_pe_1_3_2_n92,
         npu_inst_pe_1_3_2_n91, npu_inst_pe_1_3_2_n90, npu_inst_pe_1_3_2_n89,
         npu_inst_pe_1_3_2_n88, npu_inst_pe_1_3_2_n87, npu_inst_pe_1_3_2_n86,
         npu_inst_pe_1_3_2_n85, npu_inst_pe_1_3_2_n84, npu_inst_pe_1_3_2_n83,
         npu_inst_pe_1_3_2_n82, npu_inst_pe_1_3_2_n81, npu_inst_pe_1_3_2_n80,
         npu_inst_pe_1_3_2_n79, npu_inst_pe_1_3_2_n78, npu_inst_pe_1_3_2_n77,
         npu_inst_pe_1_3_2_n76, npu_inst_pe_1_3_2_n75, npu_inst_pe_1_3_2_n74,
         npu_inst_pe_1_3_2_n73, npu_inst_pe_1_3_2_n72, npu_inst_pe_1_3_2_n71,
         npu_inst_pe_1_3_2_n70, npu_inst_pe_1_3_2_n69, npu_inst_pe_1_3_2_n68,
         npu_inst_pe_1_3_2_n67, npu_inst_pe_1_3_2_n66, npu_inst_pe_1_3_2_n65,
         npu_inst_pe_1_3_2_n64, npu_inst_pe_1_3_2_n63, npu_inst_pe_1_3_2_n62,
         npu_inst_pe_1_3_2_n61, npu_inst_pe_1_3_2_n60, npu_inst_pe_1_3_2_n59,
         npu_inst_pe_1_3_2_n58, npu_inst_pe_1_3_2_n57, npu_inst_pe_1_3_2_n56,
         npu_inst_pe_1_3_2_n55, npu_inst_pe_1_3_2_n54, npu_inst_pe_1_3_2_n53,
         npu_inst_pe_1_3_2_n52, npu_inst_pe_1_3_2_n51, npu_inst_pe_1_3_2_n50,
         npu_inst_pe_1_3_2_n49, npu_inst_pe_1_3_2_n48, npu_inst_pe_1_3_2_n47,
         npu_inst_pe_1_3_2_n46, npu_inst_pe_1_3_2_n45, npu_inst_pe_1_3_2_n44,
         npu_inst_pe_1_3_2_n43, npu_inst_pe_1_3_2_n42, npu_inst_pe_1_3_2_n41,
         npu_inst_pe_1_3_2_n40, npu_inst_pe_1_3_2_n39, npu_inst_pe_1_3_2_n38,
         npu_inst_pe_1_3_2_n37, npu_inst_pe_1_3_2_n27, npu_inst_pe_1_3_2_n26,
         npu_inst_pe_1_3_2_net3886, npu_inst_pe_1_3_2_net3880,
         npu_inst_pe_1_3_2_N94, npu_inst_pe_1_3_2_N93, npu_inst_pe_1_3_2_N84,
         npu_inst_pe_1_3_2_N80, npu_inst_pe_1_3_2_N79, npu_inst_pe_1_3_2_N78,
         npu_inst_pe_1_3_2_N77, npu_inst_pe_1_3_2_N76, npu_inst_pe_1_3_2_N75,
         npu_inst_pe_1_3_2_N74, npu_inst_pe_1_3_2_N73, npu_inst_pe_1_3_2_N72,
         npu_inst_pe_1_3_2_N71, npu_inst_pe_1_3_2_N70, npu_inst_pe_1_3_2_N69,
         npu_inst_pe_1_3_2_N68, npu_inst_pe_1_3_2_N67, npu_inst_pe_1_3_2_N66,
         npu_inst_pe_1_3_2_N65, npu_inst_pe_1_3_2_int_data_0_,
         npu_inst_pe_1_3_2_int_data_1_, npu_inst_pe_1_3_2_int_q_weight_0_,
         npu_inst_pe_1_3_2_int_q_weight_1_,
         npu_inst_pe_1_3_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_2_int_q_reg_h_0__1_, npu_inst_pe_1_3_3_n118,
         npu_inst_pe_1_3_3_n117, npu_inst_pe_1_3_3_n116,
         npu_inst_pe_1_3_3_n115, npu_inst_pe_1_3_3_n114,
         npu_inst_pe_1_3_3_n113, npu_inst_pe_1_3_3_n112,
         npu_inst_pe_1_3_3_n111, npu_inst_pe_1_3_3_n110,
         npu_inst_pe_1_3_3_n109, npu_inst_pe_1_3_3_n108,
         npu_inst_pe_1_3_3_n107, npu_inst_pe_1_3_3_n106,
         npu_inst_pe_1_3_3_n105, npu_inst_pe_1_3_3_n104,
         npu_inst_pe_1_3_3_n103, npu_inst_pe_1_3_3_n102,
         npu_inst_pe_1_3_3_n101, npu_inst_pe_1_3_3_n100, npu_inst_pe_1_3_3_n99,
         npu_inst_pe_1_3_3_n98, npu_inst_pe_1_3_3_n36, npu_inst_pe_1_3_3_n35,
         npu_inst_pe_1_3_3_n34, npu_inst_pe_1_3_3_n33, npu_inst_pe_1_3_3_n32,
         npu_inst_pe_1_3_3_n31, npu_inst_pe_1_3_3_n30, npu_inst_pe_1_3_3_n29,
         npu_inst_pe_1_3_3_n28, npu_inst_pe_1_3_3_n25, npu_inst_pe_1_3_3_n24,
         npu_inst_pe_1_3_3_n23, npu_inst_pe_1_3_3_n22, npu_inst_pe_1_3_3_n21,
         npu_inst_pe_1_3_3_n20, npu_inst_pe_1_3_3_n19, npu_inst_pe_1_3_3_n18,
         npu_inst_pe_1_3_3_n17, npu_inst_pe_1_3_3_n16, npu_inst_pe_1_3_3_n15,
         npu_inst_pe_1_3_3_n14, npu_inst_pe_1_3_3_n13, npu_inst_pe_1_3_3_n12,
         npu_inst_pe_1_3_3_n11, npu_inst_pe_1_3_3_n10, npu_inst_pe_1_3_3_n9,
         npu_inst_pe_1_3_3_n8, npu_inst_pe_1_3_3_n7, npu_inst_pe_1_3_3_n6,
         npu_inst_pe_1_3_3_n5, npu_inst_pe_1_3_3_n4, npu_inst_pe_1_3_3_n3,
         npu_inst_pe_1_3_3_n2, npu_inst_pe_1_3_3_n1,
         npu_inst_pe_1_3_3_sub_77_carry_7_, npu_inst_pe_1_3_3_sub_77_carry_6_,
         npu_inst_pe_1_3_3_sub_77_carry_5_, npu_inst_pe_1_3_3_sub_77_carry_4_,
         npu_inst_pe_1_3_3_sub_77_carry_3_, npu_inst_pe_1_3_3_sub_77_carry_2_,
         npu_inst_pe_1_3_3_sub_77_carry_1_, npu_inst_pe_1_3_3_add_79_carry_7_,
         npu_inst_pe_1_3_3_add_79_carry_6_, npu_inst_pe_1_3_3_add_79_carry_5_,
         npu_inst_pe_1_3_3_add_79_carry_4_, npu_inst_pe_1_3_3_add_79_carry_3_,
         npu_inst_pe_1_3_3_add_79_carry_2_, npu_inst_pe_1_3_3_add_79_carry_1_,
         npu_inst_pe_1_3_3_n97, npu_inst_pe_1_3_3_n96, npu_inst_pe_1_3_3_n95,
         npu_inst_pe_1_3_3_n94, npu_inst_pe_1_3_3_n93, npu_inst_pe_1_3_3_n92,
         npu_inst_pe_1_3_3_n91, npu_inst_pe_1_3_3_n90, npu_inst_pe_1_3_3_n89,
         npu_inst_pe_1_3_3_n88, npu_inst_pe_1_3_3_n87, npu_inst_pe_1_3_3_n86,
         npu_inst_pe_1_3_3_n85, npu_inst_pe_1_3_3_n84, npu_inst_pe_1_3_3_n83,
         npu_inst_pe_1_3_3_n82, npu_inst_pe_1_3_3_n81, npu_inst_pe_1_3_3_n80,
         npu_inst_pe_1_3_3_n79, npu_inst_pe_1_3_3_n78, npu_inst_pe_1_3_3_n77,
         npu_inst_pe_1_3_3_n76, npu_inst_pe_1_3_3_n75, npu_inst_pe_1_3_3_n74,
         npu_inst_pe_1_3_3_n73, npu_inst_pe_1_3_3_n72, npu_inst_pe_1_3_3_n71,
         npu_inst_pe_1_3_3_n70, npu_inst_pe_1_3_3_n69, npu_inst_pe_1_3_3_n68,
         npu_inst_pe_1_3_3_n67, npu_inst_pe_1_3_3_n66, npu_inst_pe_1_3_3_n65,
         npu_inst_pe_1_3_3_n64, npu_inst_pe_1_3_3_n63, npu_inst_pe_1_3_3_n62,
         npu_inst_pe_1_3_3_n61, npu_inst_pe_1_3_3_n60, npu_inst_pe_1_3_3_n59,
         npu_inst_pe_1_3_3_n58, npu_inst_pe_1_3_3_n57, npu_inst_pe_1_3_3_n56,
         npu_inst_pe_1_3_3_n55, npu_inst_pe_1_3_3_n54, npu_inst_pe_1_3_3_n53,
         npu_inst_pe_1_3_3_n52, npu_inst_pe_1_3_3_n51, npu_inst_pe_1_3_3_n50,
         npu_inst_pe_1_3_3_n49, npu_inst_pe_1_3_3_n48, npu_inst_pe_1_3_3_n47,
         npu_inst_pe_1_3_3_n46, npu_inst_pe_1_3_3_n45, npu_inst_pe_1_3_3_n44,
         npu_inst_pe_1_3_3_n43, npu_inst_pe_1_3_3_n42, npu_inst_pe_1_3_3_n41,
         npu_inst_pe_1_3_3_n40, npu_inst_pe_1_3_3_n39, npu_inst_pe_1_3_3_n38,
         npu_inst_pe_1_3_3_n37, npu_inst_pe_1_3_3_n27, npu_inst_pe_1_3_3_n26,
         npu_inst_pe_1_3_3_net3863, npu_inst_pe_1_3_3_net3857,
         npu_inst_pe_1_3_3_N94, npu_inst_pe_1_3_3_N93, npu_inst_pe_1_3_3_N84,
         npu_inst_pe_1_3_3_N80, npu_inst_pe_1_3_3_N79, npu_inst_pe_1_3_3_N78,
         npu_inst_pe_1_3_3_N77, npu_inst_pe_1_3_3_N76, npu_inst_pe_1_3_3_N75,
         npu_inst_pe_1_3_3_N74, npu_inst_pe_1_3_3_N73, npu_inst_pe_1_3_3_N72,
         npu_inst_pe_1_3_3_N71, npu_inst_pe_1_3_3_N70, npu_inst_pe_1_3_3_N69,
         npu_inst_pe_1_3_3_N68, npu_inst_pe_1_3_3_N67, npu_inst_pe_1_3_3_N66,
         npu_inst_pe_1_3_3_N65, npu_inst_pe_1_3_3_int_data_0_,
         npu_inst_pe_1_3_3_int_data_1_, npu_inst_pe_1_3_3_int_q_weight_0_,
         npu_inst_pe_1_3_3_int_q_weight_1_,
         npu_inst_pe_1_3_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_3_int_q_reg_h_0__1_, npu_inst_pe_1_3_4_n117,
         npu_inst_pe_1_3_4_n116, npu_inst_pe_1_3_4_n115,
         npu_inst_pe_1_3_4_n114, npu_inst_pe_1_3_4_n113,
         npu_inst_pe_1_3_4_n112, npu_inst_pe_1_3_4_n111,
         npu_inst_pe_1_3_4_n110, npu_inst_pe_1_3_4_n109,
         npu_inst_pe_1_3_4_n108, npu_inst_pe_1_3_4_n107,
         npu_inst_pe_1_3_4_n106, npu_inst_pe_1_3_4_n105,
         npu_inst_pe_1_3_4_n104, npu_inst_pe_1_3_4_n103,
         npu_inst_pe_1_3_4_n102, npu_inst_pe_1_3_4_n101,
         npu_inst_pe_1_3_4_n100, npu_inst_pe_1_3_4_n99, npu_inst_pe_1_3_4_n98,
         npu_inst_pe_1_3_4_n36, npu_inst_pe_1_3_4_n35, npu_inst_pe_1_3_4_n34,
         npu_inst_pe_1_3_4_n33, npu_inst_pe_1_3_4_n32, npu_inst_pe_1_3_4_n31,
         npu_inst_pe_1_3_4_n30, npu_inst_pe_1_3_4_n29, npu_inst_pe_1_3_4_n28,
         npu_inst_pe_1_3_4_n25, npu_inst_pe_1_3_4_n24, npu_inst_pe_1_3_4_n23,
         npu_inst_pe_1_3_4_n22, npu_inst_pe_1_3_4_n21, npu_inst_pe_1_3_4_n20,
         npu_inst_pe_1_3_4_n19, npu_inst_pe_1_3_4_n18, npu_inst_pe_1_3_4_n17,
         npu_inst_pe_1_3_4_n16, npu_inst_pe_1_3_4_n15, npu_inst_pe_1_3_4_n14,
         npu_inst_pe_1_3_4_n13, npu_inst_pe_1_3_4_n12, npu_inst_pe_1_3_4_n11,
         npu_inst_pe_1_3_4_n10, npu_inst_pe_1_3_4_n9, npu_inst_pe_1_3_4_n8,
         npu_inst_pe_1_3_4_n7, npu_inst_pe_1_3_4_n6, npu_inst_pe_1_3_4_n5,
         npu_inst_pe_1_3_4_n4, npu_inst_pe_1_3_4_n3, npu_inst_pe_1_3_4_n2,
         npu_inst_pe_1_3_4_n1, npu_inst_pe_1_3_4_sub_77_carry_7_,
         npu_inst_pe_1_3_4_sub_77_carry_6_, npu_inst_pe_1_3_4_sub_77_carry_5_,
         npu_inst_pe_1_3_4_sub_77_carry_4_, npu_inst_pe_1_3_4_sub_77_carry_3_,
         npu_inst_pe_1_3_4_sub_77_carry_2_, npu_inst_pe_1_3_4_sub_77_carry_1_,
         npu_inst_pe_1_3_4_add_79_carry_7_, npu_inst_pe_1_3_4_add_79_carry_6_,
         npu_inst_pe_1_3_4_add_79_carry_5_, npu_inst_pe_1_3_4_add_79_carry_4_,
         npu_inst_pe_1_3_4_add_79_carry_3_, npu_inst_pe_1_3_4_add_79_carry_2_,
         npu_inst_pe_1_3_4_add_79_carry_1_, npu_inst_pe_1_3_4_n97,
         npu_inst_pe_1_3_4_n96, npu_inst_pe_1_3_4_n95, npu_inst_pe_1_3_4_n94,
         npu_inst_pe_1_3_4_n93, npu_inst_pe_1_3_4_n92, npu_inst_pe_1_3_4_n91,
         npu_inst_pe_1_3_4_n90, npu_inst_pe_1_3_4_n89, npu_inst_pe_1_3_4_n88,
         npu_inst_pe_1_3_4_n87, npu_inst_pe_1_3_4_n86, npu_inst_pe_1_3_4_n85,
         npu_inst_pe_1_3_4_n84, npu_inst_pe_1_3_4_n83, npu_inst_pe_1_3_4_n82,
         npu_inst_pe_1_3_4_n81, npu_inst_pe_1_3_4_n80, npu_inst_pe_1_3_4_n79,
         npu_inst_pe_1_3_4_n78, npu_inst_pe_1_3_4_n77, npu_inst_pe_1_3_4_n76,
         npu_inst_pe_1_3_4_n75, npu_inst_pe_1_3_4_n74, npu_inst_pe_1_3_4_n73,
         npu_inst_pe_1_3_4_n72, npu_inst_pe_1_3_4_n71, npu_inst_pe_1_3_4_n70,
         npu_inst_pe_1_3_4_n69, npu_inst_pe_1_3_4_n68, npu_inst_pe_1_3_4_n67,
         npu_inst_pe_1_3_4_n66, npu_inst_pe_1_3_4_n65, npu_inst_pe_1_3_4_n64,
         npu_inst_pe_1_3_4_n63, npu_inst_pe_1_3_4_n62, npu_inst_pe_1_3_4_n61,
         npu_inst_pe_1_3_4_n60, npu_inst_pe_1_3_4_n59, npu_inst_pe_1_3_4_n58,
         npu_inst_pe_1_3_4_n57, npu_inst_pe_1_3_4_n56, npu_inst_pe_1_3_4_n55,
         npu_inst_pe_1_3_4_n54, npu_inst_pe_1_3_4_n53, npu_inst_pe_1_3_4_n52,
         npu_inst_pe_1_3_4_n51, npu_inst_pe_1_3_4_n50, npu_inst_pe_1_3_4_n49,
         npu_inst_pe_1_3_4_n48, npu_inst_pe_1_3_4_n47, npu_inst_pe_1_3_4_n46,
         npu_inst_pe_1_3_4_n45, npu_inst_pe_1_3_4_n44, npu_inst_pe_1_3_4_n43,
         npu_inst_pe_1_3_4_n42, npu_inst_pe_1_3_4_n41, npu_inst_pe_1_3_4_n40,
         npu_inst_pe_1_3_4_n39, npu_inst_pe_1_3_4_n38, npu_inst_pe_1_3_4_n37,
         npu_inst_pe_1_3_4_n27, npu_inst_pe_1_3_4_n26,
         npu_inst_pe_1_3_4_net3840, npu_inst_pe_1_3_4_net3834,
         npu_inst_pe_1_3_4_N94, npu_inst_pe_1_3_4_N93, npu_inst_pe_1_3_4_N84,
         npu_inst_pe_1_3_4_N80, npu_inst_pe_1_3_4_N79, npu_inst_pe_1_3_4_N78,
         npu_inst_pe_1_3_4_N77, npu_inst_pe_1_3_4_N76, npu_inst_pe_1_3_4_N75,
         npu_inst_pe_1_3_4_N74, npu_inst_pe_1_3_4_N73, npu_inst_pe_1_3_4_N72,
         npu_inst_pe_1_3_4_N71, npu_inst_pe_1_3_4_N70, npu_inst_pe_1_3_4_N69,
         npu_inst_pe_1_3_4_N68, npu_inst_pe_1_3_4_N67, npu_inst_pe_1_3_4_N66,
         npu_inst_pe_1_3_4_N65, npu_inst_pe_1_3_4_int_data_0_,
         npu_inst_pe_1_3_4_int_data_1_, npu_inst_pe_1_3_4_int_q_weight_0_,
         npu_inst_pe_1_3_4_int_q_weight_1_,
         npu_inst_pe_1_3_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_4_int_q_reg_h_0__1_, npu_inst_pe_1_3_5_n118,
         npu_inst_pe_1_3_5_n117, npu_inst_pe_1_3_5_n116,
         npu_inst_pe_1_3_5_n115, npu_inst_pe_1_3_5_n114,
         npu_inst_pe_1_3_5_n113, npu_inst_pe_1_3_5_n112,
         npu_inst_pe_1_3_5_n111, npu_inst_pe_1_3_5_n110,
         npu_inst_pe_1_3_5_n109, npu_inst_pe_1_3_5_n108,
         npu_inst_pe_1_3_5_n107, npu_inst_pe_1_3_5_n106,
         npu_inst_pe_1_3_5_n105, npu_inst_pe_1_3_5_n104,
         npu_inst_pe_1_3_5_n103, npu_inst_pe_1_3_5_n102,
         npu_inst_pe_1_3_5_n101, npu_inst_pe_1_3_5_n100, npu_inst_pe_1_3_5_n99,
         npu_inst_pe_1_3_5_n98, npu_inst_pe_1_3_5_n36, npu_inst_pe_1_3_5_n35,
         npu_inst_pe_1_3_5_n34, npu_inst_pe_1_3_5_n33, npu_inst_pe_1_3_5_n32,
         npu_inst_pe_1_3_5_n31, npu_inst_pe_1_3_5_n30, npu_inst_pe_1_3_5_n29,
         npu_inst_pe_1_3_5_n28, npu_inst_pe_1_3_5_n25, npu_inst_pe_1_3_5_n24,
         npu_inst_pe_1_3_5_n23, npu_inst_pe_1_3_5_n22, npu_inst_pe_1_3_5_n21,
         npu_inst_pe_1_3_5_n20, npu_inst_pe_1_3_5_n19, npu_inst_pe_1_3_5_n18,
         npu_inst_pe_1_3_5_n17, npu_inst_pe_1_3_5_n16, npu_inst_pe_1_3_5_n15,
         npu_inst_pe_1_3_5_n14, npu_inst_pe_1_3_5_n13, npu_inst_pe_1_3_5_n12,
         npu_inst_pe_1_3_5_n11, npu_inst_pe_1_3_5_n10, npu_inst_pe_1_3_5_n9,
         npu_inst_pe_1_3_5_n8, npu_inst_pe_1_3_5_n7, npu_inst_pe_1_3_5_n6,
         npu_inst_pe_1_3_5_n5, npu_inst_pe_1_3_5_n4, npu_inst_pe_1_3_5_n3,
         npu_inst_pe_1_3_5_n2, npu_inst_pe_1_3_5_n1,
         npu_inst_pe_1_3_5_sub_77_carry_7_, npu_inst_pe_1_3_5_sub_77_carry_6_,
         npu_inst_pe_1_3_5_sub_77_carry_5_, npu_inst_pe_1_3_5_sub_77_carry_4_,
         npu_inst_pe_1_3_5_sub_77_carry_3_, npu_inst_pe_1_3_5_sub_77_carry_2_,
         npu_inst_pe_1_3_5_sub_77_carry_1_, npu_inst_pe_1_3_5_add_79_carry_7_,
         npu_inst_pe_1_3_5_add_79_carry_6_, npu_inst_pe_1_3_5_add_79_carry_5_,
         npu_inst_pe_1_3_5_add_79_carry_4_, npu_inst_pe_1_3_5_add_79_carry_3_,
         npu_inst_pe_1_3_5_add_79_carry_2_, npu_inst_pe_1_3_5_add_79_carry_1_,
         npu_inst_pe_1_3_5_n97, npu_inst_pe_1_3_5_n96, npu_inst_pe_1_3_5_n95,
         npu_inst_pe_1_3_5_n94, npu_inst_pe_1_3_5_n93, npu_inst_pe_1_3_5_n92,
         npu_inst_pe_1_3_5_n91, npu_inst_pe_1_3_5_n90, npu_inst_pe_1_3_5_n89,
         npu_inst_pe_1_3_5_n88, npu_inst_pe_1_3_5_n87, npu_inst_pe_1_3_5_n86,
         npu_inst_pe_1_3_5_n85, npu_inst_pe_1_3_5_n84, npu_inst_pe_1_3_5_n83,
         npu_inst_pe_1_3_5_n82, npu_inst_pe_1_3_5_n81, npu_inst_pe_1_3_5_n80,
         npu_inst_pe_1_3_5_n79, npu_inst_pe_1_3_5_n78, npu_inst_pe_1_3_5_n77,
         npu_inst_pe_1_3_5_n76, npu_inst_pe_1_3_5_n75, npu_inst_pe_1_3_5_n74,
         npu_inst_pe_1_3_5_n73, npu_inst_pe_1_3_5_n72, npu_inst_pe_1_3_5_n71,
         npu_inst_pe_1_3_5_n70, npu_inst_pe_1_3_5_n69, npu_inst_pe_1_3_5_n68,
         npu_inst_pe_1_3_5_n67, npu_inst_pe_1_3_5_n66, npu_inst_pe_1_3_5_n65,
         npu_inst_pe_1_3_5_n64, npu_inst_pe_1_3_5_n63, npu_inst_pe_1_3_5_n62,
         npu_inst_pe_1_3_5_n61, npu_inst_pe_1_3_5_n60, npu_inst_pe_1_3_5_n59,
         npu_inst_pe_1_3_5_n58, npu_inst_pe_1_3_5_n57, npu_inst_pe_1_3_5_n56,
         npu_inst_pe_1_3_5_n55, npu_inst_pe_1_3_5_n54, npu_inst_pe_1_3_5_n53,
         npu_inst_pe_1_3_5_n52, npu_inst_pe_1_3_5_n51, npu_inst_pe_1_3_5_n50,
         npu_inst_pe_1_3_5_n49, npu_inst_pe_1_3_5_n48, npu_inst_pe_1_3_5_n47,
         npu_inst_pe_1_3_5_n46, npu_inst_pe_1_3_5_n45, npu_inst_pe_1_3_5_n44,
         npu_inst_pe_1_3_5_n43, npu_inst_pe_1_3_5_n42, npu_inst_pe_1_3_5_n41,
         npu_inst_pe_1_3_5_n40, npu_inst_pe_1_3_5_n39, npu_inst_pe_1_3_5_n38,
         npu_inst_pe_1_3_5_n37, npu_inst_pe_1_3_5_n27, npu_inst_pe_1_3_5_n26,
         npu_inst_pe_1_3_5_net3817, npu_inst_pe_1_3_5_net3811,
         npu_inst_pe_1_3_5_N94, npu_inst_pe_1_3_5_N93, npu_inst_pe_1_3_5_N84,
         npu_inst_pe_1_3_5_N80, npu_inst_pe_1_3_5_N79, npu_inst_pe_1_3_5_N78,
         npu_inst_pe_1_3_5_N77, npu_inst_pe_1_3_5_N76, npu_inst_pe_1_3_5_N75,
         npu_inst_pe_1_3_5_N74, npu_inst_pe_1_3_5_N73, npu_inst_pe_1_3_5_N72,
         npu_inst_pe_1_3_5_N71, npu_inst_pe_1_3_5_N70, npu_inst_pe_1_3_5_N69,
         npu_inst_pe_1_3_5_N68, npu_inst_pe_1_3_5_N67, npu_inst_pe_1_3_5_N66,
         npu_inst_pe_1_3_5_N65, npu_inst_pe_1_3_5_int_data_0_,
         npu_inst_pe_1_3_5_int_data_1_, npu_inst_pe_1_3_5_int_q_weight_0_,
         npu_inst_pe_1_3_5_int_q_weight_1_,
         npu_inst_pe_1_3_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_5_int_q_reg_h_0__1_, npu_inst_pe_1_3_6_n118,
         npu_inst_pe_1_3_6_n117, npu_inst_pe_1_3_6_n116,
         npu_inst_pe_1_3_6_n115, npu_inst_pe_1_3_6_n114,
         npu_inst_pe_1_3_6_n113, npu_inst_pe_1_3_6_n112,
         npu_inst_pe_1_3_6_n111, npu_inst_pe_1_3_6_n110,
         npu_inst_pe_1_3_6_n109, npu_inst_pe_1_3_6_n108,
         npu_inst_pe_1_3_6_n107, npu_inst_pe_1_3_6_n106,
         npu_inst_pe_1_3_6_n105, npu_inst_pe_1_3_6_n104,
         npu_inst_pe_1_3_6_n103, npu_inst_pe_1_3_6_n102,
         npu_inst_pe_1_3_6_n101, npu_inst_pe_1_3_6_n100, npu_inst_pe_1_3_6_n99,
         npu_inst_pe_1_3_6_n98, npu_inst_pe_1_3_6_n36, npu_inst_pe_1_3_6_n35,
         npu_inst_pe_1_3_6_n34, npu_inst_pe_1_3_6_n33, npu_inst_pe_1_3_6_n32,
         npu_inst_pe_1_3_6_n31, npu_inst_pe_1_3_6_n30, npu_inst_pe_1_3_6_n29,
         npu_inst_pe_1_3_6_n28, npu_inst_pe_1_3_6_n25, npu_inst_pe_1_3_6_n24,
         npu_inst_pe_1_3_6_n23, npu_inst_pe_1_3_6_n22, npu_inst_pe_1_3_6_n21,
         npu_inst_pe_1_3_6_n20, npu_inst_pe_1_3_6_n19, npu_inst_pe_1_3_6_n18,
         npu_inst_pe_1_3_6_n17, npu_inst_pe_1_3_6_n16, npu_inst_pe_1_3_6_n15,
         npu_inst_pe_1_3_6_n14, npu_inst_pe_1_3_6_n13, npu_inst_pe_1_3_6_n12,
         npu_inst_pe_1_3_6_n11, npu_inst_pe_1_3_6_n10, npu_inst_pe_1_3_6_n9,
         npu_inst_pe_1_3_6_n8, npu_inst_pe_1_3_6_n7, npu_inst_pe_1_3_6_n6,
         npu_inst_pe_1_3_6_n5, npu_inst_pe_1_3_6_n4, npu_inst_pe_1_3_6_n3,
         npu_inst_pe_1_3_6_n2, npu_inst_pe_1_3_6_n1,
         npu_inst_pe_1_3_6_sub_77_carry_7_, npu_inst_pe_1_3_6_sub_77_carry_6_,
         npu_inst_pe_1_3_6_sub_77_carry_5_, npu_inst_pe_1_3_6_sub_77_carry_4_,
         npu_inst_pe_1_3_6_sub_77_carry_3_, npu_inst_pe_1_3_6_sub_77_carry_2_,
         npu_inst_pe_1_3_6_sub_77_carry_1_, npu_inst_pe_1_3_6_add_79_carry_7_,
         npu_inst_pe_1_3_6_add_79_carry_6_, npu_inst_pe_1_3_6_add_79_carry_5_,
         npu_inst_pe_1_3_6_add_79_carry_4_, npu_inst_pe_1_3_6_add_79_carry_3_,
         npu_inst_pe_1_3_6_add_79_carry_2_, npu_inst_pe_1_3_6_add_79_carry_1_,
         npu_inst_pe_1_3_6_n97, npu_inst_pe_1_3_6_n96, npu_inst_pe_1_3_6_n95,
         npu_inst_pe_1_3_6_n94, npu_inst_pe_1_3_6_n93, npu_inst_pe_1_3_6_n92,
         npu_inst_pe_1_3_6_n91, npu_inst_pe_1_3_6_n90, npu_inst_pe_1_3_6_n89,
         npu_inst_pe_1_3_6_n88, npu_inst_pe_1_3_6_n87, npu_inst_pe_1_3_6_n86,
         npu_inst_pe_1_3_6_n85, npu_inst_pe_1_3_6_n84, npu_inst_pe_1_3_6_n83,
         npu_inst_pe_1_3_6_n82, npu_inst_pe_1_3_6_n81, npu_inst_pe_1_3_6_n80,
         npu_inst_pe_1_3_6_n79, npu_inst_pe_1_3_6_n78, npu_inst_pe_1_3_6_n77,
         npu_inst_pe_1_3_6_n76, npu_inst_pe_1_3_6_n75, npu_inst_pe_1_3_6_n74,
         npu_inst_pe_1_3_6_n73, npu_inst_pe_1_3_6_n72, npu_inst_pe_1_3_6_n71,
         npu_inst_pe_1_3_6_n70, npu_inst_pe_1_3_6_n69, npu_inst_pe_1_3_6_n68,
         npu_inst_pe_1_3_6_n67, npu_inst_pe_1_3_6_n66, npu_inst_pe_1_3_6_n65,
         npu_inst_pe_1_3_6_n64, npu_inst_pe_1_3_6_n63, npu_inst_pe_1_3_6_n62,
         npu_inst_pe_1_3_6_n61, npu_inst_pe_1_3_6_n60, npu_inst_pe_1_3_6_n59,
         npu_inst_pe_1_3_6_n58, npu_inst_pe_1_3_6_n57, npu_inst_pe_1_3_6_n56,
         npu_inst_pe_1_3_6_n55, npu_inst_pe_1_3_6_n54, npu_inst_pe_1_3_6_n53,
         npu_inst_pe_1_3_6_n52, npu_inst_pe_1_3_6_n51, npu_inst_pe_1_3_6_n50,
         npu_inst_pe_1_3_6_n49, npu_inst_pe_1_3_6_n48, npu_inst_pe_1_3_6_n47,
         npu_inst_pe_1_3_6_n46, npu_inst_pe_1_3_6_n45, npu_inst_pe_1_3_6_n44,
         npu_inst_pe_1_3_6_n43, npu_inst_pe_1_3_6_n42, npu_inst_pe_1_3_6_n41,
         npu_inst_pe_1_3_6_n40, npu_inst_pe_1_3_6_n39, npu_inst_pe_1_3_6_n38,
         npu_inst_pe_1_3_6_n37, npu_inst_pe_1_3_6_n27, npu_inst_pe_1_3_6_n26,
         npu_inst_pe_1_3_6_net3794, npu_inst_pe_1_3_6_net3788,
         npu_inst_pe_1_3_6_N94, npu_inst_pe_1_3_6_N93, npu_inst_pe_1_3_6_N84,
         npu_inst_pe_1_3_6_N80, npu_inst_pe_1_3_6_N79, npu_inst_pe_1_3_6_N78,
         npu_inst_pe_1_3_6_N77, npu_inst_pe_1_3_6_N76, npu_inst_pe_1_3_6_N75,
         npu_inst_pe_1_3_6_N74, npu_inst_pe_1_3_6_N73, npu_inst_pe_1_3_6_N72,
         npu_inst_pe_1_3_6_N71, npu_inst_pe_1_3_6_N70, npu_inst_pe_1_3_6_N69,
         npu_inst_pe_1_3_6_N68, npu_inst_pe_1_3_6_N67, npu_inst_pe_1_3_6_N66,
         npu_inst_pe_1_3_6_N65, npu_inst_pe_1_3_6_int_data_0_,
         npu_inst_pe_1_3_6_int_data_1_, npu_inst_pe_1_3_6_int_q_weight_0_,
         npu_inst_pe_1_3_6_int_q_weight_1_,
         npu_inst_pe_1_3_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_6_int_q_reg_h_0__1_, npu_inst_pe_1_3_7_n118,
         npu_inst_pe_1_3_7_n117, npu_inst_pe_1_3_7_n116,
         npu_inst_pe_1_3_7_n115, npu_inst_pe_1_3_7_n114,
         npu_inst_pe_1_3_7_n113, npu_inst_pe_1_3_7_n112,
         npu_inst_pe_1_3_7_n111, npu_inst_pe_1_3_7_n110,
         npu_inst_pe_1_3_7_n109, npu_inst_pe_1_3_7_n108,
         npu_inst_pe_1_3_7_n107, npu_inst_pe_1_3_7_n106,
         npu_inst_pe_1_3_7_n105, npu_inst_pe_1_3_7_n104,
         npu_inst_pe_1_3_7_n103, npu_inst_pe_1_3_7_n102,
         npu_inst_pe_1_3_7_n101, npu_inst_pe_1_3_7_n100, npu_inst_pe_1_3_7_n99,
         npu_inst_pe_1_3_7_n98, npu_inst_pe_1_3_7_n36, npu_inst_pe_1_3_7_n35,
         npu_inst_pe_1_3_7_n34, npu_inst_pe_1_3_7_n33, npu_inst_pe_1_3_7_n32,
         npu_inst_pe_1_3_7_n31, npu_inst_pe_1_3_7_n30, npu_inst_pe_1_3_7_n29,
         npu_inst_pe_1_3_7_n28, npu_inst_pe_1_3_7_n25, npu_inst_pe_1_3_7_n24,
         npu_inst_pe_1_3_7_n23, npu_inst_pe_1_3_7_n22, npu_inst_pe_1_3_7_n21,
         npu_inst_pe_1_3_7_n20, npu_inst_pe_1_3_7_n19, npu_inst_pe_1_3_7_n18,
         npu_inst_pe_1_3_7_n17, npu_inst_pe_1_3_7_n16, npu_inst_pe_1_3_7_n15,
         npu_inst_pe_1_3_7_n14, npu_inst_pe_1_3_7_n13, npu_inst_pe_1_3_7_n12,
         npu_inst_pe_1_3_7_n11, npu_inst_pe_1_3_7_n10, npu_inst_pe_1_3_7_n9,
         npu_inst_pe_1_3_7_n8, npu_inst_pe_1_3_7_n7, npu_inst_pe_1_3_7_n6,
         npu_inst_pe_1_3_7_n5, npu_inst_pe_1_3_7_n4, npu_inst_pe_1_3_7_n3,
         npu_inst_pe_1_3_7_n2, npu_inst_pe_1_3_7_n1,
         npu_inst_pe_1_3_7_sub_77_carry_7_, npu_inst_pe_1_3_7_sub_77_carry_6_,
         npu_inst_pe_1_3_7_sub_77_carry_5_, npu_inst_pe_1_3_7_sub_77_carry_4_,
         npu_inst_pe_1_3_7_sub_77_carry_3_, npu_inst_pe_1_3_7_sub_77_carry_2_,
         npu_inst_pe_1_3_7_sub_77_carry_1_, npu_inst_pe_1_3_7_add_79_carry_7_,
         npu_inst_pe_1_3_7_add_79_carry_6_, npu_inst_pe_1_3_7_add_79_carry_5_,
         npu_inst_pe_1_3_7_add_79_carry_4_, npu_inst_pe_1_3_7_add_79_carry_3_,
         npu_inst_pe_1_3_7_add_79_carry_2_, npu_inst_pe_1_3_7_add_79_carry_1_,
         npu_inst_pe_1_3_7_n97, npu_inst_pe_1_3_7_n96, npu_inst_pe_1_3_7_n95,
         npu_inst_pe_1_3_7_n94, npu_inst_pe_1_3_7_n93, npu_inst_pe_1_3_7_n92,
         npu_inst_pe_1_3_7_n91, npu_inst_pe_1_3_7_n90, npu_inst_pe_1_3_7_n89,
         npu_inst_pe_1_3_7_n88, npu_inst_pe_1_3_7_n87, npu_inst_pe_1_3_7_n86,
         npu_inst_pe_1_3_7_n85, npu_inst_pe_1_3_7_n84, npu_inst_pe_1_3_7_n83,
         npu_inst_pe_1_3_7_n82, npu_inst_pe_1_3_7_n81, npu_inst_pe_1_3_7_n80,
         npu_inst_pe_1_3_7_n79, npu_inst_pe_1_3_7_n78, npu_inst_pe_1_3_7_n77,
         npu_inst_pe_1_3_7_n76, npu_inst_pe_1_3_7_n75, npu_inst_pe_1_3_7_n74,
         npu_inst_pe_1_3_7_n73, npu_inst_pe_1_3_7_n72, npu_inst_pe_1_3_7_n71,
         npu_inst_pe_1_3_7_n70, npu_inst_pe_1_3_7_n69, npu_inst_pe_1_3_7_n68,
         npu_inst_pe_1_3_7_n67, npu_inst_pe_1_3_7_n66, npu_inst_pe_1_3_7_n65,
         npu_inst_pe_1_3_7_n64, npu_inst_pe_1_3_7_n63, npu_inst_pe_1_3_7_n62,
         npu_inst_pe_1_3_7_n61, npu_inst_pe_1_3_7_n60, npu_inst_pe_1_3_7_n59,
         npu_inst_pe_1_3_7_n58, npu_inst_pe_1_3_7_n57, npu_inst_pe_1_3_7_n56,
         npu_inst_pe_1_3_7_n55, npu_inst_pe_1_3_7_n54, npu_inst_pe_1_3_7_n53,
         npu_inst_pe_1_3_7_n52, npu_inst_pe_1_3_7_n51, npu_inst_pe_1_3_7_n50,
         npu_inst_pe_1_3_7_n49, npu_inst_pe_1_3_7_n48, npu_inst_pe_1_3_7_n47,
         npu_inst_pe_1_3_7_n46, npu_inst_pe_1_3_7_n45, npu_inst_pe_1_3_7_n44,
         npu_inst_pe_1_3_7_n43, npu_inst_pe_1_3_7_n42, npu_inst_pe_1_3_7_n41,
         npu_inst_pe_1_3_7_n40, npu_inst_pe_1_3_7_n39, npu_inst_pe_1_3_7_n38,
         npu_inst_pe_1_3_7_n37, npu_inst_pe_1_3_7_n27, npu_inst_pe_1_3_7_n26,
         npu_inst_pe_1_3_7_net3771, npu_inst_pe_1_3_7_net3765,
         npu_inst_pe_1_3_7_N94, npu_inst_pe_1_3_7_N93, npu_inst_pe_1_3_7_N84,
         npu_inst_pe_1_3_7_N80, npu_inst_pe_1_3_7_N79, npu_inst_pe_1_3_7_N78,
         npu_inst_pe_1_3_7_N77, npu_inst_pe_1_3_7_N76, npu_inst_pe_1_3_7_N75,
         npu_inst_pe_1_3_7_N74, npu_inst_pe_1_3_7_N73, npu_inst_pe_1_3_7_N72,
         npu_inst_pe_1_3_7_N71, npu_inst_pe_1_3_7_N70, npu_inst_pe_1_3_7_N69,
         npu_inst_pe_1_3_7_N68, npu_inst_pe_1_3_7_N67, npu_inst_pe_1_3_7_N66,
         npu_inst_pe_1_3_7_N65, npu_inst_pe_1_3_7_int_data_0_,
         npu_inst_pe_1_3_7_int_data_1_, npu_inst_pe_1_3_7_int_q_weight_0_,
         npu_inst_pe_1_3_7_int_q_weight_1_,
         npu_inst_pe_1_3_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_3_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_3_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_3_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_3_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_3_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_3_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_3_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_3_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_3_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_3_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_3_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_3_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_3_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_3_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_3_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_3_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_3_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_3_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_3_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_3_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_3_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_3_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_3_7_int_q_reg_h_0__1_, npu_inst_pe_1_4_0_n118,
         npu_inst_pe_1_4_0_n117, npu_inst_pe_1_4_0_n116,
         npu_inst_pe_1_4_0_n115, npu_inst_pe_1_4_0_n114,
         npu_inst_pe_1_4_0_n113, npu_inst_pe_1_4_0_n112,
         npu_inst_pe_1_4_0_n111, npu_inst_pe_1_4_0_n110,
         npu_inst_pe_1_4_0_n109, npu_inst_pe_1_4_0_n108,
         npu_inst_pe_1_4_0_n107, npu_inst_pe_1_4_0_n106,
         npu_inst_pe_1_4_0_n105, npu_inst_pe_1_4_0_n104,
         npu_inst_pe_1_4_0_n103, npu_inst_pe_1_4_0_n102,
         npu_inst_pe_1_4_0_n101, npu_inst_pe_1_4_0_n100, npu_inst_pe_1_4_0_n99,
         npu_inst_pe_1_4_0_n98, npu_inst_pe_1_4_0_n36, npu_inst_pe_1_4_0_n35,
         npu_inst_pe_1_4_0_n34, npu_inst_pe_1_4_0_n33, npu_inst_pe_1_4_0_n32,
         npu_inst_pe_1_4_0_n31, npu_inst_pe_1_4_0_n30, npu_inst_pe_1_4_0_n29,
         npu_inst_pe_1_4_0_n28, npu_inst_pe_1_4_0_n25, npu_inst_pe_1_4_0_n24,
         npu_inst_pe_1_4_0_n23, npu_inst_pe_1_4_0_n22, npu_inst_pe_1_4_0_n21,
         npu_inst_pe_1_4_0_n20, npu_inst_pe_1_4_0_n19, npu_inst_pe_1_4_0_n18,
         npu_inst_pe_1_4_0_n17, npu_inst_pe_1_4_0_n16, npu_inst_pe_1_4_0_n15,
         npu_inst_pe_1_4_0_n14, npu_inst_pe_1_4_0_n13, npu_inst_pe_1_4_0_n12,
         npu_inst_pe_1_4_0_n11, npu_inst_pe_1_4_0_n10, npu_inst_pe_1_4_0_n9,
         npu_inst_pe_1_4_0_n8, npu_inst_pe_1_4_0_n7, npu_inst_pe_1_4_0_n6,
         npu_inst_pe_1_4_0_n5, npu_inst_pe_1_4_0_n4, npu_inst_pe_1_4_0_n3,
         npu_inst_pe_1_4_0_n2, npu_inst_pe_1_4_0_n1,
         npu_inst_pe_1_4_0_sub_77_carry_7_, npu_inst_pe_1_4_0_sub_77_carry_6_,
         npu_inst_pe_1_4_0_sub_77_carry_5_, npu_inst_pe_1_4_0_sub_77_carry_4_,
         npu_inst_pe_1_4_0_sub_77_carry_3_, npu_inst_pe_1_4_0_sub_77_carry_2_,
         npu_inst_pe_1_4_0_sub_77_carry_1_, npu_inst_pe_1_4_0_add_79_carry_7_,
         npu_inst_pe_1_4_0_add_79_carry_6_, npu_inst_pe_1_4_0_add_79_carry_5_,
         npu_inst_pe_1_4_0_add_79_carry_4_, npu_inst_pe_1_4_0_add_79_carry_3_,
         npu_inst_pe_1_4_0_add_79_carry_2_, npu_inst_pe_1_4_0_add_79_carry_1_,
         npu_inst_pe_1_4_0_n97, npu_inst_pe_1_4_0_n96, npu_inst_pe_1_4_0_n95,
         npu_inst_pe_1_4_0_n94, npu_inst_pe_1_4_0_n93, npu_inst_pe_1_4_0_n92,
         npu_inst_pe_1_4_0_n91, npu_inst_pe_1_4_0_n90, npu_inst_pe_1_4_0_n89,
         npu_inst_pe_1_4_0_n88, npu_inst_pe_1_4_0_n87, npu_inst_pe_1_4_0_n86,
         npu_inst_pe_1_4_0_n85, npu_inst_pe_1_4_0_n84, npu_inst_pe_1_4_0_n83,
         npu_inst_pe_1_4_0_n82, npu_inst_pe_1_4_0_n81, npu_inst_pe_1_4_0_n80,
         npu_inst_pe_1_4_0_n79, npu_inst_pe_1_4_0_n78, npu_inst_pe_1_4_0_n77,
         npu_inst_pe_1_4_0_n76, npu_inst_pe_1_4_0_n75, npu_inst_pe_1_4_0_n74,
         npu_inst_pe_1_4_0_n73, npu_inst_pe_1_4_0_n72, npu_inst_pe_1_4_0_n71,
         npu_inst_pe_1_4_0_n70, npu_inst_pe_1_4_0_n69, npu_inst_pe_1_4_0_n68,
         npu_inst_pe_1_4_0_n67, npu_inst_pe_1_4_0_n66, npu_inst_pe_1_4_0_n65,
         npu_inst_pe_1_4_0_n64, npu_inst_pe_1_4_0_n63, npu_inst_pe_1_4_0_n62,
         npu_inst_pe_1_4_0_n61, npu_inst_pe_1_4_0_n60, npu_inst_pe_1_4_0_n59,
         npu_inst_pe_1_4_0_n58, npu_inst_pe_1_4_0_n57, npu_inst_pe_1_4_0_n56,
         npu_inst_pe_1_4_0_n55, npu_inst_pe_1_4_0_n54, npu_inst_pe_1_4_0_n53,
         npu_inst_pe_1_4_0_n52, npu_inst_pe_1_4_0_n51, npu_inst_pe_1_4_0_n50,
         npu_inst_pe_1_4_0_n49, npu_inst_pe_1_4_0_n48, npu_inst_pe_1_4_0_n47,
         npu_inst_pe_1_4_0_n46, npu_inst_pe_1_4_0_n45, npu_inst_pe_1_4_0_n44,
         npu_inst_pe_1_4_0_n43, npu_inst_pe_1_4_0_n42, npu_inst_pe_1_4_0_n41,
         npu_inst_pe_1_4_0_n40, npu_inst_pe_1_4_0_n39, npu_inst_pe_1_4_0_n38,
         npu_inst_pe_1_4_0_n37, npu_inst_pe_1_4_0_n27, npu_inst_pe_1_4_0_n26,
         npu_inst_pe_1_4_0_net3748, npu_inst_pe_1_4_0_net3742,
         npu_inst_pe_1_4_0_N94, npu_inst_pe_1_4_0_N93, npu_inst_pe_1_4_0_N84,
         npu_inst_pe_1_4_0_N80, npu_inst_pe_1_4_0_N79, npu_inst_pe_1_4_0_N78,
         npu_inst_pe_1_4_0_N77, npu_inst_pe_1_4_0_N76, npu_inst_pe_1_4_0_N75,
         npu_inst_pe_1_4_0_N74, npu_inst_pe_1_4_0_N73, npu_inst_pe_1_4_0_N72,
         npu_inst_pe_1_4_0_N71, npu_inst_pe_1_4_0_N70, npu_inst_pe_1_4_0_N69,
         npu_inst_pe_1_4_0_N68, npu_inst_pe_1_4_0_N67, npu_inst_pe_1_4_0_N66,
         npu_inst_pe_1_4_0_N65, npu_inst_pe_1_4_0_int_data_0_,
         npu_inst_pe_1_4_0_int_data_1_, npu_inst_pe_1_4_0_int_q_weight_0_,
         npu_inst_pe_1_4_0_int_q_weight_1_,
         npu_inst_pe_1_4_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_0_int_q_reg_h_0__1_, npu_inst_pe_1_4_0_o_data_h_0_,
         npu_inst_pe_1_4_0_o_data_h_1_, npu_inst_pe_1_4_1_n118,
         npu_inst_pe_1_4_1_n117, npu_inst_pe_1_4_1_n116,
         npu_inst_pe_1_4_1_n115, npu_inst_pe_1_4_1_n114,
         npu_inst_pe_1_4_1_n113, npu_inst_pe_1_4_1_n112,
         npu_inst_pe_1_4_1_n111, npu_inst_pe_1_4_1_n110,
         npu_inst_pe_1_4_1_n109, npu_inst_pe_1_4_1_n108,
         npu_inst_pe_1_4_1_n107, npu_inst_pe_1_4_1_n106,
         npu_inst_pe_1_4_1_n105, npu_inst_pe_1_4_1_n104,
         npu_inst_pe_1_4_1_n103, npu_inst_pe_1_4_1_n102,
         npu_inst_pe_1_4_1_n101, npu_inst_pe_1_4_1_n100, npu_inst_pe_1_4_1_n99,
         npu_inst_pe_1_4_1_n98, npu_inst_pe_1_4_1_n36, npu_inst_pe_1_4_1_n35,
         npu_inst_pe_1_4_1_n34, npu_inst_pe_1_4_1_n33, npu_inst_pe_1_4_1_n32,
         npu_inst_pe_1_4_1_n31, npu_inst_pe_1_4_1_n30, npu_inst_pe_1_4_1_n29,
         npu_inst_pe_1_4_1_n28, npu_inst_pe_1_4_1_n25, npu_inst_pe_1_4_1_n24,
         npu_inst_pe_1_4_1_n23, npu_inst_pe_1_4_1_n22, npu_inst_pe_1_4_1_n21,
         npu_inst_pe_1_4_1_n20, npu_inst_pe_1_4_1_n19, npu_inst_pe_1_4_1_n18,
         npu_inst_pe_1_4_1_n17, npu_inst_pe_1_4_1_n16, npu_inst_pe_1_4_1_n15,
         npu_inst_pe_1_4_1_n14, npu_inst_pe_1_4_1_n13, npu_inst_pe_1_4_1_n12,
         npu_inst_pe_1_4_1_n11, npu_inst_pe_1_4_1_n10, npu_inst_pe_1_4_1_n9,
         npu_inst_pe_1_4_1_n8, npu_inst_pe_1_4_1_n7, npu_inst_pe_1_4_1_n6,
         npu_inst_pe_1_4_1_n5, npu_inst_pe_1_4_1_n4, npu_inst_pe_1_4_1_n3,
         npu_inst_pe_1_4_1_n2, npu_inst_pe_1_4_1_n1,
         npu_inst_pe_1_4_1_sub_77_carry_7_, npu_inst_pe_1_4_1_sub_77_carry_6_,
         npu_inst_pe_1_4_1_sub_77_carry_5_, npu_inst_pe_1_4_1_sub_77_carry_4_,
         npu_inst_pe_1_4_1_sub_77_carry_3_, npu_inst_pe_1_4_1_sub_77_carry_2_,
         npu_inst_pe_1_4_1_sub_77_carry_1_, npu_inst_pe_1_4_1_add_79_carry_7_,
         npu_inst_pe_1_4_1_add_79_carry_6_, npu_inst_pe_1_4_1_add_79_carry_5_,
         npu_inst_pe_1_4_1_add_79_carry_4_, npu_inst_pe_1_4_1_add_79_carry_3_,
         npu_inst_pe_1_4_1_add_79_carry_2_, npu_inst_pe_1_4_1_add_79_carry_1_,
         npu_inst_pe_1_4_1_n97, npu_inst_pe_1_4_1_n96, npu_inst_pe_1_4_1_n95,
         npu_inst_pe_1_4_1_n94, npu_inst_pe_1_4_1_n93, npu_inst_pe_1_4_1_n92,
         npu_inst_pe_1_4_1_n91, npu_inst_pe_1_4_1_n90, npu_inst_pe_1_4_1_n89,
         npu_inst_pe_1_4_1_n88, npu_inst_pe_1_4_1_n87, npu_inst_pe_1_4_1_n86,
         npu_inst_pe_1_4_1_n85, npu_inst_pe_1_4_1_n84, npu_inst_pe_1_4_1_n83,
         npu_inst_pe_1_4_1_n82, npu_inst_pe_1_4_1_n81, npu_inst_pe_1_4_1_n80,
         npu_inst_pe_1_4_1_n79, npu_inst_pe_1_4_1_n78, npu_inst_pe_1_4_1_n77,
         npu_inst_pe_1_4_1_n76, npu_inst_pe_1_4_1_n75, npu_inst_pe_1_4_1_n74,
         npu_inst_pe_1_4_1_n73, npu_inst_pe_1_4_1_n72, npu_inst_pe_1_4_1_n71,
         npu_inst_pe_1_4_1_n70, npu_inst_pe_1_4_1_n69, npu_inst_pe_1_4_1_n68,
         npu_inst_pe_1_4_1_n67, npu_inst_pe_1_4_1_n66, npu_inst_pe_1_4_1_n65,
         npu_inst_pe_1_4_1_n64, npu_inst_pe_1_4_1_n63, npu_inst_pe_1_4_1_n62,
         npu_inst_pe_1_4_1_n61, npu_inst_pe_1_4_1_n60, npu_inst_pe_1_4_1_n59,
         npu_inst_pe_1_4_1_n58, npu_inst_pe_1_4_1_n57, npu_inst_pe_1_4_1_n56,
         npu_inst_pe_1_4_1_n55, npu_inst_pe_1_4_1_n54, npu_inst_pe_1_4_1_n53,
         npu_inst_pe_1_4_1_n52, npu_inst_pe_1_4_1_n51, npu_inst_pe_1_4_1_n50,
         npu_inst_pe_1_4_1_n49, npu_inst_pe_1_4_1_n48, npu_inst_pe_1_4_1_n47,
         npu_inst_pe_1_4_1_n46, npu_inst_pe_1_4_1_n45, npu_inst_pe_1_4_1_n44,
         npu_inst_pe_1_4_1_n43, npu_inst_pe_1_4_1_n42, npu_inst_pe_1_4_1_n41,
         npu_inst_pe_1_4_1_n40, npu_inst_pe_1_4_1_n39, npu_inst_pe_1_4_1_n38,
         npu_inst_pe_1_4_1_n37, npu_inst_pe_1_4_1_n27, npu_inst_pe_1_4_1_n26,
         npu_inst_pe_1_4_1_net3725, npu_inst_pe_1_4_1_net3719,
         npu_inst_pe_1_4_1_N94, npu_inst_pe_1_4_1_N93, npu_inst_pe_1_4_1_N84,
         npu_inst_pe_1_4_1_N80, npu_inst_pe_1_4_1_N79, npu_inst_pe_1_4_1_N78,
         npu_inst_pe_1_4_1_N77, npu_inst_pe_1_4_1_N76, npu_inst_pe_1_4_1_N75,
         npu_inst_pe_1_4_1_N74, npu_inst_pe_1_4_1_N73, npu_inst_pe_1_4_1_N72,
         npu_inst_pe_1_4_1_N71, npu_inst_pe_1_4_1_N70, npu_inst_pe_1_4_1_N69,
         npu_inst_pe_1_4_1_N68, npu_inst_pe_1_4_1_N67, npu_inst_pe_1_4_1_N66,
         npu_inst_pe_1_4_1_N65, npu_inst_pe_1_4_1_int_data_0_,
         npu_inst_pe_1_4_1_int_data_1_, npu_inst_pe_1_4_1_int_q_weight_0_,
         npu_inst_pe_1_4_1_int_q_weight_1_,
         npu_inst_pe_1_4_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_1_int_q_reg_h_0__1_, npu_inst_pe_1_4_2_n118,
         npu_inst_pe_1_4_2_n117, npu_inst_pe_1_4_2_n116,
         npu_inst_pe_1_4_2_n115, npu_inst_pe_1_4_2_n114,
         npu_inst_pe_1_4_2_n113, npu_inst_pe_1_4_2_n112,
         npu_inst_pe_1_4_2_n111, npu_inst_pe_1_4_2_n110,
         npu_inst_pe_1_4_2_n109, npu_inst_pe_1_4_2_n108,
         npu_inst_pe_1_4_2_n107, npu_inst_pe_1_4_2_n106,
         npu_inst_pe_1_4_2_n105, npu_inst_pe_1_4_2_n104,
         npu_inst_pe_1_4_2_n103, npu_inst_pe_1_4_2_n102,
         npu_inst_pe_1_4_2_n101, npu_inst_pe_1_4_2_n100, npu_inst_pe_1_4_2_n99,
         npu_inst_pe_1_4_2_n98, npu_inst_pe_1_4_2_n36, npu_inst_pe_1_4_2_n35,
         npu_inst_pe_1_4_2_n34, npu_inst_pe_1_4_2_n33, npu_inst_pe_1_4_2_n32,
         npu_inst_pe_1_4_2_n31, npu_inst_pe_1_4_2_n30, npu_inst_pe_1_4_2_n29,
         npu_inst_pe_1_4_2_n28, npu_inst_pe_1_4_2_n25, npu_inst_pe_1_4_2_n24,
         npu_inst_pe_1_4_2_n23, npu_inst_pe_1_4_2_n22, npu_inst_pe_1_4_2_n21,
         npu_inst_pe_1_4_2_n20, npu_inst_pe_1_4_2_n19, npu_inst_pe_1_4_2_n18,
         npu_inst_pe_1_4_2_n17, npu_inst_pe_1_4_2_n16, npu_inst_pe_1_4_2_n15,
         npu_inst_pe_1_4_2_n14, npu_inst_pe_1_4_2_n13, npu_inst_pe_1_4_2_n12,
         npu_inst_pe_1_4_2_n11, npu_inst_pe_1_4_2_n10, npu_inst_pe_1_4_2_n9,
         npu_inst_pe_1_4_2_n8, npu_inst_pe_1_4_2_n7, npu_inst_pe_1_4_2_n6,
         npu_inst_pe_1_4_2_n5, npu_inst_pe_1_4_2_n4, npu_inst_pe_1_4_2_n3,
         npu_inst_pe_1_4_2_n2, npu_inst_pe_1_4_2_n1,
         npu_inst_pe_1_4_2_sub_77_carry_7_, npu_inst_pe_1_4_2_sub_77_carry_6_,
         npu_inst_pe_1_4_2_sub_77_carry_5_, npu_inst_pe_1_4_2_sub_77_carry_4_,
         npu_inst_pe_1_4_2_sub_77_carry_3_, npu_inst_pe_1_4_2_sub_77_carry_2_,
         npu_inst_pe_1_4_2_sub_77_carry_1_, npu_inst_pe_1_4_2_add_79_carry_7_,
         npu_inst_pe_1_4_2_add_79_carry_6_, npu_inst_pe_1_4_2_add_79_carry_5_,
         npu_inst_pe_1_4_2_add_79_carry_4_, npu_inst_pe_1_4_2_add_79_carry_3_,
         npu_inst_pe_1_4_2_add_79_carry_2_, npu_inst_pe_1_4_2_add_79_carry_1_,
         npu_inst_pe_1_4_2_n97, npu_inst_pe_1_4_2_n96, npu_inst_pe_1_4_2_n95,
         npu_inst_pe_1_4_2_n94, npu_inst_pe_1_4_2_n93, npu_inst_pe_1_4_2_n92,
         npu_inst_pe_1_4_2_n91, npu_inst_pe_1_4_2_n90, npu_inst_pe_1_4_2_n89,
         npu_inst_pe_1_4_2_n88, npu_inst_pe_1_4_2_n87, npu_inst_pe_1_4_2_n86,
         npu_inst_pe_1_4_2_n85, npu_inst_pe_1_4_2_n84, npu_inst_pe_1_4_2_n83,
         npu_inst_pe_1_4_2_n82, npu_inst_pe_1_4_2_n81, npu_inst_pe_1_4_2_n80,
         npu_inst_pe_1_4_2_n79, npu_inst_pe_1_4_2_n78, npu_inst_pe_1_4_2_n77,
         npu_inst_pe_1_4_2_n76, npu_inst_pe_1_4_2_n75, npu_inst_pe_1_4_2_n74,
         npu_inst_pe_1_4_2_n73, npu_inst_pe_1_4_2_n72, npu_inst_pe_1_4_2_n71,
         npu_inst_pe_1_4_2_n70, npu_inst_pe_1_4_2_n69, npu_inst_pe_1_4_2_n68,
         npu_inst_pe_1_4_2_n67, npu_inst_pe_1_4_2_n66, npu_inst_pe_1_4_2_n65,
         npu_inst_pe_1_4_2_n64, npu_inst_pe_1_4_2_n63, npu_inst_pe_1_4_2_n62,
         npu_inst_pe_1_4_2_n61, npu_inst_pe_1_4_2_n60, npu_inst_pe_1_4_2_n59,
         npu_inst_pe_1_4_2_n58, npu_inst_pe_1_4_2_n57, npu_inst_pe_1_4_2_n56,
         npu_inst_pe_1_4_2_n55, npu_inst_pe_1_4_2_n54, npu_inst_pe_1_4_2_n53,
         npu_inst_pe_1_4_2_n52, npu_inst_pe_1_4_2_n51, npu_inst_pe_1_4_2_n50,
         npu_inst_pe_1_4_2_n49, npu_inst_pe_1_4_2_n48, npu_inst_pe_1_4_2_n47,
         npu_inst_pe_1_4_2_n46, npu_inst_pe_1_4_2_n45, npu_inst_pe_1_4_2_n44,
         npu_inst_pe_1_4_2_n43, npu_inst_pe_1_4_2_n42, npu_inst_pe_1_4_2_n41,
         npu_inst_pe_1_4_2_n40, npu_inst_pe_1_4_2_n39, npu_inst_pe_1_4_2_n38,
         npu_inst_pe_1_4_2_n37, npu_inst_pe_1_4_2_n27, npu_inst_pe_1_4_2_n26,
         npu_inst_pe_1_4_2_net3702, npu_inst_pe_1_4_2_net3696,
         npu_inst_pe_1_4_2_N94, npu_inst_pe_1_4_2_N93, npu_inst_pe_1_4_2_N84,
         npu_inst_pe_1_4_2_N80, npu_inst_pe_1_4_2_N79, npu_inst_pe_1_4_2_N78,
         npu_inst_pe_1_4_2_N77, npu_inst_pe_1_4_2_N76, npu_inst_pe_1_4_2_N75,
         npu_inst_pe_1_4_2_N74, npu_inst_pe_1_4_2_N73, npu_inst_pe_1_4_2_N72,
         npu_inst_pe_1_4_2_N71, npu_inst_pe_1_4_2_N70, npu_inst_pe_1_4_2_N69,
         npu_inst_pe_1_4_2_N68, npu_inst_pe_1_4_2_N67, npu_inst_pe_1_4_2_N66,
         npu_inst_pe_1_4_2_N65, npu_inst_pe_1_4_2_int_data_0_,
         npu_inst_pe_1_4_2_int_data_1_, npu_inst_pe_1_4_2_int_q_weight_0_,
         npu_inst_pe_1_4_2_int_q_weight_1_,
         npu_inst_pe_1_4_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_2_int_q_reg_h_0__1_, npu_inst_pe_1_4_3_n118,
         npu_inst_pe_1_4_3_n117, npu_inst_pe_1_4_3_n116,
         npu_inst_pe_1_4_3_n115, npu_inst_pe_1_4_3_n114,
         npu_inst_pe_1_4_3_n113, npu_inst_pe_1_4_3_n112,
         npu_inst_pe_1_4_3_n111, npu_inst_pe_1_4_3_n110,
         npu_inst_pe_1_4_3_n109, npu_inst_pe_1_4_3_n108,
         npu_inst_pe_1_4_3_n107, npu_inst_pe_1_4_3_n106,
         npu_inst_pe_1_4_3_n105, npu_inst_pe_1_4_3_n104,
         npu_inst_pe_1_4_3_n103, npu_inst_pe_1_4_3_n102,
         npu_inst_pe_1_4_3_n101, npu_inst_pe_1_4_3_n100, npu_inst_pe_1_4_3_n99,
         npu_inst_pe_1_4_3_n98, npu_inst_pe_1_4_3_n36, npu_inst_pe_1_4_3_n35,
         npu_inst_pe_1_4_3_n34, npu_inst_pe_1_4_3_n33, npu_inst_pe_1_4_3_n32,
         npu_inst_pe_1_4_3_n31, npu_inst_pe_1_4_3_n30, npu_inst_pe_1_4_3_n29,
         npu_inst_pe_1_4_3_n28, npu_inst_pe_1_4_3_n25, npu_inst_pe_1_4_3_n24,
         npu_inst_pe_1_4_3_n23, npu_inst_pe_1_4_3_n22, npu_inst_pe_1_4_3_n21,
         npu_inst_pe_1_4_3_n20, npu_inst_pe_1_4_3_n19, npu_inst_pe_1_4_3_n18,
         npu_inst_pe_1_4_3_n17, npu_inst_pe_1_4_3_n16, npu_inst_pe_1_4_3_n15,
         npu_inst_pe_1_4_3_n14, npu_inst_pe_1_4_3_n13, npu_inst_pe_1_4_3_n12,
         npu_inst_pe_1_4_3_n11, npu_inst_pe_1_4_3_n10, npu_inst_pe_1_4_3_n9,
         npu_inst_pe_1_4_3_n8, npu_inst_pe_1_4_3_n7, npu_inst_pe_1_4_3_n6,
         npu_inst_pe_1_4_3_n5, npu_inst_pe_1_4_3_n4, npu_inst_pe_1_4_3_n3,
         npu_inst_pe_1_4_3_n2, npu_inst_pe_1_4_3_n1,
         npu_inst_pe_1_4_3_sub_77_carry_7_, npu_inst_pe_1_4_3_sub_77_carry_6_,
         npu_inst_pe_1_4_3_sub_77_carry_5_, npu_inst_pe_1_4_3_sub_77_carry_4_,
         npu_inst_pe_1_4_3_sub_77_carry_3_, npu_inst_pe_1_4_3_sub_77_carry_2_,
         npu_inst_pe_1_4_3_sub_77_carry_1_, npu_inst_pe_1_4_3_add_79_carry_7_,
         npu_inst_pe_1_4_3_add_79_carry_6_, npu_inst_pe_1_4_3_add_79_carry_5_,
         npu_inst_pe_1_4_3_add_79_carry_4_, npu_inst_pe_1_4_3_add_79_carry_3_,
         npu_inst_pe_1_4_3_add_79_carry_2_, npu_inst_pe_1_4_3_add_79_carry_1_,
         npu_inst_pe_1_4_3_n97, npu_inst_pe_1_4_3_n96, npu_inst_pe_1_4_3_n95,
         npu_inst_pe_1_4_3_n94, npu_inst_pe_1_4_3_n93, npu_inst_pe_1_4_3_n92,
         npu_inst_pe_1_4_3_n91, npu_inst_pe_1_4_3_n90, npu_inst_pe_1_4_3_n89,
         npu_inst_pe_1_4_3_n88, npu_inst_pe_1_4_3_n87, npu_inst_pe_1_4_3_n86,
         npu_inst_pe_1_4_3_n85, npu_inst_pe_1_4_3_n84, npu_inst_pe_1_4_3_n83,
         npu_inst_pe_1_4_3_n82, npu_inst_pe_1_4_3_n81, npu_inst_pe_1_4_3_n80,
         npu_inst_pe_1_4_3_n79, npu_inst_pe_1_4_3_n78, npu_inst_pe_1_4_3_n77,
         npu_inst_pe_1_4_3_n76, npu_inst_pe_1_4_3_n75, npu_inst_pe_1_4_3_n74,
         npu_inst_pe_1_4_3_n73, npu_inst_pe_1_4_3_n72, npu_inst_pe_1_4_3_n71,
         npu_inst_pe_1_4_3_n70, npu_inst_pe_1_4_3_n69, npu_inst_pe_1_4_3_n68,
         npu_inst_pe_1_4_3_n67, npu_inst_pe_1_4_3_n66, npu_inst_pe_1_4_3_n65,
         npu_inst_pe_1_4_3_n64, npu_inst_pe_1_4_3_n63, npu_inst_pe_1_4_3_n62,
         npu_inst_pe_1_4_3_n61, npu_inst_pe_1_4_3_n60, npu_inst_pe_1_4_3_n59,
         npu_inst_pe_1_4_3_n58, npu_inst_pe_1_4_3_n57, npu_inst_pe_1_4_3_n56,
         npu_inst_pe_1_4_3_n55, npu_inst_pe_1_4_3_n54, npu_inst_pe_1_4_3_n53,
         npu_inst_pe_1_4_3_n52, npu_inst_pe_1_4_3_n51, npu_inst_pe_1_4_3_n50,
         npu_inst_pe_1_4_3_n49, npu_inst_pe_1_4_3_n48, npu_inst_pe_1_4_3_n47,
         npu_inst_pe_1_4_3_n46, npu_inst_pe_1_4_3_n45, npu_inst_pe_1_4_3_n44,
         npu_inst_pe_1_4_3_n43, npu_inst_pe_1_4_3_n42, npu_inst_pe_1_4_3_n41,
         npu_inst_pe_1_4_3_n40, npu_inst_pe_1_4_3_n39, npu_inst_pe_1_4_3_n38,
         npu_inst_pe_1_4_3_n37, npu_inst_pe_1_4_3_n27, npu_inst_pe_1_4_3_n26,
         npu_inst_pe_1_4_3_net3679, npu_inst_pe_1_4_3_net3673,
         npu_inst_pe_1_4_3_N94, npu_inst_pe_1_4_3_N93, npu_inst_pe_1_4_3_N84,
         npu_inst_pe_1_4_3_N80, npu_inst_pe_1_4_3_N79, npu_inst_pe_1_4_3_N78,
         npu_inst_pe_1_4_3_N77, npu_inst_pe_1_4_3_N76, npu_inst_pe_1_4_3_N75,
         npu_inst_pe_1_4_3_N74, npu_inst_pe_1_4_3_N73, npu_inst_pe_1_4_3_N72,
         npu_inst_pe_1_4_3_N71, npu_inst_pe_1_4_3_N70, npu_inst_pe_1_4_3_N69,
         npu_inst_pe_1_4_3_N68, npu_inst_pe_1_4_3_N67, npu_inst_pe_1_4_3_N66,
         npu_inst_pe_1_4_3_N65, npu_inst_pe_1_4_3_int_data_0_,
         npu_inst_pe_1_4_3_int_data_1_, npu_inst_pe_1_4_3_int_q_weight_0_,
         npu_inst_pe_1_4_3_int_q_weight_1_,
         npu_inst_pe_1_4_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_3_int_q_reg_h_0__1_, npu_inst_pe_1_4_4_n118,
         npu_inst_pe_1_4_4_n117, npu_inst_pe_1_4_4_n116,
         npu_inst_pe_1_4_4_n115, npu_inst_pe_1_4_4_n114,
         npu_inst_pe_1_4_4_n113, npu_inst_pe_1_4_4_n112,
         npu_inst_pe_1_4_4_n111, npu_inst_pe_1_4_4_n110,
         npu_inst_pe_1_4_4_n109, npu_inst_pe_1_4_4_n108,
         npu_inst_pe_1_4_4_n107, npu_inst_pe_1_4_4_n106,
         npu_inst_pe_1_4_4_n105, npu_inst_pe_1_4_4_n104,
         npu_inst_pe_1_4_4_n103, npu_inst_pe_1_4_4_n102,
         npu_inst_pe_1_4_4_n101, npu_inst_pe_1_4_4_n100, npu_inst_pe_1_4_4_n99,
         npu_inst_pe_1_4_4_n98, npu_inst_pe_1_4_4_n36, npu_inst_pe_1_4_4_n35,
         npu_inst_pe_1_4_4_n34, npu_inst_pe_1_4_4_n33, npu_inst_pe_1_4_4_n32,
         npu_inst_pe_1_4_4_n31, npu_inst_pe_1_4_4_n30, npu_inst_pe_1_4_4_n29,
         npu_inst_pe_1_4_4_n28, npu_inst_pe_1_4_4_n25, npu_inst_pe_1_4_4_n24,
         npu_inst_pe_1_4_4_n23, npu_inst_pe_1_4_4_n22, npu_inst_pe_1_4_4_n21,
         npu_inst_pe_1_4_4_n20, npu_inst_pe_1_4_4_n19, npu_inst_pe_1_4_4_n18,
         npu_inst_pe_1_4_4_n17, npu_inst_pe_1_4_4_n16, npu_inst_pe_1_4_4_n15,
         npu_inst_pe_1_4_4_n14, npu_inst_pe_1_4_4_n13, npu_inst_pe_1_4_4_n12,
         npu_inst_pe_1_4_4_n11, npu_inst_pe_1_4_4_n10, npu_inst_pe_1_4_4_n9,
         npu_inst_pe_1_4_4_n8, npu_inst_pe_1_4_4_n7, npu_inst_pe_1_4_4_n6,
         npu_inst_pe_1_4_4_n5, npu_inst_pe_1_4_4_n4, npu_inst_pe_1_4_4_n3,
         npu_inst_pe_1_4_4_n2, npu_inst_pe_1_4_4_n1,
         npu_inst_pe_1_4_4_sub_77_carry_7_, npu_inst_pe_1_4_4_sub_77_carry_6_,
         npu_inst_pe_1_4_4_sub_77_carry_5_, npu_inst_pe_1_4_4_sub_77_carry_4_,
         npu_inst_pe_1_4_4_sub_77_carry_3_, npu_inst_pe_1_4_4_sub_77_carry_2_,
         npu_inst_pe_1_4_4_sub_77_carry_1_, npu_inst_pe_1_4_4_add_79_carry_7_,
         npu_inst_pe_1_4_4_add_79_carry_6_, npu_inst_pe_1_4_4_add_79_carry_5_,
         npu_inst_pe_1_4_4_add_79_carry_4_, npu_inst_pe_1_4_4_add_79_carry_3_,
         npu_inst_pe_1_4_4_add_79_carry_2_, npu_inst_pe_1_4_4_add_79_carry_1_,
         npu_inst_pe_1_4_4_n97, npu_inst_pe_1_4_4_n96, npu_inst_pe_1_4_4_n95,
         npu_inst_pe_1_4_4_n94, npu_inst_pe_1_4_4_n93, npu_inst_pe_1_4_4_n92,
         npu_inst_pe_1_4_4_n91, npu_inst_pe_1_4_4_n90, npu_inst_pe_1_4_4_n89,
         npu_inst_pe_1_4_4_n88, npu_inst_pe_1_4_4_n87, npu_inst_pe_1_4_4_n86,
         npu_inst_pe_1_4_4_n85, npu_inst_pe_1_4_4_n84, npu_inst_pe_1_4_4_n83,
         npu_inst_pe_1_4_4_n82, npu_inst_pe_1_4_4_n81, npu_inst_pe_1_4_4_n80,
         npu_inst_pe_1_4_4_n79, npu_inst_pe_1_4_4_n78, npu_inst_pe_1_4_4_n77,
         npu_inst_pe_1_4_4_n76, npu_inst_pe_1_4_4_n75, npu_inst_pe_1_4_4_n74,
         npu_inst_pe_1_4_4_n73, npu_inst_pe_1_4_4_n72, npu_inst_pe_1_4_4_n71,
         npu_inst_pe_1_4_4_n70, npu_inst_pe_1_4_4_n69, npu_inst_pe_1_4_4_n68,
         npu_inst_pe_1_4_4_n67, npu_inst_pe_1_4_4_n66, npu_inst_pe_1_4_4_n65,
         npu_inst_pe_1_4_4_n64, npu_inst_pe_1_4_4_n63, npu_inst_pe_1_4_4_n62,
         npu_inst_pe_1_4_4_n61, npu_inst_pe_1_4_4_n60, npu_inst_pe_1_4_4_n59,
         npu_inst_pe_1_4_4_n58, npu_inst_pe_1_4_4_n57, npu_inst_pe_1_4_4_n56,
         npu_inst_pe_1_4_4_n55, npu_inst_pe_1_4_4_n54, npu_inst_pe_1_4_4_n53,
         npu_inst_pe_1_4_4_n52, npu_inst_pe_1_4_4_n51, npu_inst_pe_1_4_4_n50,
         npu_inst_pe_1_4_4_n49, npu_inst_pe_1_4_4_n48, npu_inst_pe_1_4_4_n47,
         npu_inst_pe_1_4_4_n46, npu_inst_pe_1_4_4_n45, npu_inst_pe_1_4_4_n44,
         npu_inst_pe_1_4_4_n43, npu_inst_pe_1_4_4_n42, npu_inst_pe_1_4_4_n41,
         npu_inst_pe_1_4_4_n40, npu_inst_pe_1_4_4_n39, npu_inst_pe_1_4_4_n38,
         npu_inst_pe_1_4_4_n37, npu_inst_pe_1_4_4_n27, npu_inst_pe_1_4_4_n26,
         npu_inst_pe_1_4_4_net3656, npu_inst_pe_1_4_4_net3650,
         npu_inst_pe_1_4_4_N94, npu_inst_pe_1_4_4_N93, npu_inst_pe_1_4_4_N84,
         npu_inst_pe_1_4_4_N80, npu_inst_pe_1_4_4_N79, npu_inst_pe_1_4_4_N78,
         npu_inst_pe_1_4_4_N77, npu_inst_pe_1_4_4_N76, npu_inst_pe_1_4_4_N75,
         npu_inst_pe_1_4_4_N74, npu_inst_pe_1_4_4_N73, npu_inst_pe_1_4_4_N72,
         npu_inst_pe_1_4_4_N71, npu_inst_pe_1_4_4_N70, npu_inst_pe_1_4_4_N69,
         npu_inst_pe_1_4_4_N68, npu_inst_pe_1_4_4_N67, npu_inst_pe_1_4_4_N66,
         npu_inst_pe_1_4_4_N65, npu_inst_pe_1_4_4_int_data_0_,
         npu_inst_pe_1_4_4_int_data_1_, npu_inst_pe_1_4_4_int_q_weight_0_,
         npu_inst_pe_1_4_4_int_q_weight_1_,
         npu_inst_pe_1_4_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_4_int_q_reg_h_0__1_, npu_inst_pe_1_4_5_n118,
         npu_inst_pe_1_4_5_n117, npu_inst_pe_1_4_5_n116,
         npu_inst_pe_1_4_5_n115, npu_inst_pe_1_4_5_n114,
         npu_inst_pe_1_4_5_n113, npu_inst_pe_1_4_5_n112,
         npu_inst_pe_1_4_5_n111, npu_inst_pe_1_4_5_n110,
         npu_inst_pe_1_4_5_n109, npu_inst_pe_1_4_5_n108,
         npu_inst_pe_1_4_5_n107, npu_inst_pe_1_4_5_n106,
         npu_inst_pe_1_4_5_n105, npu_inst_pe_1_4_5_n104,
         npu_inst_pe_1_4_5_n103, npu_inst_pe_1_4_5_n102,
         npu_inst_pe_1_4_5_n101, npu_inst_pe_1_4_5_n100, npu_inst_pe_1_4_5_n99,
         npu_inst_pe_1_4_5_n98, npu_inst_pe_1_4_5_n36, npu_inst_pe_1_4_5_n35,
         npu_inst_pe_1_4_5_n34, npu_inst_pe_1_4_5_n33, npu_inst_pe_1_4_5_n32,
         npu_inst_pe_1_4_5_n31, npu_inst_pe_1_4_5_n30, npu_inst_pe_1_4_5_n29,
         npu_inst_pe_1_4_5_n28, npu_inst_pe_1_4_5_n25, npu_inst_pe_1_4_5_n24,
         npu_inst_pe_1_4_5_n23, npu_inst_pe_1_4_5_n22, npu_inst_pe_1_4_5_n21,
         npu_inst_pe_1_4_5_n20, npu_inst_pe_1_4_5_n19, npu_inst_pe_1_4_5_n18,
         npu_inst_pe_1_4_5_n17, npu_inst_pe_1_4_5_n16, npu_inst_pe_1_4_5_n15,
         npu_inst_pe_1_4_5_n14, npu_inst_pe_1_4_5_n13, npu_inst_pe_1_4_5_n12,
         npu_inst_pe_1_4_5_n11, npu_inst_pe_1_4_5_n10, npu_inst_pe_1_4_5_n9,
         npu_inst_pe_1_4_5_n8, npu_inst_pe_1_4_5_n7, npu_inst_pe_1_4_5_n6,
         npu_inst_pe_1_4_5_n5, npu_inst_pe_1_4_5_n4, npu_inst_pe_1_4_5_n3,
         npu_inst_pe_1_4_5_n2, npu_inst_pe_1_4_5_n1,
         npu_inst_pe_1_4_5_sub_77_carry_7_, npu_inst_pe_1_4_5_sub_77_carry_6_,
         npu_inst_pe_1_4_5_sub_77_carry_5_, npu_inst_pe_1_4_5_sub_77_carry_4_,
         npu_inst_pe_1_4_5_sub_77_carry_3_, npu_inst_pe_1_4_5_sub_77_carry_2_,
         npu_inst_pe_1_4_5_sub_77_carry_1_, npu_inst_pe_1_4_5_add_79_carry_7_,
         npu_inst_pe_1_4_5_add_79_carry_6_, npu_inst_pe_1_4_5_add_79_carry_5_,
         npu_inst_pe_1_4_5_add_79_carry_4_, npu_inst_pe_1_4_5_add_79_carry_3_,
         npu_inst_pe_1_4_5_add_79_carry_2_, npu_inst_pe_1_4_5_add_79_carry_1_,
         npu_inst_pe_1_4_5_n97, npu_inst_pe_1_4_5_n96, npu_inst_pe_1_4_5_n95,
         npu_inst_pe_1_4_5_n94, npu_inst_pe_1_4_5_n93, npu_inst_pe_1_4_5_n92,
         npu_inst_pe_1_4_5_n91, npu_inst_pe_1_4_5_n90, npu_inst_pe_1_4_5_n89,
         npu_inst_pe_1_4_5_n88, npu_inst_pe_1_4_5_n87, npu_inst_pe_1_4_5_n86,
         npu_inst_pe_1_4_5_n85, npu_inst_pe_1_4_5_n84, npu_inst_pe_1_4_5_n83,
         npu_inst_pe_1_4_5_n82, npu_inst_pe_1_4_5_n81, npu_inst_pe_1_4_5_n80,
         npu_inst_pe_1_4_5_n79, npu_inst_pe_1_4_5_n78, npu_inst_pe_1_4_5_n77,
         npu_inst_pe_1_4_5_n76, npu_inst_pe_1_4_5_n75, npu_inst_pe_1_4_5_n74,
         npu_inst_pe_1_4_5_n73, npu_inst_pe_1_4_5_n72, npu_inst_pe_1_4_5_n71,
         npu_inst_pe_1_4_5_n70, npu_inst_pe_1_4_5_n69, npu_inst_pe_1_4_5_n68,
         npu_inst_pe_1_4_5_n67, npu_inst_pe_1_4_5_n66, npu_inst_pe_1_4_5_n65,
         npu_inst_pe_1_4_5_n64, npu_inst_pe_1_4_5_n63, npu_inst_pe_1_4_5_n62,
         npu_inst_pe_1_4_5_n61, npu_inst_pe_1_4_5_n60, npu_inst_pe_1_4_5_n59,
         npu_inst_pe_1_4_5_n58, npu_inst_pe_1_4_5_n57, npu_inst_pe_1_4_5_n56,
         npu_inst_pe_1_4_5_n55, npu_inst_pe_1_4_5_n54, npu_inst_pe_1_4_5_n53,
         npu_inst_pe_1_4_5_n52, npu_inst_pe_1_4_5_n51, npu_inst_pe_1_4_5_n50,
         npu_inst_pe_1_4_5_n49, npu_inst_pe_1_4_5_n48, npu_inst_pe_1_4_5_n47,
         npu_inst_pe_1_4_5_n46, npu_inst_pe_1_4_5_n45, npu_inst_pe_1_4_5_n44,
         npu_inst_pe_1_4_5_n43, npu_inst_pe_1_4_5_n42, npu_inst_pe_1_4_5_n41,
         npu_inst_pe_1_4_5_n40, npu_inst_pe_1_4_5_n39, npu_inst_pe_1_4_5_n38,
         npu_inst_pe_1_4_5_n37, npu_inst_pe_1_4_5_n27, npu_inst_pe_1_4_5_n26,
         npu_inst_pe_1_4_5_net3633, npu_inst_pe_1_4_5_net3627,
         npu_inst_pe_1_4_5_N94, npu_inst_pe_1_4_5_N93, npu_inst_pe_1_4_5_N84,
         npu_inst_pe_1_4_5_N80, npu_inst_pe_1_4_5_N79, npu_inst_pe_1_4_5_N78,
         npu_inst_pe_1_4_5_N77, npu_inst_pe_1_4_5_N76, npu_inst_pe_1_4_5_N75,
         npu_inst_pe_1_4_5_N74, npu_inst_pe_1_4_5_N73, npu_inst_pe_1_4_5_N72,
         npu_inst_pe_1_4_5_N71, npu_inst_pe_1_4_5_N70, npu_inst_pe_1_4_5_N69,
         npu_inst_pe_1_4_5_N68, npu_inst_pe_1_4_5_N67, npu_inst_pe_1_4_5_N66,
         npu_inst_pe_1_4_5_N65, npu_inst_pe_1_4_5_int_data_0_,
         npu_inst_pe_1_4_5_int_data_1_, npu_inst_pe_1_4_5_int_q_weight_0_,
         npu_inst_pe_1_4_5_int_q_weight_1_,
         npu_inst_pe_1_4_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_5_int_q_reg_h_0__1_, npu_inst_pe_1_4_6_n118,
         npu_inst_pe_1_4_6_n117, npu_inst_pe_1_4_6_n116,
         npu_inst_pe_1_4_6_n115, npu_inst_pe_1_4_6_n114,
         npu_inst_pe_1_4_6_n113, npu_inst_pe_1_4_6_n112,
         npu_inst_pe_1_4_6_n111, npu_inst_pe_1_4_6_n110,
         npu_inst_pe_1_4_6_n109, npu_inst_pe_1_4_6_n108,
         npu_inst_pe_1_4_6_n107, npu_inst_pe_1_4_6_n106,
         npu_inst_pe_1_4_6_n105, npu_inst_pe_1_4_6_n104,
         npu_inst_pe_1_4_6_n103, npu_inst_pe_1_4_6_n102,
         npu_inst_pe_1_4_6_n101, npu_inst_pe_1_4_6_n100, npu_inst_pe_1_4_6_n99,
         npu_inst_pe_1_4_6_n98, npu_inst_pe_1_4_6_n36, npu_inst_pe_1_4_6_n35,
         npu_inst_pe_1_4_6_n34, npu_inst_pe_1_4_6_n33, npu_inst_pe_1_4_6_n32,
         npu_inst_pe_1_4_6_n31, npu_inst_pe_1_4_6_n30, npu_inst_pe_1_4_6_n29,
         npu_inst_pe_1_4_6_n28, npu_inst_pe_1_4_6_n25, npu_inst_pe_1_4_6_n24,
         npu_inst_pe_1_4_6_n23, npu_inst_pe_1_4_6_n22, npu_inst_pe_1_4_6_n21,
         npu_inst_pe_1_4_6_n20, npu_inst_pe_1_4_6_n19, npu_inst_pe_1_4_6_n18,
         npu_inst_pe_1_4_6_n17, npu_inst_pe_1_4_6_n16, npu_inst_pe_1_4_6_n15,
         npu_inst_pe_1_4_6_n14, npu_inst_pe_1_4_6_n13, npu_inst_pe_1_4_6_n12,
         npu_inst_pe_1_4_6_n11, npu_inst_pe_1_4_6_n10, npu_inst_pe_1_4_6_n9,
         npu_inst_pe_1_4_6_n8, npu_inst_pe_1_4_6_n7, npu_inst_pe_1_4_6_n6,
         npu_inst_pe_1_4_6_n5, npu_inst_pe_1_4_6_n4, npu_inst_pe_1_4_6_n3,
         npu_inst_pe_1_4_6_n2, npu_inst_pe_1_4_6_n1,
         npu_inst_pe_1_4_6_sub_77_carry_7_, npu_inst_pe_1_4_6_sub_77_carry_6_,
         npu_inst_pe_1_4_6_sub_77_carry_5_, npu_inst_pe_1_4_6_sub_77_carry_4_,
         npu_inst_pe_1_4_6_sub_77_carry_3_, npu_inst_pe_1_4_6_sub_77_carry_2_,
         npu_inst_pe_1_4_6_sub_77_carry_1_, npu_inst_pe_1_4_6_add_79_carry_7_,
         npu_inst_pe_1_4_6_add_79_carry_6_, npu_inst_pe_1_4_6_add_79_carry_5_,
         npu_inst_pe_1_4_6_add_79_carry_4_, npu_inst_pe_1_4_6_add_79_carry_3_,
         npu_inst_pe_1_4_6_add_79_carry_2_, npu_inst_pe_1_4_6_add_79_carry_1_,
         npu_inst_pe_1_4_6_n97, npu_inst_pe_1_4_6_n96, npu_inst_pe_1_4_6_n95,
         npu_inst_pe_1_4_6_n94, npu_inst_pe_1_4_6_n93, npu_inst_pe_1_4_6_n92,
         npu_inst_pe_1_4_6_n91, npu_inst_pe_1_4_6_n90, npu_inst_pe_1_4_6_n89,
         npu_inst_pe_1_4_6_n88, npu_inst_pe_1_4_6_n87, npu_inst_pe_1_4_6_n86,
         npu_inst_pe_1_4_6_n85, npu_inst_pe_1_4_6_n84, npu_inst_pe_1_4_6_n83,
         npu_inst_pe_1_4_6_n82, npu_inst_pe_1_4_6_n81, npu_inst_pe_1_4_6_n80,
         npu_inst_pe_1_4_6_n79, npu_inst_pe_1_4_6_n78, npu_inst_pe_1_4_6_n77,
         npu_inst_pe_1_4_6_n76, npu_inst_pe_1_4_6_n75, npu_inst_pe_1_4_6_n74,
         npu_inst_pe_1_4_6_n73, npu_inst_pe_1_4_6_n72, npu_inst_pe_1_4_6_n71,
         npu_inst_pe_1_4_6_n70, npu_inst_pe_1_4_6_n69, npu_inst_pe_1_4_6_n68,
         npu_inst_pe_1_4_6_n67, npu_inst_pe_1_4_6_n66, npu_inst_pe_1_4_6_n65,
         npu_inst_pe_1_4_6_n64, npu_inst_pe_1_4_6_n63, npu_inst_pe_1_4_6_n62,
         npu_inst_pe_1_4_6_n61, npu_inst_pe_1_4_6_n60, npu_inst_pe_1_4_6_n59,
         npu_inst_pe_1_4_6_n58, npu_inst_pe_1_4_6_n57, npu_inst_pe_1_4_6_n56,
         npu_inst_pe_1_4_6_n55, npu_inst_pe_1_4_6_n54, npu_inst_pe_1_4_6_n53,
         npu_inst_pe_1_4_6_n52, npu_inst_pe_1_4_6_n51, npu_inst_pe_1_4_6_n50,
         npu_inst_pe_1_4_6_n49, npu_inst_pe_1_4_6_n48, npu_inst_pe_1_4_6_n47,
         npu_inst_pe_1_4_6_n46, npu_inst_pe_1_4_6_n45, npu_inst_pe_1_4_6_n44,
         npu_inst_pe_1_4_6_n43, npu_inst_pe_1_4_6_n42, npu_inst_pe_1_4_6_n41,
         npu_inst_pe_1_4_6_n40, npu_inst_pe_1_4_6_n39, npu_inst_pe_1_4_6_n38,
         npu_inst_pe_1_4_6_n37, npu_inst_pe_1_4_6_n27, npu_inst_pe_1_4_6_n26,
         npu_inst_pe_1_4_6_net3610, npu_inst_pe_1_4_6_net3604,
         npu_inst_pe_1_4_6_N94, npu_inst_pe_1_4_6_N93, npu_inst_pe_1_4_6_N84,
         npu_inst_pe_1_4_6_N80, npu_inst_pe_1_4_6_N79, npu_inst_pe_1_4_6_N78,
         npu_inst_pe_1_4_6_N77, npu_inst_pe_1_4_6_N76, npu_inst_pe_1_4_6_N75,
         npu_inst_pe_1_4_6_N74, npu_inst_pe_1_4_6_N73, npu_inst_pe_1_4_6_N72,
         npu_inst_pe_1_4_6_N71, npu_inst_pe_1_4_6_N70, npu_inst_pe_1_4_6_N69,
         npu_inst_pe_1_4_6_N68, npu_inst_pe_1_4_6_N67, npu_inst_pe_1_4_6_N66,
         npu_inst_pe_1_4_6_N65, npu_inst_pe_1_4_6_int_data_0_,
         npu_inst_pe_1_4_6_int_data_1_, npu_inst_pe_1_4_6_int_q_weight_0_,
         npu_inst_pe_1_4_6_int_q_weight_1_,
         npu_inst_pe_1_4_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_6_int_q_reg_h_0__1_, npu_inst_pe_1_4_7_n118,
         npu_inst_pe_1_4_7_n117, npu_inst_pe_1_4_7_n116,
         npu_inst_pe_1_4_7_n115, npu_inst_pe_1_4_7_n114,
         npu_inst_pe_1_4_7_n113, npu_inst_pe_1_4_7_n112,
         npu_inst_pe_1_4_7_n111, npu_inst_pe_1_4_7_n110,
         npu_inst_pe_1_4_7_n109, npu_inst_pe_1_4_7_n108,
         npu_inst_pe_1_4_7_n107, npu_inst_pe_1_4_7_n106,
         npu_inst_pe_1_4_7_n105, npu_inst_pe_1_4_7_n104,
         npu_inst_pe_1_4_7_n103, npu_inst_pe_1_4_7_n102,
         npu_inst_pe_1_4_7_n101, npu_inst_pe_1_4_7_n100, npu_inst_pe_1_4_7_n99,
         npu_inst_pe_1_4_7_n98, npu_inst_pe_1_4_7_n36, npu_inst_pe_1_4_7_n35,
         npu_inst_pe_1_4_7_n34, npu_inst_pe_1_4_7_n33, npu_inst_pe_1_4_7_n32,
         npu_inst_pe_1_4_7_n31, npu_inst_pe_1_4_7_n30, npu_inst_pe_1_4_7_n29,
         npu_inst_pe_1_4_7_n28, npu_inst_pe_1_4_7_n25, npu_inst_pe_1_4_7_n24,
         npu_inst_pe_1_4_7_n23, npu_inst_pe_1_4_7_n22, npu_inst_pe_1_4_7_n21,
         npu_inst_pe_1_4_7_n20, npu_inst_pe_1_4_7_n19, npu_inst_pe_1_4_7_n18,
         npu_inst_pe_1_4_7_n17, npu_inst_pe_1_4_7_n16, npu_inst_pe_1_4_7_n15,
         npu_inst_pe_1_4_7_n14, npu_inst_pe_1_4_7_n13, npu_inst_pe_1_4_7_n12,
         npu_inst_pe_1_4_7_n11, npu_inst_pe_1_4_7_n10, npu_inst_pe_1_4_7_n9,
         npu_inst_pe_1_4_7_n8, npu_inst_pe_1_4_7_n7, npu_inst_pe_1_4_7_n6,
         npu_inst_pe_1_4_7_n5, npu_inst_pe_1_4_7_n4, npu_inst_pe_1_4_7_n3,
         npu_inst_pe_1_4_7_n2, npu_inst_pe_1_4_7_n1,
         npu_inst_pe_1_4_7_sub_77_carry_7_, npu_inst_pe_1_4_7_sub_77_carry_6_,
         npu_inst_pe_1_4_7_sub_77_carry_5_, npu_inst_pe_1_4_7_sub_77_carry_4_,
         npu_inst_pe_1_4_7_sub_77_carry_3_, npu_inst_pe_1_4_7_sub_77_carry_2_,
         npu_inst_pe_1_4_7_sub_77_carry_1_, npu_inst_pe_1_4_7_add_79_carry_7_,
         npu_inst_pe_1_4_7_add_79_carry_6_, npu_inst_pe_1_4_7_add_79_carry_5_,
         npu_inst_pe_1_4_7_add_79_carry_4_, npu_inst_pe_1_4_7_add_79_carry_3_,
         npu_inst_pe_1_4_7_add_79_carry_2_, npu_inst_pe_1_4_7_add_79_carry_1_,
         npu_inst_pe_1_4_7_n97, npu_inst_pe_1_4_7_n96, npu_inst_pe_1_4_7_n95,
         npu_inst_pe_1_4_7_n94, npu_inst_pe_1_4_7_n93, npu_inst_pe_1_4_7_n92,
         npu_inst_pe_1_4_7_n91, npu_inst_pe_1_4_7_n90, npu_inst_pe_1_4_7_n89,
         npu_inst_pe_1_4_7_n88, npu_inst_pe_1_4_7_n87, npu_inst_pe_1_4_7_n86,
         npu_inst_pe_1_4_7_n85, npu_inst_pe_1_4_7_n84, npu_inst_pe_1_4_7_n83,
         npu_inst_pe_1_4_7_n82, npu_inst_pe_1_4_7_n81, npu_inst_pe_1_4_7_n80,
         npu_inst_pe_1_4_7_n79, npu_inst_pe_1_4_7_n78, npu_inst_pe_1_4_7_n77,
         npu_inst_pe_1_4_7_n76, npu_inst_pe_1_4_7_n75, npu_inst_pe_1_4_7_n74,
         npu_inst_pe_1_4_7_n73, npu_inst_pe_1_4_7_n72, npu_inst_pe_1_4_7_n71,
         npu_inst_pe_1_4_7_n70, npu_inst_pe_1_4_7_n69, npu_inst_pe_1_4_7_n68,
         npu_inst_pe_1_4_7_n67, npu_inst_pe_1_4_7_n66, npu_inst_pe_1_4_7_n65,
         npu_inst_pe_1_4_7_n64, npu_inst_pe_1_4_7_n63, npu_inst_pe_1_4_7_n62,
         npu_inst_pe_1_4_7_n61, npu_inst_pe_1_4_7_n60, npu_inst_pe_1_4_7_n59,
         npu_inst_pe_1_4_7_n58, npu_inst_pe_1_4_7_n57, npu_inst_pe_1_4_7_n56,
         npu_inst_pe_1_4_7_n55, npu_inst_pe_1_4_7_n54, npu_inst_pe_1_4_7_n53,
         npu_inst_pe_1_4_7_n52, npu_inst_pe_1_4_7_n51, npu_inst_pe_1_4_7_n50,
         npu_inst_pe_1_4_7_n49, npu_inst_pe_1_4_7_n48, npu_inst_pe_1_4_7_n47,
         npu_inst_pe_1_4_7_n46, npu_inst_pe_1_4_7_n45, npu_inst_pe_1_4_7_n44,
         npu_inst_pe_1_4_7_n43, npu_inst_pe_1_4_7_n42, npu_inst_pe_1_4_7_n41,
         npu_inst_pe_1_4_7_n40, npu_inst_pe_1_4_7_n39, npu_inst_pe_1_4_7_n38,
         npu_inst_pe_1_4_7_n37, npu_inst_pe_1_4_7_n27, npu_inst_pe_1_4_7_n26,
         npu_inst_pe_1_4_7_net3587, npu_inst_pe_1_4_7_net3581,
         npu_inst_pe_1_4_7_N94, npu_inst_pe_1_4_7_N93, npu_inst_pe_1_4_7_N84,
         npu_inst_pe_1_4_7_N80, npu_inst_pe_1_4_7_N79, npu_inst_pe_1_4_7_N78,
         npu_inst_pe_1_4_7_N77, npu_inst_pe_1_4_7_N76, npu_inst_pe_1_4_7_N75,
         npu_inst_pe_1_4_7_N74, npu_inst_pe_1_4_7_N73, npu_inst_pe_1_4_7_N72,
         npu_inst_pe_1_4_7_N71, npu_inst_pe_1_4_7_N70, npu_inst_pe_1_4_7_N69,
         npu_inst_pe_1_4_7_N68, npu_inst_pe_1_4_7_N67, npu_inst_pe_1_4_7_N66,
         npu_inst_pe_1_4_7_N65, npu_inst_pe_1_4_7_int_data_0_,
         npu_inst_pe_1_4_7_int_data_1_, npu_inst_pe_1_4_7_int_q_weight_0_,
         npu_inst_pe_1_4_7_int_q_weight_1_,
         npu_inst_pe_1_4_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_4_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_4_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_4_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_4_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_4_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_4_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_4_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_4_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_4_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_4_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_4_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_4_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_4_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_4_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_4_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_4_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_4_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_4_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_4_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_4_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_4_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_4_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_4_7_int_q_reg_h_0__1_, npu_inst_pe_1_5_0_n117,
         npu_inst_pe_1_5_0_n116, npu_inst_pe_1_5_0_n115,
         npu_inst_pe_1_5_0_n114, npu_inst_pe_1_5_0_n113,
         npu_inst_pe_1_5_0_n112, npu_inst_pe_1_5_0_n111,
         npu_inst_pe_1_5_0_n110, npu_inst_pe_1_5_0_n109,
         npu_inst_pe_1_5_0_n108, npu_inst_pe_1_5_0_n107,
         npu_inst_pe_1_5_0_n106, npu_inst_pe_1_5_0_n105,
         npu_inst_pe_1_5_0_n104, npu_inst_pe_1_5_0_n103,
         npu_inst_pe_1_5_0_n102, npu_inst_pe_1_5_0_n101,
         npu_inst_pe_1_5_0_n100, npu_inst_pe_1_5_0_n99, npu_inst_pe_1_5_0_n98,
         npu_inst_pe_1_5_0_n36, npu_inst_pe_1_5_0_n35, npu_inst_pe_1_5_0_n34,
         npu_inst_pe_1_5_0_n33, npu_inst_pe_1_5_0_n32, npu_inst_pe_1_5_0_n31,
         npu_inst_pe_1_5_0_n30, npu_inst_pe_1_5_0_n29, npu_inst_pe_1_5_0_n28,
         npu_inst_pe_1_5_0_n25, npu_inst_pe_1_5_0_n24, npu_inst_pe_1_5_0_n23,
         npu_inst_pe_1_5_0_n22, npu_inst_pe_1_5_0_n21, npu_inst_pe_1_5_0_n20,
         npu_inst_pe_1_5_0_n19, npu_inst_pe_1_5_0_n18, npu_inst_pe_1_5_0_n17,
         npu_inst_pe_1_5_0_n16, npu_inst_pe_1_5_0_n15, npu_inst_pe_1_5_0_n14,
         npu_inst_pe_1_5_0_n13, npu_inst_pe_1_5_0_n12, npu_inst_pe_1_5_0_n11,
         npu_inst_pe_1_5_0_n10, npu_inst_pe_1_5_0_n9, npu_inst_pe_1_5_0_n8,
         npu_inst_pe_1_5_0_n7, npu_inst_pe_1_5_0_n6, npu_inst_pe_1_5_0_n5,
         npu_inst_pe_1_5_0_n4, npu_inst_pe_1_5_0_n3, npu_inst_pe_1_5_0_n2,
         npu_inst_pe_1_5_0_n1, npu_inst_pe_1_5_0_sub_77_carry_7_,
         npu_inst_pe_1_5_0_sub_77_carry_6_, npu_inst_pe_1_5_0_sub_77_carry_5_,
         npu_inst_pe_1_5_0_sub_77_carry_4_, npu_inst_pe_1_5_0_sub_77_carry_3_,
         npu_inst_pe_1_5_0_sub_77_carry_2_, npu_inst_pe_1_5_0_sub_77_carry_1_,
         npu_inst_pe_1_5_0_add_79_carry_7_, npu_inst_pe_1_5_0_add_79_carry_6_,
         npu_inst_pe_1_5_0_add_79_carry_5_, npu_inst_pe_1_5_0_add_79_carry_4_,
         npu_inst_pe_1_5_0_add_79_carry_3_, npu_inst_pe_1_5_0_add_79_carry_2_,
         npu_inst_pe_1_5_0_add_79_carry_1_, npu_inst_pe_1_5_0_n97,
         npu_inst_pe_1_5_0_n96, npu_inst_pe_1_5_0_n95, npu_inst_pe_1_5_0_n94,
         npu_inst_pe_1_5_0_n93, npu_inst_pe_1_5_0_n92, npu_inst_pe_1_5_0_n91,
         npu_inst_pe_1_5_0_n90, npu_inst_pe_1_5_0_n89, npu_inst_pe_1_5_0_n88,
         npu_inst_pe_1_5_0_n87, npu_inst_pe_1_5_0_n86, npu_inst_pe_1_5_0_n85,
         npu_inst_pe_1_5_0_n84, npu_inst_pe_1_5_0_n83, npu_inst_pe_1_5_0_n82,
         npu_inst_pe_1_5_0_n81, npu_inst_pe_1_5_0_n80, npu_inst_pe_1_5_0_n79,
         npu_inst_pe_1_5_0_n78, npu_inst_pe_1_5_0_n77, npu_inst_pe_1_5_0_n76,
         npu_inst_pe_1_5_0_n75, npu_inst_pe_1_5_0_n74, npu_inst_pe_1_5_0_n73,
         npu_inst_pe_1_5_0_n72, npu_inst_pe_1_5_0_n71, npu_inst_pe_1_5_0_n70,
         npu_inst_pe_1_5_0_n69, npu_inst_pe_1_5_0_n68, npu_inst_pe_1_5_0_n67,
         npu_inst_pe_1_5_0_n66, npu_inst_pe_1_5_0_n65, npu_inst_pe_1_5_0_n64,
         npu_inst_pe_1_5_0_n63, npu_inst_pe_1_5_0_n62, npu_inst_pe_1_5_0_n61,
         npu_inst_pe_1_5_0_n60, npu_inst_pe_1_5_0_n59, npu_inst_pe_1_5_0_n58,
         npu_inst_pe_1_5_0_n57, npu_inst_pe_1_5_0_n56, npu_inst_pe_1_5_0_n55,
         npu_inst_pe_1_5_0_n54, npu_inst_pe_1_5_0_n53, npu_inst_pe_1_5_0_n52,
         npu_inst_pe_1_5_0_n51, npu_inst_pe_1_5_0_n50, npu_inst_pe_1_5_0_n49,
         npu_inst_pe_1_5_0_n48, npu_inst_pe_1_5_0_n47, npu_inst_pe_1_5_0_n46,
         npu_inst_pe_1_5_0_n45, npu_inst_pe_1_5_0_n44, npu_inst_pe_1_5_0_n43,
         npu_inst_pe_1_5_0_n42, npu_inst_pe_1_5_0_n41, npu_inst_pe_1_5_0_n40,
         npu_inst_pe_1_5_0_n39, npu_inst_pe_1_5_0_n38, npu_inst_pe_1_5_0_n37,
         npu_inst_pe_1_5_0_n27, npu_inst_pe_1_5_0_n26,
         npu_inst_pe_1_5_0_net3564, npu_inst_pe_1_5_0_net3558,
         npu_inst_pe_1_5_0_N94, npu_inst_pe_1_5_0_N93, npu_inst_pe_1_5_0_N84,
         npu_inst_pe_1_5_0_N80, npu_inst_pe_1_5_0_N79, npu_inst_pe_1_5_0_N78,
         npu_inst_pe_1_5_0_N77, npu_inst_pe_1_5_0_N76, npu_inst_pe_1_5_0_N75,
         npu_inst_pe_1_5_0_N74, npu_inst_pe_1_5_0_N73, npu_inst_pe_1_5_0_N72,
         npu_inst_pe_1_5_0_N71, npu_inst_pe_1_5_0_N70, npu_inst_pe_1_5_0_N69,
         npu_inst_pe_1_5_0_N68, npu_inst_pe_1_5_0_N67, npu_inst_pe_1_5_0_N66,
         npu_inst_pe_1_5_0_N65, npu_inst_pe_1_5_0_int_data_0_,
         npu_inst_pe_1_5_0_int_data_1_, npu_inst_pe_1_5_0_int_q_weight_0_,
         npu_inst_pe_1_5_0_int_q_weight_1_,
         npu_inst_pe_1_5_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_0_int_q_reg_h_0__1_, npu_inst_pe_1_5_0_o_data_h_0_,
         npu_inst_pe_1_5_0_o_data_h_1_, npu_inst_pe_1_5_1_n118,
         npu_inst_pe_1_5_1_n117, npu_inst_pe_1_5_1_n116,
         npu_inst_pe_1_5_1_n115, npu_inst_pe_1_5_1_n114,
         npu_inst_pe_1_5_1_n113, npu_inst_pe_1_5_1_n112,
         npu_inst_pe_1_5_1_n111, npu_inst_pe_1_5_1_n110,
         npu_inst_pe_1_5_1_n109, npu_inst_pe_1_5_1_n108,
         npu_inst_pe_1_5_1_n107, npu_inst_pe_1_5_1_n106,
         npu_inst_pe_1_5_1_n105, npu_inst_pe_1_5_1_n104,
         npu_inst_pe_1_5_1_n103, npu_inst_pe_1_5_1_n102,
         npu_inst_pe_1_5_1_n101, npu_inst_pe_1_5_1_n100, npu_inst_pe_1_5_1_n99,
         npu_inst_pe_1_5_1_n98, npu_inst_pe_1_5_1_n36, npu_inst_pe_1_5_1_n35,
         npu_inst_pe_1_5_1_n34, npu_inst_pe_1_5_1_n33, npu_inst_pe_1_5_1_n32,
         npu_inst_pe_1_5_1_n31, npu_inst_pe_1_5_1_n30, npu_inst_pe_1_5_1_n29,
         npu_inst_pe_1_5_1_n28, npu_inst_pe_1_5_1_n25, npu_inst_pe_1_5_1_n24,
         npu_inst_pe_1_5_1_n23, npu_inst_pe_1_5_1_n22, npu_inst_pe_1_5_1_n21,
         npu_inst_pe_1_5_1_n20, npu_inst_pe_1_5_1_n19, npu_inst_pe_1_5_1_n18,
         npu_inst_pe_1_5_1_n17, npu_inst_pe_1_5_1_n16, npu_inst_pe_1_5_1_n15,
         npu_inst_pe_1_5_1_n14, npu_inst_pe_1_5_1_n13, npu_inst_pe_1_5_1_n12,
         npu_inst_pe_1_5_1_n11, npu_inst_pe_1_5_1_n10, npu_inst_pe_1_5_1_n9,
         npu_inst_pe_1_5_1_n8, npu_inst_pe_1_5_1_n7, npu_inst_pe_1_5_1_n6,
         npu_inst_pe_1_5_1_n5, npu_inst_pe_1_5_1_n4, npu_inst_pe_1_5_1_n3,
         npu_inst_pe_1_5_1_n2, npu_inst_pe_1_5_1_n1,
         npu_inst_pe_1_5_1_sub_77_carry_7_, npu_inst_pe_1_5_1_sub_77_carry_6_,
         npu_inst_pe_1_5_1_sub_77_carry_5_, npu_inst_pe_1_5_1_sub_77_carry_4_,
         npu_inst_pe_1_5_1_sub_77_carry_3_, npu_inst_pe_1_5_1_sub_77_carry_2_,
         npu_inst_pe_1_5_1_sub_77_carry_1_, npu_inst_pe_1_5_1_add_79_carry_7_,
         npu_inst_pe_1_5_1_add_79_carry_6_, npu_inst_pe_1_5_1_add_79_carry_5_,
         npu_inst_pe_1_5_1_add_79_carry_4_, npu_inst_pe_1_5_1_add_79_carry_3_,
         npu_inst_pe_1_5_1_add_79_carry_2_, npu_inst_pe_1_5_1_add_79_carry_1_,
         npu_inst_pe_1_5_1_n97, npu_inst_pe_1_5_1_n96, npu_inst_pe_1_5_1_n95,
         npu_inst_pe_1_5_1_n94, npu_inst_pe_1_5_1_n93, npu_inst_pe_1_5_1_n92,
         npu_inst_pe_1_5_1_n91, npu_inst_pe_1_5_1_n90, npu_inst_pe_1_5_1_n89,
         npu_inst_pe_1_5_1_n88, npu_inst_pe_1_5_1_n87, npu_inst_pe_1_5_1_n86,
         npu_inst_pe_1_5_1_n85, npu_inst_pe_1_5_1_n84, npu_inst_pe_1_5_1_n83,
         npu_inst_pe_1_5_1_n82, npu_inst_pe_1_5_1_n81, npu_inst_pe_1_5_1_n80,
         npu_inst_pe_1_5_1_n79, npu_inst_pe_1_5_1_n78, npu_inst_pe_1_5_1_n77,
         npu_inst_pe_1_5_1_n76, npu_inst_pe_1_5_1_n75, npu_inst_pe_1_5_1_n74,
         npu_inst_pe_1_5_1_n73, npu_inst_pe_1_5_1_n72, npu_inst_pe_1_5_1_n71,
         npu_inst_pe_1_5_1_n70, npu_inst_pe_1_5_1_n69, npu_inst_pe_1_5_1_n68,
         npu_inst_pe_1_5_1_n67, npu_inst_pe_1_5_1_n66, npu_inst_pe_1_5_1_n65,
         npu_inst_pe_1_5_1_n64, npu_inst_pe_1_5_1_n63, npu_inst_pe_1_5_1_n62,
         npu_inst_pe_1_5_1_n61, npu_inst_pe_1_5_1_n60, npu_inst_pe_1_5_1_n59,
         npu_inst_pe_1_5_1_n58, npu_inst_pe_1_5_1_n57, npu_inst_pe_1_5_1_n56,
         npu_inst_pe_1_5_1_n55, npu_inst_pe_1_5_1_n54, npu_inst_pe_1_5_1_n53,
         npu_inst_pe_1_5_1_n52, npu_inst_pe_1_5_1_n51, npu_inst_pe_1_5_1_n50,
         npu_inst_pe_1_5_1_n49, npu_inst_pe_1_5_1_n48, npu_inst_pe_1_5_1_n47,
         npu_inst_pe_1_5_1_n46, npu_inst_pe_1_5_1_n45, npu_inst_pe_1_5_1_n44,
         npu_inst_pe_1_5_1_n43, npu_inst_pe_1_5_1_n42, npu_inst_pe_1_5_1_n41,
         npu_inst_pe_1_5_1_n40, npu_inst_pe_1_5_1_n39, npu_inst_pe_1_5_1_n38,
         npu_inst_pe_1_5_1_n37, npu_inst_pe_1_5_1_n27, npu_inst_pe_1_5_1_n26,
         npu_inst_pe_1_5_1_net3541, npu_inst_pe_1_5_1_net3535,
         npu_inst_pe_1_5_1_N94, npu_inst_pe_1_5_1_N93, npu_inst_pe_1_5_1_N84,
         npu_inst_pe_1_5_1_N80, npu_inst_pe_1_5_1_N79, npu_inst_pe_1_5_1_N78,
         npu_inst_pe_1_5_1_N77, npu_inst_pe_1_5_1_N76, npu_inst_pe_1_5_1_N75,
         npu_inst_pe_1_5_1_N74, npu_inst_pe_1_5_1_N73, npu_inst_pe_1_5_1_N72,
         npu_inst_pe_1_5_1_N71, npu_inst_pe_1_5_1_N70, npu_inst_pe_1_5_1_N69,
         npu_inst_pe_1_5_1_N68, npu_inst_pe_1_5_1_N67, npu_inst_pe_1_5_1_N66,
         npu_inst_pe_1_5_1_N65, npu_inst_pe_1_5_1_int_data_0_,
         npu_inst_pe_1_5_1_int_data_1_, npu_inst_pe_1_5_1_int_q_weight_0_,
         npu_inst_pe_1_5_1_int_q_weight_1_,
         npu_inst_pe_1_5_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_1_int_q_reg_h_0__1_, npu_inst_pe_1_5_2_n118,
         npu_inst_pe_1_5_2_n117, npu_inst_pe_1_5_2_n116,
         npu_inst_pe_1_5_2_n115, npu_inst_pe_1_5_2_n114,
         npu_inst_pe_1_5_2_n113, npu_inst_pe_1_5_2_n112,
         npu_inst_pe_1_5_2_n111, npu_inst_pe_1_5_2_n110,
         npu_inst_pe_1_5_2_n109, npu_inst_pe_1_5_2_n108,
         npu_inst_pe_1_5_2_n107, npu_inst_pe_1_5_2_n106,
         npu_inst_pe_1_5_2_n105, npu_inst_pe_1_5_2_n104,
         npu_inst_pe_1_5_2_n103, npu_inst_pe_1_5_2_n102,
         npu_inst_pe_1_5_2_n101, npu_inst_pe_1_5_2_n100, npu_inst_pe_1_5_2_n99,
         npu_inst_pe_1_5_2_n98, npu_inst_pe_1_5_2_n36, npu_inst_pe_1_5_2_n35,
         npu_inst_pe_1_5_2_n34, npu_inst_pe_1_5_2_n33, npu_inst_pe_1_5_2_n32,
         npu_inst_pe_1_5_2_n31, npu_inst_pe_1_5_2_n30, npu_inst_pe_1_5_2_n29,
         npu_inst_pe_1_5_2_n28, npu_inst_pe_1_5_2_n25, npu_inst_pe_1_5_2_n24,
         npu_inst_pe_1_5_2_n23, npu_inst_pe_1_5_2_n22, npu_inst_pe_1_5_2_n21,
         npu_inst_pe_1_5_2_n20, npu_inst_pe_1_5_2_n19, npu_inst_pe_1_5_2_n18,
         npu_inst_pe_1_5_2_n17, npu_inst_pe_1_5_2_n16, npu_inst_pe_1_5_2_n15,
         npu_inst_pe_1_5_2_n14, npu_inst_pe_1_5_2_n13, npu_inst_pe_1_5_2_n12,
         npu_inst_pe_1_5_2_n11, npu_inst_pe_1_5_2_n10, npu_inst_pe_1_5_2_n9,
         npu_inst_pe_1_5_2_n8, npu_inst_pe_1_5_2_n7, npu_inst_pe_1_5_2_n6,
         npu_inst_pe_1_5_2_n5, npu_inst_pe_1_5_2_n4, npu_inst_pe_1_5_2_n3,
         npu_inst_pe_1_5_2_n2, npu_inst_pe_1_5_2_n1,
         npu_inst_pe_1_5_2_sub_77_carry_7_, npu_inst_pe_1_5_2_sub_77_carry_6_,
         npu_inst_pe_1_5_2_sub_77_carry_5_, npu_inst_pe_1_5_2_sub_77_carry_4_,
         npu_inst_pe_1_5_2_sub_77_carry_3_, npu_inst_pe_1_5_2_sub_77_carry_2_,
         npu_inst_pe_1_5_2_sub_77_carry_1_, npu_inst_pe_1_5_2_add_79_carry_7_,
         npu_inst_pe_1_5_2_add_79_carry_6_, npu_inst_pe_1_5_2_add_79_carry_5_,
         npu_inst_pe_1_5_2_add_79_carry_4_, npu_inst_pe_1_5_2_add_79_carry_3_,
         npu_inst_pe_1_5_2_add_79_carry_2_, npu_inst_pe_1_5_2_add_79_carry_1_,
         npu_inst_pe_1_5_2_n97, npu_inst_pe_1_5_2_n96, npu_inst_pe_1_5_2_n95,
         npu_inst_pe_1_5_2_n94, npu_inst_pe_1_5_2_n93, npu_inst_pe_1_5_2_n92,
         npu_inst_pe_1_5_2_n91, npu_inst_pe_1_5_2_n90, npu_inst_pe_1_5_2_n89,
         npu_inst_pe_1_5_2_n88, npu_inst_pe_1_5_2_n87, npu_inst_pe_1_5_2_n86,
         npu_inst_pe_1_5_2_n85, npu_inst_pe_1_5_2_n84, npu_inst_pe_1_5_2_n83,
         npu_inst_pe_1_5_2_n82, npu_inst_pe_1_5_2_n81, npu_inst_pe_1_5_2_n80,
         npu_inst_pe_1_5_2_n79, npu_inst_pe_1_5_2_n78, npu_inst_pe_1_5_2_n77,
         npu_inst_pe_1_5_2_n76, npu_inst_pe_1_5_2_n75, npu_inst_pe_1_5_2_n74,
         npu_inst_pe_1_5_2_n73, npu_inst_pe_1_5_2_n72, npu_inst_pe_1_5_2_n71,
         npu_inst_pe_1_5_2_n70, npu_inst_pe_1_5_2_n69, npu_inst_pe_1_5_2_n68,
         npu_inst_pe_1_5_2_n67, npu_inst_pe_1_5_2_n66, npu_inst_pe_1_5_2_n65,
         npu_inst_pe_1_5_2_n64, npu_inst_pe_1_5_2_n63, npu_inst_pe_1_5_2_n62,
         npu_inst_pe_1_5_2_n61, npu_inst_pe_1_5_2_n60, npu_inst_pe_1_5_2_n59,
         npu_inst_pe_1_5_2_n58, npu_inst_pe_1_5_2_n57, npu_inst_pe_1_5_2_n56,
         npu_inst_pe_1_5_2_n55, npu_inst_pe_1_5_2_n54, npu_inst_pe_1_5_2_n53,
         npu_inst_pe_1_5_2_n52, npu_inst_pe_1_5_2_n51, npu_inst_pe_1_5_2_n50,
         npu_inst_pe_1_5_2_n49, npu_inst_pe_1_5_2_n48, npu_inst_pe_1_5_2_n47,
         npu_inst_pe_1_5_2_n46, npu_inst_pe_1_5_2_n45, npu_inst_pe_1_5_2_n44,
         npu_inst_pe_1_5_2_n43, npu_inst_pe_1_5_2_n42, npu_inst_pe_1_5_2_n41,
         npu_inst_pe_1_5_2_n40, npu_inst_pe_1_5_2_n39, npu_inst_pe_1_5_2_n38,
         npu_inst_pe_1_5_2_n37, npu_inst_pe_1_5_2_n27, npu_inst_pe_1_5_2_n26,
         npu_inst_pe_1_5_2_net3518, npu_inst_pe_1_5_2_net3512,
         npu_inst_pe_1_5_2_N94, npu_inst_pe_1_5_2_N93, npu_inst_pe_1_5_2_N84,
         npu_inst_pe_1_5_2_N80, npu_inst_pe_1_5_2_N79, npu_inst_pe_1_5_2_N78,
         npu_inst_pe_1_5_2_N77, npu_inst_pe_1_5_2_N76, npu_inst_pe_1_5_2_N75,
         npu_inst_pe_1_5_2_N74, npu_inst_pe_1_5_2_N73, npu_inst_pe_1_5_2_N72,
         npu_inst_pe_1_5_2_N71, npu_inst_pe_1_5_2_N70, npu_inst_pe_1_5_2_N69,
         npu_inst_pe_1_5_2_N68, npu_inst_pe_1_5_2_N67, npu_inst_pe_1_5_2_N66,
         npu_inst_pe_1_5_2_N65, npu_inst_pe_1_5_2_int_data_0_,
         npu_inst_pe_1_5_2_int_data_1_, npu_inst_pe_1_5_2_int_q_weight_0_,
         npu_inst_pe_1_5_2_int_q_weight_1_,
         npu_inst_pe_1_5_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_2_int_q_reg_h_0__1_, npu_inst_pe_1_5_3_n118,
         npu_inst_pe_1_5_3_n117, npu_inst_pe_1_5_3_n116,
         npu_inst_pe_1_5_3_n115, npu_inst_pe_1_5_3_n114,
         npu_inst_pe_1_5_3_n113, npu_inst_pe_1_5_3_n112,
         npu_inst_pe_1_5_3_n111, npu_inst_pe_1_5_3_n110,
         npu_inst_pe_1_5_3_n109, npu_inst_pe_1_5_3_n108,
         npu_inst_pe_1_5_3_n107, npu_inst_pe_1_5_3_n106,
         npu_inst_pe_1_5_3_n105, npu_inst_pe_1_5_3_n104,
         npu_inst_pe_1_5_3_n103, npu_inst_pe_1_5_3_n102,
         npu_inst_pe_1_5_3_n101, npu_inst_pe_1_5_3_n100, npu_inst_pe_1_5_3_n99,
         npu_inst_pe_1_5_3_n98, npu_inst_pe_1_5_3_n36, npu_inst_pe_1_5_3_n35,
         npu_inst_pe_1_5_3_n34, npu_inst_pe_1_5_3_n33, npu_inst_pe_1_5_3_n32,
         npu_inst_pe_1_5_3_n31, npu_inst_pe_1_5_3_n30, npu_inst_pe_1_5_3_n29,
         npu_inst_pe_1_5_3_n28, npu_inst_pe_1_5_3_n25, npu_inst_pe_1_5_3_n24,
         npu_inst_pe_1_5_3_n23, npu_inst_pe_1_5_3_n22, npu_inst_pe_1_5_3_n21,
         npu_inst_pe_1_5_3_n20, npu_inst_pe_1_5_3_n19, npu_inst_pe_1_5_3_n18,
         npu_inst_pe_1_5_3_n17, npu_inst_pe_1_5_3_n16, npu_inst_pe_1_5_3_n15,
         npu_inst_pe_1_5_3_n14, npu_inst_pe_1_5_3_n13, npu_inst_pe_1_5_3_n12,
         npu_inst_pe_1_5_3_n11, npu_inst_pe_1_5_3_n10, npu_inst_pe_1_5_3_n9,
         npu_inst_pe_1_5_3_n8, npu_inst_pe_1_5_3_n7, npu_inst_pe_1_5_3_n6,
         npu_inst_pe_1_5_3_n5, npu_inst_pe_1_5_3_n4, npu_inst_pe_1_5_3_n3,
         npu_inst_pe_1_5_3_n2, npu_inst_pe_1_5_3_n1,
         npu_inst_pe_1_5_3_sub_77_carry_7_, npu_inst_pe_1_5_3_sub_77_carry_6_,
         npu_inst_pe_1_5_3_sub_77_carry_5_, npu_inst_pe_1_5_3_sub_77_carry_4_,
         npu_inst_pe_1_5_3_sub_77_carry_3_, npu_inst_pe_1_5_3_sub_77_carry_2_,
         npu_inst_pe_1_5_3_sub_77_carry_1_, npu_inst_pe_1_5_3_add_79_carry_7_,
         npu_inst_pe_1_5_3_add_79_carry_6_, npu_inst_pe_1_5_3_add_79_carry_5_,
         npu_inst_pe_1_5_3_add_79_carry_4_, npu_inst_pe_1_5_3_add_79_carry_3_,
         npu_inst_pe_1_5_3_add_79_carry_2_, npu_inst_pe_1_5_3_add_79_carry_1_,
         npu_inst_pe_1_5_3_n97, npu_inst_pe_1_5_3_n96, npu_inst_pe_1_5_3_n95,
         npu_inst_pe_1_5_3_n94, npu_inst_pe_1_5_3_n93, npu_inst_pe_1_5_3_n92,
         npu_inst_pe_1_5_3_n91, npu_inst_pe_1_5_3_n90, npu_inst_pe_1_5_3_n89,
         npu_inst_pe_1_5_3_n88, npu_inst_pe_1_5_3_n87, npu_inst_pe_1_5_3_n86,
         npu_inst_pe_1_5_3_n85, npu_inst_pe_1_5_3_n84, npu_inst_pe_1_5_3_n83,
         npu_inst_pe_1_5_3_n82, npu_inst_pe_1_5_3_n81, npu_inst_pe_1_5_3_n80,
         npu_inst_pe_1_5_3_n79, npu_inst_pe_1_5_3_n78, npu_inst_pe_1_5_3_n77,
         npu_inst_pe_1_5_3_n76, npu_inst_pe_1_5_3_n75, npu_inst_pe_1_5_3_n74,
         npu_inst_pe_1_5_3_n73, npu_inst_pe_1_5_3_n72, npu_inst_pe_1_5_3_n71,
         npu_inst_pe_1_5_3_n70, npu_inst_pe_1_5_3_n69, npu_inst_pe_1_5_3_n68,
         npu_inst_pe_1_5_3_n67, npu_inst_pe_1_5_3_n66, npu_inst_pe_1_5_3_n65,
         npu_inst_pe_1_5_3_n64, npu_inst_pe_1_5_3_n63, npu_inst_pe_1_5_3_n62,
         npu_inst_pe_1_5_3_n61, npu_inst_pe_1_5_3_n60, npu_inst_pe_1_5_3_n59,
         npu_inst_pe_1_5_3_n58, npu_inst_pe_1_5_3_n57, npu_inst_pe_1_5_3_n56,
         npu_inst_pe_1_5_3_n55, npu_inst_pe_1_5_3_n54, npu_inst_pe_1_5_3_n53,
         npu_inst_pe_1_5_3_n52, npu_inst_pe_1_5_3_n51, npu_inst_pe_1_5_3_n50,
         npu_inst_pe_1_5_3_n49, npu_inst_pe_1_5_3_n48, npu_inst_pe_1_5_3_n47,
         npu_inst_pe_1_5_3_n46, npu_inst_pe_1_5_3_n45, npu_inst_pe_1_5_3_n44,
         npu_inst_pe_1_5_3_n43, npu_inst_pe_1_5_3_n42, npu_inst_pe_1_5_3_n41,
         npu_inst_pe_1_5_3_n40, npu_inst_pe_1_5_3_n39, npu_inst_pe_1_5_3_n38,
         npu_inst_pe_1_5_3_n37, npu_inst_pe_1_5_3_n27, npu_inst_pe_1_5_3_n26,
         npu_inst_pe_1_5_3_net3495, npu_inst_pe_1_5_3_net3489,
         npu_inst_pe_1_5_3_N94, npu_inst_pe_1_5_3_N93, npu_inst_pe_1_5_3_N84,
         npu_inst_pe_1_5_3_N80, npu_inst_pe_1_5_3_N79, npu_inst_pe_1_5_3_N78,
         npu_inst_pe_1_5_3_N77, npu_inst_pe_1_5_3_N76, npu_inst_pe_1_5_3_N75,
         npu_inst_pe_1_5_3_N74, npu_inst_pe_1_5_3_N73, npu_inst_pe_1_5_3_N72,
         npu_inst_pe_1_5_3_N71, npu_inst_pe_1_5_3_N70, npu_inst_pe_1_5_3_N69,
         npu_inst_pe_1_5_3_N68, npu_inst_pe_1_5_3_N67, npu_inst_pe_1_5_3_N66,
         npu_inst_pe_1_5_3_N65, npu_inst_pe_1_5_3_int_data_0_,
         npu_inst_pe_1_5_3_int_data_1_, npu_inst_pe_1_5_3_int_q_weight_0_,
         npu_inst_pe_1_5_3_int_q_weight_1_,
         npu_inst_pe_1_5_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_3_int_q_reg_h_0__1_, npu_inst_pe_1_5_4_n118,
         npu_inst_pe_1_5_4_n117, npu_inst_pe_1_5_4_n116,
         npu_inst_pe_1_5_4_n115, npu_inst_pe_1_5_4_n114,
         npu_inst_pe_1_5_4_n113, npu_inst_pe_1_5_4_n112,
         npu_inst_pe_1_5_4_n111, npu_inst_pe_1_5_4_n110,
         npu_inst_pe_1_5_4_n109, npu_inst_pe_1_5_4_n108,
         npu_inst_pe_1_5_4_n107, npu_inst_pe_1_5_4_n106,
         npu_inst_pe_1_5_4_n105, npu_inst_pe_1_5_4_n104,
         npu_inst_pe_1_5_4_n103, npu_inst_pe_1_5_4_n102,
         npu_inst_pe_1_5_4_n101, npu_inst_pe_1_5_4_n100, npu_inst_pe_1_5_4_n99,
         npu_inst_pe_1_5_4_n98, npu_inst_pe_1_5_4_n36, npu_inst_pe_1_5_4_n35,
         npu_inst_pe_1_5_4_n34, npu_inst_pe_1_5_4_n33, npu_inst_pe_1_5_4_n32,
         npu_inst_pe_1_5_4_n31, npu_inst_pe_1_5_4_n30, npu_inst_pe_1_5_4_n29,
         npu_inst_pe_1_5_4_n28, npu_inst_pe_1_5_4_n25, npu_inst_pe_1_5_4_n24,
         npu_inst_pe_1_5_4_n23, npu_inst_pe_1_5_4_n22, npu_inst_pe_1_5_4_n21,
         npu_inst_pe_1_5_4_n20, npu_inst_pe_1_5_4_n19, npu_inst_pe_1_5_4_n18,
         npu_inst_pe_1_5_4_n17, npu_inst_pe_1_5_4_n16, npu_inst_pe_1_5_4_n15,
         npu_inst_pe_1_5_4_n14, npu_inst_pe_1_5_4_n13, npu_inst_pe_1_5_4_n12,
         npu_inst_pe_1_5_4_n11, npu_inst_pe_1_5_4_n10, npu_inst_pe_1_5_4_n9,
         npu_inst_pe_1_5_4_n8, npu_inst_pe_1_5_4_n7, npu_inst_pe_1_5_4_n6,
         npu_inst_pe_1_5_4_n5, npu_inst_pe_1_5_4_n4, npu_inst_pe_1_5_4_n3,
         npu_inst_pe_1_5_4_n2, npu_inst_pe_1_5_4_n1,
         npu_inst_pe_1_5_4_sub_77_carry_7_, npu_inst_pe_1_5_4_sub_77_carry_6_,
         npu_inst_pe_1_5_4_sub_77_carry_5_, npu_inst_pe_1_5_4_sub_77_carry_4_,
         npu_inst_pe_1_5_4_sub_77_carry_3_, npu_inst_pe_1_5_4_sub_77_carry_2_,
         npu_inst_pe_1_5_4_sub_77_carry_1_, npu_inst_pe_1_5_4_add_79_carry_7_,
         npu_inst_pe_1_5_4_add_79_carry_6_, npu_inst_pe_1_5_4_add_79_carry_5_,
         npu_inst_pe_1_5_4_add_79_carry_4_, npu_inst_pe_1_5_4_add_79_carry_3_,
         npu_inst_pe_1_5_4_add_79_carry_2_, npu_inst_pe_1_5_4_add_79_carry_1_,
         npu_inst_pe_1_5_4_n97, npu_inst_pe_1_5_4_n96, npu_inst_pe_1_5_4_n95,
         npu_inst_pe_1_5_4_n94, npu_inst_pe_1_5_4_n93, npu_inst_pe_1_5_4_n92,
         npu_inst_pe_1_5_4_n91, npu_inst_pe_1_5_4_n90, npu_inst_pe_1_5_4_n89,
         npu_inst_pe_1_5_4_n88, npu_inst_pe_1_5_4_n87, npu_inst_pe_1_5_4_n86,
         npu_inst_pe_1_5_4_n85, npu_inst_pe_1_5_4_n84, npu_inst_pe_1_5_4_n83,
         npu_inst_pe_1_5_4_n82, npu_inst_pe_1_5_4_n81, npu_inst_pe_1_5_4_n80,
         npu_inst_pe_1_5_4_n79, npu_inst_pe_1_5_4_n78, npu_inst_pe_1_5_4_n77,
         npu_inst_pe_1_5_4_n76, npu_inst_pe_1_5_4_n75, npu_inst_pe_1_5_4_n74,
         npu_inst_pe_1_5_4_n73, npu_inst_pe_1_5_4_n72, npu_inst_pe_1_5_4_n71,
         npu_inst_pe_1_5_4_n70, npu_inst_pe_1_5_4_n69, npu_inst_pe_1_5_4_n68,
         npu_inst_pe_1_5_4_n67, npu_inst_pe_1_5_4_n66, npu_inst_pe_1_5_4_n65,
         npu_inst_pe_1_5_4_n64, npu_inst_pe_1_5_4_n63, npu_inst_pe_1_5_4_n62,
         npu_inst_pe_1_5_4_n61, npu_inst_pe_1_5_4_n60, npu_inst_pe_1_5_4_n59,
         npu_inst_pe_1_5_4_n58, npu_inst_pe_1_5_4_n57, npu_inst_pe_1_5_4_n56,
         npu_inst_pe_1_5_4_n55, npu_inst_pe_1_5_4_n54, npu_inst_pe_1_5_4_n53,
         npu_inst_pe_1_5_4_n52, npu_inst_pe_1_5_4_n51, npu_inst_pe_1_5_4_n50,
         npu_inst_pe_1_5_4_n49, npu_inst_pe_1_5_4_n48, npu_inst_pe_1_5_4_n47,
         npu_inst_pe_1_5_4_n46, npu_inst_pe_1_5_4_n45, npu_inst_pe_1_5_4_n44,
         npu_inst_pe_1_5_4_n43, npu_inst_pe_1_5_4_n42, npu_inst_pe_1_5_4_n41,
         npu_inst_pe_1_5_4_n40, npu_inst_pe_1_5_4_n39, npu_inst_pe_1_5_4_n38,
         npu_inst_pe_1_5_4_n37, npu_inst_pe_1_5_4_n27, npu_inst_pe_1_5_4_n26,
         npu_inst_pe_1_5_4_net3472, npu_inst_pe_1_5_4_net3466,
         npu_inst_pe_1_5_4_N94, npu_inst_pe_1_5_4_N93, npu_inst_pe_1_5_4_N84,
         npu_inst_pe_1_5_4_N80, npu_inst_pe_1_5_4_N79, npu_inst_pe_1_5_4_N78,
         npu_inst_pe_1_5_4_N77, npu_inst_pe_1_5_4_N76, npu_inst_pe_1_5_4_N75,
         npu_inst_pe_1_5_4_N74, npu_inst_pe_1_5_4_N73, npu_inst_pe_1_5_4_N72,
         npu_inst_pe_1_5_4_N71, npu_inst_pe_1_5_4_N70, npu_inst_pe_1_5_4_N69,
         npu_inst_pe_1_5_4_N68, npu_inst_pe_1_5_4_N67, npu_inst_pe_1_5_4_N66,
         npu_inst_pe_1_5_4_N65, npu_inst_pe_1_5_4_int_data_0_,
         npu_inst_pe_1_5_4_int_data_1_, npu_inst_pe_1_5_4_int_q_weight_0_,
         npu_inst_pe_1_5_4_int_q_weight_1_,
         npu_inst_pe_1_5_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_4_int_q_reg_h_0__1_, npu_inst_pe_1_5_5_n118,
         npu_inst_pe_1_5_5_n117, npu_inst_pe_1_5_5_n116,
         npu_inst_pe_1_5_5_n115, npu_inst_pe_1_5_5_n114,
         npu_inst_pe_1_5_5_n113, npu_inst_pe_1_5_5_n112,
         npu_inst_pe_1_5_5_n111, npu_inst_pe_1_5_5_n110,
         npu_inst_pe_1_5_5_n109, npu_inst_pe_1_5_5_n108,
         npu_inst_pe_1_5_5_n107, npu_inst_pe_1_5_5_n106,
         npu_inst_pe_1_5_5_n105, npu_inst_pe_1_5_5_n104,
         npu_inst_pe_1_5_5_n103, npu_inst_pe_1_5_5_n102,
         npu_inst_pe_1_5_5_n101, npu_inst_pe_1_5_5_n100, npu_inst_pe_1_5_5_n99,
         npu_inst_pe_1_5_5_n98, npu_inst_pe_1_5_5_n36, npu_inst_pe_1_5_5_n35,
         npu_inst_pe_1_5_5_n34, npu_inst_pe_1_5_5_n33, npu_inst_pe_1_5_5_n32,
         npu_inst_pe_1_5_5_n31, npu_inst_pe_1_5_5_n30, npu_inst_pe_1_5_5_n29,
         npu_inst_pe_1_5_5_n28, npu_inst_pe_1_5_5_n25, npu_inst_pe_1_5_5_n24,
         npu_inst_pe_1_5_5_n23, npu_inst_pe_1_5_5_n22, npu_inst_pe_1_5_5_n21,
         npu_inst_pe_1_5_5_n20, npu_inst_pe_1_5_5_n19, npu_inst_pe_1_5_5_n18,
         npu_inst_pe_1_5_5_n17, npu_inst_pe_1_5_5_n16, npu_inst_pe_1_5_5_n15,
         npu_inst_pe_1_5_5_n14, npu_inst_pe_1_5_5_n13, npu_inst_pe_1_5_5_n12,
         npu_inst_pe_1_5_5_n11, npu_inst_pe_1_5_5_n10, npu_inst_pe_1_5_5_n9,
         npu_inst_pe_1_5_5_n8, npu_inst_pe_1_5_5_n7, npu_inst_pe_1_5_5_n6,
         npu_inst_pe_1_5_5_n5, npu_inst_pe_1_5_5_n4, npu_inst_pe_1_5_5_n3,
         npu_inst_pe_1_5_5_n2, npu_inst_pe_1_5_5_n1,
         npu_inst_pe_1_5_5_sub_77_carry_7_, npu_inst_pe_1_5_5_sub_77_carry_6_,
         npu_inst_pe_1_5_5_sub_77_carry_5_, npu_inst_pe_1_5_5_sub_77_carry_4_,
         npu_inst_pe_1_5_5_sub_77_carry_3_, npu_inst_pe_1_5_5_sub_77_carry_2_,
         npu_inst_pe_1_5_5_sub_77_carry_1_, npu_inst_pe_1_5_5_add_79_carry_7_,
         npu_inst_pe_1_5_5_add_79_carry_6_, npu_inst_pe_1_5_5_add_79_carry_5_,
         npu_inst_pe_1_5_5_add_79_carry_4_, npu_inst_pe_1_5_5_add_79_carry_3_,
         npu_inst_pe_1_5_5_add_79_carry_2_, npu_inst_pe_1_5_5_add_79_carry_1_,
         npu_inst_pe_1_5_5_n97, npu_inst_pe_1_5_5_n96, npu_inst_pe_1_5_5_n95,
         npu_inst_pe_1_5_5_n94, npu_inst_pe_1_5_5_n93, npu_inst_pe_1_5_5_n92,
         npu_inst_pe_1_5_5_n91, npu_inst_pe_1_5_5_n90, npu_inst_pe_1_5_5_n89,
         npu_inst_pe_1_5_5_n88, npu_inst_pe_1_5_5_n87, npu_inst_pe_1_5_5_n86,
         npu_inst_pe_1_5_5_n85, npu_inst_pe_1_5_5_n84, npu_inst_pe_1_5_5_n83,
         npu_inst_pe_1_5_5_n82, npu_inst_pe_1_5_5_n81, npu_inst_pe_1_5_5_n80,
         npu_inst_pe_1_5_5_n79, npu_inst_pe_1_5_5_n78, npu_inst_pe_1_5_5_n77,
         npu_inst_pe_1_5_5_n76, npu_inst_pe_1_5_5_n75, npu_inst_pe_1_5_5_n74,
         npu_inst_pe_1_5_5_n73, npu_inst_pe_1_5_5_n72, npu_inst_pe_1_5_5_n71,
         npu_inst_pe_1_5_5_n70, npu_inst_pe_1_5_5_n69, npu_inst_pe_1_5_5_n68,
         npu_inst_pe_1_5_5_n67, npu_inst_pe_1_5_5_n66, npu_inst_pe_1_5_5_n65,
         npu_inst_pe_1_5_5_n64, npu_inst_pe_1_5_5_n63, npu_inst_pe_1_5_5_n62,
         npu_inst_pe_1_5_5_n61, npu_inst_pe_1_5_5_n60, npu_inst_pe_1_5_5_n59,
         npu_inst_pe_1_5_5_n58, npu_inst_pe_1_5_5_n57, npu_inst_pe_1_5_5_n56,
         npu_inst_pe_1_5_5_n55, npu_inst_pe_1_5_5_n54, npu_inst_pe_1_5_5_n53,
         npu_inst_pe_1_5_5_n52, npu_inst_pe_1_5_5_n51, npu_inst_pe_1_5_5_n50,
         npu_inst_pe_1_5_5_n49, npu_inst_pe_1_5_5_n48, npu_inst_pe_1_5_5_n47,
         npu_inst_pe_1_5_5_n46, npu_inst_pe_1_5_5_n45, npu_inst_pe_1_5_5_n44,
         npu_inst_pe_1_5_5_n43, npu_inst_pe_1_5_5_n42, npu_inst_pe_1_5_5_n41,
         npu_inst_pe_1_5_5_n40, npu_inst_pe_1_5_5_n39, npu_inst_pe_1_5_5_n38,
         npu_inst_pe_1_5_5_n37, npu_inst_pe_1_5_5_n27, npu_inst_pe_1_5_5_n26,
         npu_inst_pe_1_5_5_net3449, npu_inst_pe_1_5_5_net3443,
         npu_inst_pe_1_5_5_N94, npu_inst_pe_1_5_5_N93, npu_inst_pe_1_5_5_N84,
         npu_inst_pe_1_5_5_N80, npu_inst_pe_1_5_5_N79, npu_inst_pe_1_5_5_N78,
         npu_inst_pe_1_5_5_N77, npu_inst_pe_1_5_5_N76, npu_inst_pe_1_5_5_N75,
         npu_inst_pe_1_5_5_N74, npu_inst_pe_1_5_5_N73, npu_inst_pe_1_5_5_N72,
         npu_inst_pe_1_5_5_N71, npu_inst_pe_1_5_5_N70, npu_inst_pe_1_5_5_N69,
         npu_inst_pe_1_5_5_N68, npu_inst_pe_1_5_5_N67, npu_inst_pe_1_5_5_N66,
         npu_inst_pe_1_5_5_N65, npu_inst_pe_1_5_5_int_data_0_,
         npu_inst_pe_1_5_5_int_data_1_, npu_inst_pe_1_5_5_int_q_weight_0_,
         npu_inst_pe_1_5_5_int_q_weight_1_,
         npu_inst_pe_1_5_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_5_int_q_reg_h_0__1_, npu_inst_pe_1_5_6_n118,
         npu_inst_pe_1_5_6_n117, npu_inst_pe_1_5_6_n116,
         npu_inst_pe_1_5_6_n115, npu_inst_pe_1_5_6_n114,
         npu_inst_pe_1_5_6_n113, npu_inst_pe_1_5_6_n112,
         npu_inst_pe_1_5_6_n111, npu_inst_pe_1_5_6_n110,
         npu_inst_pe_1_5_6_n109, npu_inst_pe_1_5_6_n108,
         npu_inst_pe_1_5_6_n107, npu_inst_pe_1_5_6_n106,
         npu_inst_pe_1_5_6_n105, npu_inst_pe_1_5_6_n104,
         npu_inst_pe_1_5_6_n103, npu_inst_pe_1_5_6_n102,
         npu_inst_pe_1_5_6_n101, npu_inst_pe_1_5_6_n100, npu_inst_pe_1_5_6_n99,
         npu_inst_pe_1_5_6_n98, npu_inst_pe_1_5_6_n36, npu_inst_pe_1_5_6_n35,
         npu_inst_pe_1_5_6_n34, npu_inst_pe_1_5_6_n33, npu_inst_pe_1_5_6_n32,
         npu_inst_pe_1_5_6_n31, npu_inst_pe_1_5_6_n30, npu_inst_pe_1_5_6_n29,
         npu_inst_pe_1_5_6_n28, npu_inst_pe_1_5_6_n25, npu_inst_pe_1_5_6_n24,
         npu_inst_pe_1_5_6_n23, npu_inst_pe_1_5_6_n22, npu_inst_pe_1_5_6_n21,
         npu_inst_pe_1_5_6_n20, npu_inst_pe_1_5_6_n19, npu_inst_pe_1_5_6_n18,
         npu_inst_pe_1_5_6_n17, npu_inst_pe_1_5_6_n16, npu_inst_pe_1_5_6_n15,
         npu_inst_pe_1_5_6_n14, npu_inst_pe_1_5_6_n13, npu_inst_pe_1_5_6_n12,
         npu_inst_pe_1_5_6_n11, npu_inst_pe_1_5_6_n10, npu_inst_pe_1_5_6_n9,
         npu_inst_pe_1_5_6_n8, npu_inst_pe_1_5_6_n7, npu_inst_pe_1_5_6_n6,
         npu_inst_pe_1_5_6_n5, npu_inst_pe_1_5_6_n4, npu_inst_pe_1_5_6_n3,
         npu_inst_pe_1_5_6_n2, npu_inst_pe_1_5_6_n1,
         npu_inst_pe_1_5_6_sub_77_carry_7_, npu_inst_pe_1_5_6_sub_77_carry_6_,
         npu_inst_pe_1_5_6_sub_77_carry_5_, npu_inst_pe_1_5_6_sub_77_carry_4_,
         npu_inst_pe_1_5_6_sub_77_carry_3_, npu_inst_pe_1_5_6_sub_77_carry_2_,
         npu_inst_pe_1_5_6_sub_77_carry_1_, npu_inst_pe_1_5_6_add_79_carry_7_,
         npu_inst_pe_1_5_6_add_79_carry_6_, npu_inst_pe_1_5_6_add_79_carry_5_,
         npu_inst_pe_1_5_6_add_79_carry_4_, npu_inst_pe_1_5_6_add_79_carry_3_,
         npu_inst_pe_1_5_6_add_79_carry_2_, npu_inst_pe_1_5_6_add_79_carry_1_,
         npu_inst_pe_1_5_6_n97, npu_inst_pe_1_5_6_n96, npu_inst_pe_1_5_6_n95,
         npu_inst_pe_1_5_6_n94, npu_inst_pe_1_5_6_n93, npu_inst_pe_1_5_6_n92,
         npu_inst_pe_1_5_6_n91, npu_inst_pe_1_5_6_n90, npu_inst_pe_1_5_6_n89,
         npu_inst_pe_1_5_6_n88, npu_inst_pe_1_5_6_n87, npu_inst_pe_1_5_6_n86,
         npu_inst_pe_1_5_6_n85, npu_inst_pe_1_5_6_n84, npu_inst_pe_1_5_6_n83,
         npu_inst_pe_1_5_6_n82, npu_inst_pe_1_5_6_n81, npu_inst_pe_1_5_6_n80,
         npu_inst_pe_1_5_6_n79, npu_inst_pe_1_5_6_n78, npu_inst_pe_1_5_6_n77,
         npu_inst_pe_1_5_6_n76, npu_inst_pe_1_5_6_n75, npu_inst_pe_1_5_6_n74,
         npu_inst_pe_1_5_6_n73, npu_inst_pe_1_5_6_n72, npu_inst_pe_1_5_6_n71,
         npu_inst_pe_1_5_6_n70, npu_inst_pe_1_5_6_n69, npu_inst_pe_1_5_6_n68,
         npu_inst_pe_1_5_6_n67, npu_inst_pe_1_5_6_n66, npu_inst_pe_1_5_6_n65,
         npu_inst_pe_1_5_6_n64, npu_inst_pe_1_5_6_n63, npu_inst_pe_1_5_6_n62,
         npu_inst_pe_1_5_6_n61, npu_inst_pe_1_5_6_n60, npu_inst_pe_1_5_6_n59,
         npu_inst_pe_1_5_6_n58, npu_inst_pe_1_5_6_n57, npu_inst_pe_1_5_6_n56,
         npu_inst_pe_1_5_6_n55, npu_inst_pe_1_5_6_n54, npu_inst_pe_1_5_6_n53,
         npu_inst_pe_1_5_6_n52, npu_inst_pe_1_5_6_n51, npu_inst_pe_1_5_6_n50,
         npu_inst_pe_1_5_6_n49, npu_inst_pe_1_5_6_n48, npu_inst_pe_1_5_6_n47,
         npu_inst_pe_1_5_6_n46, npu_inst_pe_1_5_6_n45, npu_inst_pe_1_5_6_n44,
         npu_inst_pe_1_5_6_n43, npu_inst_pe_1_5_6_n42, npu_inst_pe_1_5_6_n41,
         npu_inst_pe_1_5_6_n40, npu_inst_pe_1_5_6_n39, npu_inst_pe_1_5_6_n38,
         npu_inst_pe_1_5_6_n37, npu_inst_pe_1_5_6_n27, npu_inst_pe_1_5_6_n26,
         npu_inst_pe_1_5_6_net3426, npu_inst_pe_1_5_6_net3420,
         npu_inst_pe_1_5_6_N94, npu_inst_pe_1_5_6_N93, npu_inst_pe_1_5_6_N84,
         npu_inst_pe_1_5_6_N80, npu_inst_pe_1_5_6_N79, npu_inst_pe_1_5_6_N78,
         npu_inst_pe_1_5_6_N77, npu_inst_pe_1_5_6_N76, npu_inst_pe_1_5_6_N75,
         npu_inst_pe_1_5_6_N74, npu_inst_pe_1_5_6_N73, npu_inst_pe_1_5_6_N72,
         npu_inst_pe_1_5_6_N71, npu_inst_pe_1_5_6_N70, npu_inst_pe_1_5_6_N69,
         npu_inst_pe_1_5_6_N68, npu_inst_pe_1_5_6_N67, npu_inst_pe_1_5_6_N66,
         npu_inst_pe_1_5_6_N65, npu_inst_pe_1_5_6_int_data_0_,
         npu_inst_pe_1_5_6_int_data_1_, npu_inst_pe_1_5_6_int_q_weight_0_,
         npu_inst_pe_1_5_6_int_q_weight_1_,
         npu_inst_pe_1_5_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_6_int_q_reg_h_0__1_, npu_inst_pe_1_5_7_n118,
         npu_inst_pe_1_5_7_n117, npu_inst_pe_1_5_7_n116,
         npu_inst_pe_1_5_7_n115, npu_inst_pe_1_5_7_n114,
         npu_inst_pe_1_5_7_n113, npu_inst_pe_1_5_7_n112,
         npu_inst_pe_1_5_7_n111, npu_inst_pe_1_5_7_n110,
         npu_inst_pe_1_5_7_n109, npu_inst_pe_1_5_7_n108,
         npu_inst_pe_1_5_7_n107, npu_inst_pe_1_5_7_n106,
         npu_inst_pe_1_5_7_n105, npu_inst_pe_1_5_7_n104,
         npu_inst_pe_1_5_7_n103, npu_inst_pe_1_5_7_n102,
         npu_inst_pe_1_5_7_n101, npu_inst_pe_1_5_7_n100, npu_inst_pe_1_5_7_n99,
         npu_inst_pe_1_5_7_n98, npu_inst_pe_1_5_7_n36, npu_inst_pe_1_5_7_n35,
         npu_inst_pe_1_5_7_n34, npu_inst_pe_1_5_7_n33, npu_inst_pe_1_5_7_n32,
         npu_inst_pe_1_5_7_n31, npu_inst_pe_1_5_7_n30, npu_inst_pe_1_5_7_n29,
         npu_inst_pe_1_5_7_n28, npu_inst_pe_1_5_7_n25, npu_inst_pe_1_5_7_n24,
         npu_inst_pe_1_5_7_n23, npu_inst_pe_1_5_7_n22, npu_inst_pe_1_5_7_n21,
         npu_inst_pe_1_5_7_n20, npu_inst_pe_1_5_7_n19, npu_inst_pe_1_5_7_n18,
         npu_inst_pe_1_5_7_n17, npu_inst_pe_1_5_7_n16, npu_inst_pe_1_5_7_n15,
         npu_inst_pe_1_5_7_n14, npu_inst_pe_1_5_7_n13, npu_inst_pe_1_5_7_n12,
         npu_inst_pe_1_5_7_n11, npu_inst_pe_1_5_7_n10, npu_inst_pe_1_5_7_n9,
         npu_inst_pe_1_5_7_n8, npu_inst_pe_1_5_7_n7, npu_inst_pe_1_5_7_n6,
         npu_inst_pe_1_5_7_n5, npu_inst_pe_1_5_7_n4, npu_inst_pe_1_5_7_n3,
         npu_inst_pe_1_5_7_n2, npu_inst_pe_1_5_7_n1,
         npu_inst_pe_1_5_7_sub_77_carry_7_, npu_inst_pe_1_5_7_sub_77_carry_6_,
         npu_inst_pe_1_5_7_sub_77_carry_5_, npu_inst_pe_1_5_7_sub_77_carry_4_,
         npu_inst_pe_1_5_7_sub_77_carry_3_, npu_inst_pe_1_5_7_sub_77_carry_2_,
         npu_inst_pe_1_5_7_sub_77_carry_1_, npu_inst_pe_1_5_7_add_79_carry_7_,
         npu_inst_pe_1_5_7_add_79_carry_6_, npu_inst_pe_1_5_7_add_79_carry_5_,
         npu_inst_pe_1_5_7_add_79_carry_4_, npu_inst_pe_1_5_7_add_79_carry_3_,
         npu_inst_pe_1_5_7_add_79_carry_2_, npu_inst_pe_1_5_7_add_79_carry_1_,
         npu_inst_pe_1_5_7_n97, npu_inst_pe_1_5_7_n96, npu_inst_pe_1_5_7_n95,
         npu_inst_pe_1_5_7_n94, npu_inst_pe_1_5_7_n93, npu_inst_pe_1_5_7_n92,
         npu_inst_pe_1_5_7_n91, npu_inst_pe_1_5_7_n90, npu_inst_pe_1_5_7_n89,
         npu_inst_pe_1_5_7_n88, npu_inst_pe_1_5_7_n87, npu_inst_pe_1_5_7_n86,
         npu_inst_pe_1_5_7_n85, npu_inst_pe_1_5_7_n84, npu_inst_pe_1_5_7_n83,
         npu_inst_pe_1_5_7_n82, npu_inst_pe_1_5_7_n81, npu_inst_pe_1_5_7_n80,
         npu_inst_pe_1_5_7_n79, npu_inst_pe_1_5_7_n78, npu_inst_pe_1_5_7_n77,
         npu_inst_pe_1_5_7_n76, npu_inst_pe_1_5_7_n75, npu_inst_pe_1_5_7_n74,
         npu_inst_pe_1_5_7_n73, npu_inst_pe_1_5_7_n72, npu_inst_pe_1_5_7_n71,
         npu_inst_pe_1_5_7_n70, npu_inst_pe_1_5_7_n69, npu_inst_pe_1_5_7_n68,
         npu_inst_pe_1_5_7_n67, npu_inst_pe_1_5_7_n66, npu_inst_pe_1_5_7_n65,
         npu_inst_pe_1_5_7_n64, npu_inst_pe_1_5_7_n63, npu_inst_pe_1_5_7_n62,
         npu_inst_pe_1_5_7_n61, npu_inst_pe_1_5_7_n60, npu_inst_pe_1_5_7_n59,
         npu_inst_pe_1_5_7_n58, npu_inst_pe_1_5_7_n57, npu_inst_pe_1_5_7_n56,
         npu_inst_pe_1_5_7_n55, npu_inst_pe_1_5_7_n54, npu_inst_pe_1_5_7_n53,
         npu_inst_pe_1_5_7_n52, npu_inst_pe_1_5_7_n51, npu_inst_pe_1_5_7_n50,
         npu_inst_pe_1_5_7_n49, npu_inst_pe_1_5_7_n48, npu_inst_pe_1_5_7_n47,
         npu_inst_pe_1_5_7_n46, npu_inst_pe_1_5_7_n45, npu_inst_pe_1_5_7_n44,
         npu_inst_pe_1_5_7_n43, npu_inst_pe_1_5_7_n42, npu_inst_pe_1_5_7_n41,
         npu_inst_pe_1_5_7_n40, npu_inst_pe_1_5_7_n39, npu_inst_pe_1_5_7_n38,
         npu_inst_pe_1_5_7_n37, npu_inst_pe_1_5_7_n27, npu_inst_pe_1_5_7_n26,
         npu_inst_pe_1_5_7_net3403, npu_inst_pe_1_5_7_net3397,
         npu_inst_pe_1_5_7_N94, npu_inst_pe_1_5_7_N93, npu_inst_pe_1_5_7_N84,
         npu_inst_pe_1_5_7_N80, npu_inst_pe_1_5_7_N79, npu_inst_pe_1_5_7_N78,
         npu_inst_pe_1_5_7_N77, npu_inst_pe_1_5_7_N76, npu_inst_pe_1_5_7_N75,
         npu_inst_pe_1_5_7_N74, npu_inst_pe_1_5_7_N73, npu_inst_pe_1_5_7_N72,
         npu_inst_pe_1_5_7_N71, npu_inst_pe_1_5_7_N70, npu_inst_pe_1_5_7_N69,
         npu_inst_pe_1_5_7_N68, npu_inst_pe_1_5_7_N67, npu_inst_pe_1_5_7_N66,
         npu_inst_pe_1_5_7_N65, npu_inst_pe_1_5_7_int_data_0_,
         npu_inst_pe_1_5_7_int_data_1_, npu_inst_pe_1_5_7_int_q_weight_0_,
         npu_inst_pe_1_5_7_int_q_weight_1_,
         npu_inst_pe_1_5_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_5_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_5_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_5_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_5_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_5_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_5_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_5_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_5_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_5_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_5_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_5_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_5_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_5_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_5_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_5_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_5_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_5_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_5_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_5_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_5_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_5_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_5_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_5_7_int_q_reg_h_0__1_, npu_inst_pe_1_6_0_n118,
         npu_inst_pe_1_6_0_n117, npu_inst_pe_1_6_0_n116,
         npu_inst_pe_1_6_0_n115, npu_inst_pe_1_6_0_n114,
         npu_inst_pe_1_6_0_n113, npu_inst_pe_1_6_0_n112,
         npu_inst_pe_1_6_0_n111, npu_inst_pe_1_6_0_n110,
         npu_inst_pe_1_6_0_n109, npu_inst_pe_1_6_0_n108,
         npu_inst_pe_1_6_0_n107, npu_inst_pe_1_6_0_n106,
         npu_inst_pe_1_6_0_n105, npu_inst_pe_1_6_0_n104,
         npu_inst_pe_1_6_0_n103, npu_inst_pe_1_6_0_n102,
         npu_inst_pe_1_6_0_n101, npu_inst_pe_1_6_0_n100, npu_inst_pe_1_6_0_n99,
         npu_inst_pe_1_6_0_n98, npu_inst_pe_1_6_0_n36, npu_inst_pe_1_6_0_n35,
         npu_inst_pe_1_6_0_n34, npu_inst_pe_1_6_0_n33, npu_inst_pe_1_6_0_n32,
         npu_inst_pe_1_6_0_n31, npu_inst_pe_1_6_0_n30, npu_inst_pe_1_6_0_n29,
         npu_inst_pe_1_6_0_n28, npu_inst_pe_1_6_0_n25, npu_inst_pe_1_6_0_n24,
         npu_inst_pe_1_6_0_n23, npu_inst_pe_1_6_0_n22, npu_inst_pe_1_6_0_n21,
         npu_inst_pe_1_6_0_n20, npu_inst_pe_1_6_0_n19, npu_inst_pe_1_6_0_n18,
         npu_inst_pe_1_6_0_n17, npu_inst_pe_1_6_0_n16, npu_inst_pe_1_6_0_n15,
         npu_inst_pe_1_6_0_n14, npu_inst_pe_1_6_0_n13, npu_inst_pe_1_6_0_n12,
         npu_inst_pe_1_6_0_n11, npu_inst_pe_1_6_0_n10, npu_inst_pe_1_6_0_n9,
         npu_inst_pe_1_6_0_n8, npu_inst_pe_1_6_0_n7, npu_inst_pe_1_6_0_n6,
         npu_inst_pe_1_6_0_n5, npu_inst_pe_1_6_0_n4, npu_inst_pe_1_6_0_n3,
         npu_inst_pe_1_6_0_n2, npu_inst_pe_1_6_0_n1,
         npu_inst_pe_1_6_0_sub_77_carry_7_, npu_inst_pe_1_6_0_sub_77_carry_6_,
         npu_inst_pe_1_6_0_sub_77_carry_5_, npu_inst_pe_1_6_0_sub_77_carry_4_,
         npu_inst_pe_1_6_0_sub_77_carry_3_, npu_inst_pe_1_6_0_sub_77_carry_2_,
         npu_inst_pe_1_6_0_sub_77_carry_1_, npu_inst_pe_1_6_0_add_79_carry_7_,
         npu_inst_pe_1_6_0_add_79_carry_6_, npu_inst_pe_1_6_0_add_79_carry_5_,
         npu_inst_pe_1_6_0_add_79_carry_4_, npu_inst_pe_1_6_0_add_79_carry_3_,
         npu_inst_pe_1_6_0_add_79_carry_2_, npu_inst_pe_1_6_0_add_79_carry_1_,
         npu_inst_pe_1_6_0_n97, npu_inst_pe_1_6_0_n96, npu_inst_pe_1_6_0_n95,
         npu_inst_pe_1_6_0_n94, npu_inst_pe_1_6_0_n93, npu_inst_pe_1_6_0_n92,
         npu_inst_pe_1_6_0_n91, npu_inst_pe_1_6_0_n90, npu_inst_pe_1_6_0_n89,
         npu_inst_pe_1_6_0_n88, npu_inst_pe_1_6_0_n87, npu_inst_pe_1_6_0_n86,
         npu_inst_pe_1_6_0_n85, npu_inst_pe_1_6_0_n84, npu_inst_pe_1_6_0_n83,
         npu_inst_pe_1_6_0_n82, npu_inst_pe_1_6_0_n81, npu_inst_pe_1_6_0_n80,
         npu_inst_pe_1_6_0_n79, npu_inst_pe_1_6_0_n78, npu_inst_pe_1_6_0_n77,
         npu_inst_pe_1_6_0_n76, npu_inst_pe_1_6_0_n75, npu_inst_pe_1_6_0_n74,
         npu_inst_pe_1_6_0_n73, npu_inst_pe_1_6_0_n72, npu_inst_pe_1_6_0_n71,
         npu_inst_pe_1_6_0_n70, npu_inst_pe_1_6_0_n69, npu_inst_pe_1_6_0_n68,
         npu_inst_pe_1_6_0_n67, npu_inst_pe_1_6_0_n66, npu_inst_pe_1_6_0_n65,
         npu_inst_pe_1_6_0_n64, npu_inst_pe_1_6_0_n63, npu_inst_pe_1_6_0_n62,
         npu_inst_pe_1_6_0_n61, npu_inst_pe_1_6_0_n60, npu_inst_pe_1_6_0_n59,
         npu_inst_pe_1_6_0_n58, npu_inst_pe_1_6_0_n57, npu_inst_pe_1_6_0_n56,
         npu_inst_pe_1_6_0_n55, npu_inst_pe_1_6_0_n54, npu_inst_pe_1_6_0_n53,
         npu_inst_pe_1_6_0_n52, npu_inst_pe_1_6_0_n51, npu_inst_pe_1_6_0_n50,
         npu_inst_pe_1_6_0_n49, npu_inst_pe_1_6_0_n48, npu_inst_pe_1_6_0_n47,
         npu_inst_pe_1_6_0_n46, npu_inst_pe_1_6_0_n45, npu_inst_pe_1_6_0_n44,
         npu_inst_pe_1_6_0_n43, npu_inst_pe_1_6_0_n42, npu_inst_pe_1_6_0_n41,
         npu_inst_pe_1_6_0_n40, npu_inst_pe_1_6_0_n39, npu_inst_pe_1_6_0_n38,
         npu_inst_pe_1_6_0_n37, npu_inst_pe_1_6_0_n27, npu_inst_pe_1_6_0_n26,
         npu_inst_pe_1_6_0_net3380, npu_inst_pe_1_6_0_net3374,
         npu_inst_pe_1_6_0_N94, npu_inst_pe_1_6_0_N93, npu_inst_pe_1_6_0_N84,
         npu_inst_pe_1_6_0_N80, npu_inst_pe_1_6_0_N79, npu_inst_pe_1_6_0_N78,
         npu_inst_pe_1_6_0_N77, npu_inst_pe_1_6_0_N76, npu_inst_pe_1_6_0_N75,
         npu_inst_pe_1_6_0_N74, npu_inst_pe_1_6_0_N73, npu_inst_pe_1_6_0_N72,
         npu_inst_pe_1_6_0_N71, npu_inst_pe_1_6_0_N70, npu_inst_pe_1_6_0_N69,
         npu_inst_pe_1_6_0_N68, npu_inst_pe_1_6_0_N67, npu_inst_pe_1_6_0_N66,
         npu_inst_pe_1_6_0_N65, npu_inst_pe_1_6_0_int_data_0_,
         npu_inst_pe_1_6_0_int_data_1_, npu_inst_pe_1_6_0_int_q_weight_0_,
         npu_inst_pe_1_6_0_int_q_weight_1_,
         npu_inst_pe_1_6_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_0_int_q_reg_h_0__1_, npu_inst_pe_1_6_0_o_data_h_0_,
         npu_inst_pe_1_6_0_o_data_h_1_, npu_inst_pe_1_6_1_n118,
         npu_inst_pe_1_6_1_n117, npu_inst_pe_1_6_1_n116,
         npu_inst_pe_1_6_1_n115, npu_inst_pe_1_6_1_n114,
         npu_inst_pe_1_6_1_n113, npu_inst_pe_1_6_1_n112,
         npu_inst_pe_1_6_1_n111, npu_inst_pe_1_6_1_n110,
         npu_inst_pe_1_6_1_n109, npu_inst_pe_1_6_1_n108,
         npu_inst_pe_1_6_1_n107, npu_inst_pe_1_6_1_n106,
         npu_inst_pe_1_6_1_n105, npu_inst_pe_1_6_1_n104,
         npu_inst_pe_1_6_1_n103, npu_inst_pe_1_6_1_n102,
         npu_inst_pe_1_6_1_n101, npu_inst_pe_1_6_1_n100, npu_inst_pe_1_6_1_n99,
         npu_inst_pe_1_6_1_n98, npu_inst_pe_1_6_1_n36, npu_inst_pe_1_6_1_n35,
         npu_inst_pe_1_6_1_n34, npu_inst_pe_1_6_1_n33, npu_inst_pe_1_6_1_n32,
         npu_inst_pe_1_6_1_n31, npu_inst_pe_1_6_1_n30, npu_inst_pe_1_6_1_n29,
         npu_inst_pe_1_6_1_n28, npu_inst_pe_1_6_1_n25, npu_inst_pe_1_6_1_n24,
         npu_inst_pe_1_6_1_n23, npu_inst_pe_1_6_1_n22, npu_inst_pe_1_6_1_n21,
         npu_inst_pe_1_6_1_n20, npu_inst_pe_1_6_1_n19, npu_inst_pe_1_6_1_n18,
         npu_inst_pe_1_6_1_n17, npu_inst_pe_1_6_1_n16, npu_inst_pe_1_6_1_n15,
         npu_inst_pe_1_6_1_n14, npu_inst_pe_1_6_1_n13, npu_inst_pe_1_6_1_n12,
         npu_inst_pe_1_6_1_n11, npu_inst_pe_1_6_1_n10, npu_inst_pe_1_6_1_n9,
         npu_inst_pe_1_6_1_n8, npu_inst_pe_1_6_1_n7, npu_inst_pe_1_6_1_n6,
         npu_inst_pe_1_6_1_n5, npu_inst_pe_1_6_1_n4, npu_inst_pe_1_6_1_n3,
         npu_inst_pe_1_6_1_n2, npu_inst_pe_1_6_1_n1,
         npu_inst_pe_1_6_1_sub_77_carry_7_, npu_inst_pe_1_6_1_sub_77_carry_6_,
         npu_inst_pe_1_6_1_sub_77_carry_5_, npu_inst_pe_1_6_1_sub_77_carry_4_,
         npu_inst_pe_1_6_1_sub_77_carry_3_, npu_inst_pe_1_6_1_sub_77_carry_2_,
         npu_inst_pe_1_6_1_sub_77_carry_1_, npu_inst_pe_1_6_1_add_79_carry_7_,
         npu_inst_pe_1_6_1_add_79_carry_6_, npu_inst_pe_1_6_1_add_79_carry_5_,
         npu_inst_pe_1_6_1_add_79_carry_4_, npu_inst_pe_1_6_1_add_79_carry_3_,
         npu_inst_pe_1_6_1_add_79_carry_2_, npu_inst_pe_1_6_1_add_79_carry_1_,
         npu_inst_pe_1_6_1_n97, npu_inst_pe_1_6_1_n96, npu_inst_pe_1_6_1_n95,
         npu_inst_pe_1_6_1_n94, npu_inst_pe_1_6_1_n93, npu_inst_pe_1_6_1_n92,
         npu_inst_pe_1_6_1_n91, npu_inst_pe_1_6_1_n90, npu_inst_pe_1_6_1_n89,
         npu_inst_pe_1_6_1_n88, npu_inst_pe_1_6_1_n87, npu_inst_pe_1_6_1_n86,
         npu_inst_pe_1_6_1_n85, npu_inst_pe_1_6_1_n84, npu_inst_pe_1_6_1_n83,
         npu_inst_pe_1_6_1_n82, npu_inst_pe_1_6_1_n81, npu_inst_pe_1_6_1_n80,
         npu_inst_pe_1_6_1_n79, npu_inst_pe_1_6_1_n78, npu_inst_pe_1_6_1_n77,
         npu_inst_pe_1_6_1_n76, npu_inst_pe_1_6_1_n75, npu_inst_pe_1_6_1_n74,
         npu_inst_pe_1_6_1_n73, npu_inst_pe_1_6_1_n72, npu_inst_pe_1_6_1_n71,
         npu_inst_pe_1_6_1_n70, npu_inst_pe_1_6_1_n69, npu_inst_pe_1_6_1_n68,
         npu_inst_pe_1_6_1_n67, npu_inst_pe_1_6_1_n66, npu_inst_pe_1_6_1_n65,
         npu_inst_pe_1_6_1_n64, npu_inst_pe_1_6_1_n63, npu_inst_pe_1_6_1_n62,
         npu_inst_pe_1_6_1_n61, npu_inst_pe_1_6_1_n60, npu_inst_pe_1_6_1_n59,
         npu_inst_pe_1_6_1_n58, npu_inst_pe_1_6_1_n57, npu_inst_pe_1_6_1_n56,
         npu_inst_pe_1_6_1_n55, npu_inst_pe_1_6_1_n54, npu_inst_pe_1_6_1_n53,
         npu_inst_pe_1_6_1_n52, npu_inst_pe_1_6_1_n51, npu_inst_pe_1_6_1_n50,
         npu_inst_pe_1_6_1_n49, npu_inst_pe_1_6_1_n48, npu_inst_pe_1_6_1_n47,
         npu_inst_pe_1_6_1_n46, npu_inst_pe_1_6_1_n45, npu_inst_pe_1_6_1_n44,
         npu_inst_pe_1_6_1_n43, npu_inst_pe_1_6_1_n42, npu_inst_pe_1_6_1_n41,
         npu_inst_pe_1_6_1_n40, npu_inst_pe_1_6_1_n39, npu_inst_pe_1_6_1_n38,
         npu_inst_pe_1_6_1_n37, npu_inst_pe_1_6_1_n27, npu_inst_pe_1_6_1_n26,
         npu_inst_pe_1_6_1_net3357, npu_inst_pe_1_6_1_net3351,
         npu_inst_pe_1_6_1_N94, npu_inst_pe_1_6_1_N93, npu_inst_pe_1_6_1_N84,
         npu_inst_pe_1_6_1_N80, npu_inst_pe_1_6_1_N79, npu_inst_pe_1_6_1_N78,
         npu_inst_pe_1_6_1_N77, npu_inst_pe_1_6_1_N76, npu_inst_pe_1_6_1_N75,
         npu_inst_pe_1_6_1_N74, npu_inst_pe_1_6_1_N73, npu_inst_pe_1_6_1_N72,
         npu_inst_pe_1_6_1_N71, npu_inst_pe_1_6_1_N70, npu_inst_pe_1_6_1_N69,
         npu_inst_pe_1_6_1_N68, npu_inst_pe_1_6_1_N67, npu_inst_pe_1_6_1_N66,
         npu_inst_pe_1_6_1_N65, npu_inst_pe_1_6_1_int_data_0_,
         npu_inst_pe_1_6_1_int_data_1_, npu_inst_pe_1_6_1_int_q_weight_0_,
         npu_inst_pe_1_6_1_int_q_weight_1_,
         npu_inst_pe_1_6_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_1_int_q_reg_h_0__1_, npu_inst_pe_1_6_2_n118,
         npu_inst_pe_1_6_2_n117, npu_inst_pe_1_6_2_n116,
         npu_inst_pe_1_6_2_n115, npu_inst_pe_1_6_2_n114,
         npu_inst_pe_1_6_2_n113, npu_inst_pe_1_6_2_n112,
         npu_inst_pe_1_6_2_n111, npu_inst_pe_1_6_2_n110,
         npu_inst_pe_1_6_2_n109, npu_inst_pe_1_6_2_n108,
         npu_inst_pe_1_6_2_n107, npu_inst_pe_1_6_2_n106,
         npu_inst_pe_1_6_2_n105, npu_inst_pe_1_6_2_n104,
         npu_inst_pe_1_6_2_n103, npu_inst_pe_1_6_2_n102,
         npu_inst_pe_1_6_2_n101, npu_inst_pe_1_6_2_n100, npu_inst_pe_1_6_2_n99,
         npu_inst_pe_1_6_2_n98, npu_inst_pe_1_6_2_n36, npu_inst_pe_1_6_2_n35,
         npu_inst_pe_1_6_2_n34, npu_inst_pe_1_6_2_n33, npu_inst_pe_1_6_2_n32,
         npu_inst_pe_1_6_2_n31, npu_inst_pe_1_6_2_n30, npu_inst_pe_1_6_2_n29,
         npu_inst_pe_1_6_2_n28, npu_inst_pe_1_6_2_n25, npu_inst_pe_1_6_2_n24,
         npu_inst_pe_1_6_2_n23, npu_inst_pe_1_6_2_n22, npu_inst_pe_1_6_2_n21,
         npu_inst_pe_1_6_2_n20, npu_inst_pe_1_6_2_n19, npu_inst_pe_1_6_2_n18,
         npu_inst_pe_1_6_2_n17, npu_inst_pe_1_6_2_n16, npu_inst_pe_1_6_2_n15,
         npu_inst_pe_1_6_2_n14, npu_inst_pe_1_6_2_n13, npu_inst_pe_1_6_2_n12,
         npu_inst_pe_1_6_2_n11, npu_inst_pe_1_6_2_n10, npu_inst_pe_1_6_2_n9,
         npu_inst_pe_1_6_2_n8, npu_inst_pe_1_6_2_n7, npu_inst_pe_1_6_2_n6,
         npu_inst_pe_1_6_2_n5, npu_inst_pe_1_6_2_n4, npu_inst_pe_1_6_2_n3,
         npu_inst_pe_1_6_2_n2, npu_inst_pe_1_6_2_n1,
         npu_inst_pe_1_6_2_sub_77_carry_7_, npu_inst_pe_1_6_2_sub_77_carry_6_,
         npu_inst_pe_1_6_2_sub_77_carry_5_, npu_inst_pe_1_6_2_sub_77_carry_4_,
         npu_inst_pe_1_6_2_sub_77_carry_3_, npu_inst_pe_1_6_2_sub_77_carry_2_,
         npu_inst_pe_1_6_2_sub_77_carry_1_, npu_inst_pe_1_6_2_add_79_carry_7_,
         npu_inst_pe_1_6_2_add_79_carry_6_, npu_inst_pe_1_6_2_add_79_carry_5_,
         npu_inst_pe_1_6_2_add_79_carry_4_, npu_inst_pe_1_6_2_add_79_carry_3_,
         npu_inst_pe_1_6_2_add_79_carry_2_, npu_inst_pe_1_6_2_add_79_carry_1_,
         npu_inst_pe_1_6_2_n97, npu_inst_pe_1_6_2_n96, npu_inst_pe_1_6_2_n95,
         npu_inst_pe_1_6_2_n94, npu_inst_pe_1_6_2_n93, npu_inst_pe_1_6_2_n92,
         npu_inst_pe_1_6_2_n91, npu_inst_pe_1_6_2_n90, npu_inst_pe_1_6_2_n89,
         npu_inst_pe_1_6_2_n88, npu_inst_pe_1_6_2_n87, npu_inst_pe_1_6_2_n86,
         npu_inst_pe_1_6_2_n85, npu_inst_pe_1_6_2_n84, npu_inst_pe_1_6_2_n83,
         npu_inst_pe_1_6_2_n82, npu_inst_pe_1_6_2_n81, npu_inst_pe_1_6_2_n80,
         npu_inst_pe_1_6_2_n79, npu_inst_pe_1_6_2_n78, npu_inst_pe_1_6_2_n77,
         npu_inst_pe_1_6_2_n76, npu_inst_pe_1_6_2_n75, npu_inst_pe_1_6_2_n74,
         npu_inst_pe_1_6_2_n73, npu_inst_pe_1_6_2_n72, npu_inst_pe_1_6_2_n71,
         npu_inst_pe_1_6_2_n70, npu_inst_pe_1_6_2_n69, npu_inst_pe_1_6_2_n68,
         npu_inst_pe_1_6_2_n67, npu_inst_pe_1_6_2_n66, npu_inst_pe_1_6_2_n65,
         npu_inst_pe_1_6_2_n64, npu_inst_pe_1_6_2_n63, npu_inst_pe_1_6_2_n62,
         npu_inst_pe_1_6_2_n61, npu_inst_pe_1_6_2_n60, npu_inst_pe_1_6_2_n59,
         npu_inst_pe_1_6_2_n58, npu_inst_pe_1_6_2_n57, npu_inst_pe_1_6_2_n56,
         npu_inst_pe_1_6_2_n55, npu_inst_pe_1_6_2_n54, npu_inst_pe_1_6_2_n53,
         npu_inst_pe_1_6_2_n52, npu_inst_pe_1_6_2_n51, npu_inst_pe_1_6_2_n50,
         npu_inst_pe_1_6_2_n49, npu_inst_pe_1_6_2_n48, npu_inst_pe_1_6_2_n47,
         npu_inst_pe_1_6_2_n46, npu_inst_pe_1_6_2_n45, npu_inst_pe_1_6_2_n44,
         npu_inst_pe_1_6_2_n43, npu_inst_pe_1_6_2_n42, npu_inst_pe_1_6_2_n41,
         npu_inst_pe_1_6_2_n40, npu_inst_pe_1_6_2_n39, npu_inst_pe_1_6_2_n38,
         npu_inst_pe_1_6_2_n37, npu_inst_pe_1_6_2_n27, npu_inst_pe_1_6_2_n26,
         npu_inst_pe_1_6_2_net3334, npu_inst_pe_1_6_2_net3328,
         npu_inst_pe_1_6_2_N94, npu_inst_pe_1_6_2_N93, npu_inst_pe_1_6_2_N84,
         npu_inst_pe_1_6_2_N80, npu_inst_pe_1_6_2_N79, npu_inst_pe_1_6_2_N78,
         npu_inst_pe_1_6_2_N77, npu_inst_pe_1_6_2_N76, npu_inst_pe_1_6_2_N75,
         npu_inst_pe_1_6_2_N74, npu_inst_pe_1_6_2_N73, npu_inst_pe_1_6_2_N72,
         npu_inst_pe_1_6_2_N71, npu_inst_pe_1_6_2_N70, npu_inst_pe_1_6_2_N69,
         npu_inst_pe_1_6_2_N68, npu_inst_pe_1_6_2_N67, npu_inst_pe_1_6_2_N66,
         npu_inst_pe_1_6_2_N65, npu_inst_pe_1_6_2_int_data_0_,
         npu_inst_pe_1_6_2_int_data_1_, npu_inst_pe_1_6_2_int_q_weight_0_,
         npu_inst_pe_1_6_2_int_q_weight_1_,
         npu_inst_pe_1_6_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_2_int_q_reg_h_0__1_, npu_inst_pe_1_6_3_n118,
         npu_inst_pe_1_6_3_n117, npu_inst_pe_1_6_3_n116,
         npu_inst_pe_1_6_3_n115, npu_inst_pe_1_6_3_n114,
         npu_inst_pe_1_6_3_n113, npu_inst_pe_1_6_3_n112,
         npu_inst_pe_1_6_3_n111, npu_inst_pe_1_6_3_n110,
         npu_inst_pe_1_6_3_n109, npu_inst_pe_1_6_3_n108,
         npu_inst_pe_1_6_3_n107, npu_inst_pe_1_6_3_n106,
         npu_inst_pe_1_6_3_n105, npu_inst_pe_1_6_3_n104,
         npu_inst_pe_1_6_3_n103, npu_inst_pe_1_6_3_n102,
         npu_inst_pe_1_6_3_n101, npu_inst_pe_1_6_3_n100, npu_inst_pe_1_6_3_n99,
         npu_inst_pe_1_6_3_n98, npu_inst_pe_1_6_3_n36, npu_inst_pe_1_6_3_n35,
         npu_inst_pe_1_6_3_n34, npu_inst_pe_1_6_3_n33, npu_inst_pe_1_6_3_n32,
         npu_inst_pe_1_6_3_n31, npu_inst_pe_1_6_3_n30, npu_inst_pe_1_6_3_n29,
         npu_inst_pe_1_6_3_n28, npu_inst_pe_1_6_3_n25, npu_inst_pe_1_6_3_n24,
         npu_inst_pe_1_6_3_n23, npu_inst_pe_1_6_3_n22, npu_inst_pe_1_6_3_n21,
         npu_inst_pe_1_6_3_n20, npu_inst_pe_1_6_3_n19, npu_inst_pe_1_6_3_n18,
         npu_inst_pe_1_6_3_n17, npu_inst_pe_1_6_3_n16, npu_inst_pe_1_6_3_n15,
         npu_inst_pe_1_6_3_n14, npu_inst_pe_1_6_3_n13, npu_inst_pe_1_6_3_n12,
         npu_inst_pe_1_6_3_n11, npu_inst_pe_1_6_3_n10, npu_inst_pe_1_6_3_n9,
         npu_inst_pe_1_6_3_n8, npu_inst_pe_1_6_3_n7, npu_inst_pe_1_6_3_n6,
         npu_inst_pe_1_6_3_n5, npu_inst_pe_1_6_3_n4, npu_inst_pe_1_6_3_n3,
         npu_inst_pe_1_6_3_n2, npu_inst_pe_1_6_3_n1,
         npu_inst_pe_1_6_3_sub_77_carry_7_, npu_inst_pe_1_6_3_sub_77_carry_6_,
         npu_inst_pe_1_6_3_sub_77_carry_5_, npu_inst_pe_1_6_3_sub_77_carry_4_,
         npu_inst_pe_1_6_3_sub_77_carry_3_, npu_inst_pe_1_6_3_sub_77_carry_2_,
         npu_inst_pe_1_6_3_sub_77_carry_1_, npu_inst_pe_1_6_3_add_79_carry_7_,
         npu_inst_pe_1_6_3_add_79_carry_6_, npu_inst_pe_1_6_3_add_79_carry_5_,
         npu_inst_pe_1_6_3_add_79_carry_4_, npu_inst_pe_1_6_3_add_79_carry_3_,
         npu_inst_pe_1_6_3_add_79_carry_2_, npu_inst_pe_1_6_3_add_79_carry_1_,
         npu_inst_pe_1_6_3_n97, npu_inst_pe_1_6_3_n96, npu_inst_pe_1_6_3_n95,
         npu_inst_pe_1_6_3_n94, npu_inst_pe_1_6_3_n93, npu_inst_pe_1_6_3_n92,
         npu_inst_pe_1_6_3_n91, npu_inst_pe_1_6_3_n90, npu_inst_pe_1_6_3_n89,
         npu_inst_pe_1_6_3_n88, npu_inst_pe_1_6_3_n87, npu_inst_pe_1_6_3_n86,
         npu_inst_pe_1_6_3_n85, npu_inst_pe_1_6_3_n84, npu_inst_pe_1_6_3_n83,
         npu_inst_pe_1_6_3_n82, npu_inst_pe_1_6_3_n81, npu_inst_pe_1_6_3_n80,
         npu_inst_pe_1_6_3_n79, npu_inst_pe_1_6_3_n78, npu_inst_pe_1_6_3_n77,
         npu_inst_pe_1_6_3_n76, npu_inst_pe_1_6_3_n75, npu_inst_pe_1_6_3_n74,
         npu_inst_pe_1_6_3_n73, npu_inst_pe_1_6_3_n72, npu_inst_pe_1_6_3_n71,
         npu_inst_pe_1_6_3_n70, npu_inst_pe_1_6_3_n69, npu_inst_pe_1_6_3_n68,
         npu_inst_pe_1_6_3_n67, npu_inst_pe_1_6_3_n66, npu_inst_pe_1_6_3_n65,
         npu_inst_pe_1_6_3_n64, npu_inst_pe_1_6_3_n63, npu_inst_pe_1_6_3_n62,
         npu_inst_pe_1_6_3_n61, npu_inst_pe_1_6_3_n60, npu_inst_pe_1_6_3_n59,
         npu_inst_pe_1_6_3_n58, npu_inst_pe_1_6_3_n57, npu_inst_pe_1_6_3_n56,
         npu_inst_pe_1_6_3_n55, npu_inst_pe_1_6_3_n54, npu_inst_pe_1_6_3_n53,
         npu_inst_pe_1_6_3_n52, npu_inst_pe_1_6_3_n51, npu_inst_pe_1_6_3_n50,
         npu_inst_pe_1_6_3_n49, npu_inst_pe_1_6_3_n48, npu_inst_pe_1_6_3_n47,
         npu_inst_pe_1_6_3_n46, npu_inst_pe_1_6_3_n45, npu_inst_pe_1_6_3_n44,
         npu_inst_pe_1_6_3_n43, npu_inst_pe_1_6_3_n42, npu_inst_pe_1_6_3_n41,
         npu_inst_pe_1_6_3_n40, npu_inst_pe_1_6_3_n39, npu_inst_pe_1_6_3_n38,
         npu_inst_pe_1_6_3_n37, npu_inst_pe_1_6_3_n27, npu_inst_pe_1_6_3_n26,
         npu_inst_pe_1_6_3_net3311, npu_inst_pe_1_6_3_net3305,
         npu_inst_pe_1_6_3_N94, npu_inst_pe_1_6_3_N93, npu_inst_pe_1_6_3_N84,
         npu_inst_pe_1_6_3_N80, npu_inst_pe_1_6_3_N79, npu_inst_pe_1_6_3_N78,
         npu_inst_pe_1_6_3_N77, npu_inst_pe_1_6_3_N76, npu_inst_pe_1_6_3_N75,
         npu_inst_pe_1_6_3_N74, npu_inst_pe_1_6_3_N73, npu_inst_pe_1_6_3_N72,
         npu_inst_pe_1_6_3_N71, npu_inst_pe_1_6_3_N70, npu_inst_pe_1_6_3_N69,
         npu_inst_pe_1_6_3_N68, npu_inst_pe_1_6_3_N67, npu_inst_pe_1_6_3_N66,
         npu_inst_pe_1_6_3_N65, npu_inst_pe_1_6_3_int_data_0_,
         npu_inst_pe_1_6_3_int_data_1_, npu_inst_pe_1_6_3_int_q_weight_0_,
         npu_inst_pe_1_6_3_int_q_weight_1_,
         npu_inst_pe_1_6_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_3_int_q_reg_h_0__1_, npu_inst_pe_1_6_4_n117,
         npu_inst_pe_1_6_4_n116, npu_inst_pe_1_6_4_n115,
         npu_inst_pe_1_6_4_n114, npu_inst_pe_1_6_4_n113,
         npu_inst_pe_1_6_4_n112, npu_inst_pe_1_6_4_n111,
         npu_inst_pe_1_6_4_n110, npu_inst_pe_1_6_4_n109,
         npu_inst_pe_1_6_4_n108, npu_inst_pe_1_6_4_n107,
         npu_inst_pe_1_6_4_n106, npu_inst_pe_1_6_4_n105,
         npu_inst_pe_1_6_4_n104, npu_inst_pe_1_6_4_n103,
         npu_inst_pe_1_6_4_n102, npu_inst_pe_1_6_4_n101,
         npu_inst_pe_1_6_4_n100, npu_inst_pe_1_6_4_n99, npu_inst_pe_1_6_4_n98,
         npu_inst_pe_1_6_4_n36, npu_inst_pe_1_6_4_n35, npu_inst_pe_1_6_4_n34,
         npu_inst_pe_1_6_4_n33, npu_inst_pe_1_6_4_n32, npu_inst_pe_1_6_4_n31,
         npu_inst_pe_1_6_4_n30, npu_inst_pe_1_6_4_n29, npu_inst_pe_1_6_4_n28,
         npu_inst_pe_1_6_4_n25, npu_inst_pe_1_6_4_n24, npu_inst_pe_1_6_4_n23,
         npu_inst_pe_1_6_4_n22, npu_inst_pe_1_6_4_n21, npu_inst_pe_1_6_4_n20,
         npu_inst_pe_1_6_4_n19, npu_inst_pe_1_6_4_n18, npu_inst_pe_1_6_4_n17,
         npu_inst_pe_1_6_4_n16, npu_inst_pe_1_6_4_n15, npu_inst_pe_1_6_4_n14,
         npu_inst_pe_1_6_4_n13, npu_inst_pe_1_6_4_n12, npu_inst_pe_1_6_4_n11,
         npu_inst_pe_1_6_4_n10, npu_inst_pe_1_6_4_n9, npu_inst_pe_1_6_4_n8,
         npu_inst_pe_1_6_4_n7, npu_inst_pe_1_6_4_n6, npu_inst_pe_1_6_4_n5,
         npu_inst_pe_1_6_4_n4, npu_inst_pe_1_6_4_n3, npu_inst_pe_1_6_4_n2,
         npu_inst_pe_1_6_4_n1, npu_inst_pe_1_6_4_sub_77_carry_7_,
         npu_inst_pe_1_6_4_sub_77_carry_6_, npu_inst_pe_1_6_4_sub_77_carry_5_,
         npu_inst_pe_1_6_4_sub_77_carry_4_, npu_inst_pe_1_6_4_sub_77_carry_3_,
         npu_inst_pe_1_6_4_sub_77_carry_2_, npu_inst_pe_1_6_4_sub_77_carry_1_,
         npu_inst_pe_1_6_4_add_79_carry_7_, npu_inst_pe_1_6_4_add_79_carry_6_,
         npu_inst_pe_1_6_4_add_79_carry_5_, npu_inst_pe_1_6_4_add_79_carry_4_,
         npu_inst_pe_1_6_4_add_79_carry_3_, npu_inst_pe_1_6_4_add_79_carry_2_,
         npu_inst_pe_1_6_4_add_79_carry_1_, npu_inst_pe_1_6_4_n97,
         npu_inst_pe_1_6_4_n96, npu_inst_pe_1_6_4_n95, npu_inst_pe_1_6_4_n94,
         npu_inst_pe_1_6_4_n93, npu_inst_pe_1_6_4_n92, npu_inst_pe_1_6_4_n91,
         npu_inst_pe_1_6_4_n90, npu_inst_pe_1_6_4_n89, npu_inst_pe_1_6_4_n88,
         npu_inst_pe_1_6_4_n87, npu_inst_pe_1_6_4_n86, npu_inst_pe_1_6_4_n85,
         npu_inst_pe_1_6_4_n84, npu_inst_pe_1_6_4_n83, npu_inst_pe_1_6_4_n82,
         npu_inst_pe_1_6_4_n81, npu_inst_pe_1_6_4_n80, npu_inst_pe_1_6_4_n79,
         npu_inst_pe_1_6_4_n78, npu_inst_pe_1_6_4_n77, npu_inst_pe_1_6_4_n76,
         npu_inst_pe_1_6_4_n75, npu_inst_pe_1_6_4_n74, npu_inst_pe_1_6_4_n73,
         npu_inst_pe_1_6_4_n72, npu_inst_pe_1_6_4_n71, npu_inst_pe_1_6_4_n70,
         npu_inst_pe_1_6_4_n69, npu_inst_pe_1_6_4_n68, npu_inst_pe_1_6_4_n67,
         npu_inst_pe_1_6_4_n66, npu_inst_pe_1_6_4_n65, npu_inst_pe_1_6_4_n64,
         npu_inst_pe_1_6_4_n63, npu_inst_pe_1_6_4_n62, npu_inst_pe_1_6_4_n61,
         npu_inst_pe_1_6_4_n60, npu_inst_pe_1_6_4_n59, npu_inst_pe_1_6_4_n58,
         npu_inst_pe_1_6_4_n57, npu_inst_pe_1_6_4_n56, npu_inst_pe_1_6_4_n55,
         npu_inst_pe_1_6_4_n54, npu_inst_pe_1_6_4_n53, npu_inst_pe_1_6_4_n52,
         npu_inst_pe_1_6_4_n51, npu_inst_pe_1_6_4_n50, npu_inst_pe_1_6_4_n49,
         npu_inst_pe_1_6_4_n48, npu_inst_pe_1_6_4_n47, npu_inst_pe_1_6_4_n46,
         npu_inst_pe_1_6_4_n45, npu_inst_pe_1_6_4_n44, npu_inst_pe_1_6_4_n43,
         npu_inst_pe_1_6_4_n42, npu_inst_pe_1_6_4_n41, npu_inst_pe_1_6_4_n40,
         npu_inst_pe_1_6_4_n39, npu_inst_pe_1_6_4_n38, npu_inst_pe_1_6_4_n37,
         npu_inst_pe_1_6_4_n27, npu_inst_pe_1_6_4_n26,
         npu_inst_pe_1_6_4_net3288, npu_inst_pe_1_6_4_net3282,
         npu_inst_pe_1_6_4_N94, npu_inst_pe_1_6_4_N93, npu_inst_pe_1_6_4_N84,
         npu_inst_pe_1_6_4_N80, npu_inst_pe_1_6_4_N79, npu_inst_pe_1_6_4_N78,
         npu_inst_pe_1_6_4_N77, npu_inst_pe_1_6_4_N76, npu_inst_pe_1_6_4_N75,
         npu_inst_pe_1_6_4_N74, npu_inst_pe_1_6_4_N73, npu_inst_pe_1_6_4_N72,
         npu_inst_pe_1_6_4_N71, npu_inst_pe_1_6_4_N70, npu_inst_pe_1_6_4_N69,
         npu_inst_pe_1_6_4_N68, npu_inst_pe_1_6_4_N67, npu_inst_pe_1_6_4_N66,
         npu_inst_pe_1_6_4_N65, npu_inst_pe_1_6_4_int_data_0_,
         npu_inst_pe_1_6_4_int_data_1_, npu_inst_pe_1_6_4_int_q_weight_0_,
         npu_inst_pe_1_6_4_int_q_weight_1_,
         npu_inst_pe_1_6_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_4_int_q_reg_h_0__1_, npu_inst_pe_1_6_5_n118,
         npu_inst_pe_1_6_5_n117, npu_inst_pe_1_6_5_n116,
         npu_inst_pe_1_6_5_n115, npu_inst_pe_1_6_5_n114,
         npu_inst_pe_1_6_5_n113, npu_inst_pe_1_6_5_n112,
         npu_inst_pe_1_6_5_n111, npu_inst_pe_1_6_5_n110,
         npu_inst_pe_1_6_5_n109, npu_inst_pe_1_6_5_n108,
         npu_inst_pe_1_6_5_n107, npu_inst_pe_1_6_5_n106,
         npu_inst_pe_1_6_5_n105, npu_inst_pe_1_6_5_n104,
         npu_inst_pe_1_6_5_n103, npu_inst_pe_1_6_5_n102,
         npu_inst_pe_1_6_5_n101, npu_inst_pe_1_6_5_n100, npu_inst_pe_1_6_5_n99,
         npu_inst_pe_1_6_5_n98, npu_inst_pe_1_6_5_n36, npu_inst_pe_1_6_5_n35,
         npu_inst_pe_1_6_5_n34, npu_inst_pe_1_6_5_n33, npu_inst_pe_1_6_5_n32,
         npu_inst_pe_1_6_5_n31, npu_inst_pe_1_6_5_n30, npu_inst_pe_1_6_5_n29,
         npu_inst_pe_1_6_5_n28, npu_inst_pe_1_6_5_n25, npu_inst_pe_1_6_5_n24,
         npu_inst_pe_1_6_5_n23, npu_inst_pe_1_6_5_n22, npu_inst_pe_1_6_5_n21,
         npu_inst_pe_1_6_5_n20, npu_inst_pe_1_6_5_n19, npu_inst_pe_1_6_5_n18,
         npu_inst_pe_1_6_5_n17, npu_inst_pe_1_6_5_n16, npu_inst_pe_1_6_5_n15,
         npu_inst_pe_1_6_5_n14, npu_inst_pe_1_6_5_n13, npu_inst_pe_1_6_5_n12,
         npu_inst_pe_1_6_5_n11, npu_inst_pe_1_6_5_n10, npu_inst_pe_1_6_5_n9,
         npu_inst_pe_1_6_5_n8, npu_inst_pe_1_6_5_n7, npu_inst_pe_1_6_5_n6,
         npu_inst_pe_1_6_5_n5, npu_inst_pe_1_6_5_n4, npu_inst_pe_1_6_5_n3,
         npu_inst_pe_1_6_5_n2, npu_inst_pe_1_6_5_n1,
         npu_inst_pe_1_6_5_sub_77_carry_7_, npu_inst_pe_1_6_5_sub_77_carry_6_,
         npu_inst_pe_1_6_5_sub_77_carry_5_, npu_inst_pe_1_6_5_sub_77_carry_4_,
         npu_inst_pe_1_6_5_sub_77_carry_3_, npu_inst_pe_1_6_5_sub_77_carry_2_,
         npu_inst_pe_1_6_5_sub_77_carry_1_, npu_inst_pe_1_6_5_add_79_carry_7_,
         npu_inst_pe_1_6_5_add_79_carry_6_, npu_inst_pe_1_6_5_add_79_carry_5_,
         npu_inst_pe_1_6_5_add_79_carry_4_, npu_inst_pe_1_6_5_add_79_carry_3_,
         npu_inst_pe_1_6_5_add_79_carry_2_, npu_inst_pe_1_6_5_add_79_carry_1_,
         npu_inst_pe_1_6_5_n97, npu_inst_pe_1_6_5_n96, npu_inst_pe_1_6_5_n95,
         npu_inst_pe_1_6_5_n94, npu_inst_pe_1_6_5_n93, npu_inst_pe_1_6_5_n92,
         npu_inst_pe_1_6_5_n91, npu_inst_pe_1_6_5_n90, npu_inst_pe_1_6_5_n89,
         npu_inst_pe_1_6_5_n88, npu_inst_pe_1_6_5_n87, npu_inst_pe_1_6_5_n86,
         npu_inst_pe_1_6_5_n85, npu_inst_pe_1_6_5_n84, npu_inst_pe_1_6_5_n83,
         npu_inst_pe_1_6_5_n82, npu_inst_pe_1_6_5_n81, npu_inst_pe_1_6_5_n80,
         npu_inst_pe_1_6_5_n79, npu_inst_pe_1_6_5_n78, npu_inst_pe_1_6_5_n77,
         npu_inst_pe_1_6_5_n76, npu_inst_pe_1_6_5_n75, npu_inst_pe_1_6_5_n74,
         npu_inst_pe_1_6_5_n73, npu_inst_pe_1_6_5_n72, npu_inst_pe_1_6_5_n71,
         npu_inst_pe_1_6_5_n70, npu_inst_pe_1_6_5_n69, npu_inst_pe_1_6_5_n68,
         npu_inst_pe_1_6_5_n67, npu_inst_pe_1_6_5_n66, npu_inst_pe_1_6_5_n65,
         npu_inst_pe_1_6_5_n64, npu_inst_pe_1_6_5_n63, npu_inst_pe_1_6_5_n62,
         npu_inst_pe_1_6_5_n61, npu_inst_pe_1_6_5_n60, npu_inst_pe_1_6_5_n59,
         npu_inst_pe_1_6_5_n58, npu_inst_pe_1_6_5_n57, npu_inst_pe_1_6_5_n56,
         npu_inst_pe_1_6_5_n55, npu_inst_pe_1_6_5_n54, npu_inst_pe_1_6_5_n53,
         npu_inst_pe_1_6_5_n52, npu_inst_pe_1_6_5_n51, npu_inst_pe_1_6_5_n50,
         npu_inst_pe_1_6_5_n49, npu_inst_pe_1_6_5_n48, npu_inst_pe_1_6_5_n47,
         npu_inst_pe_1_6_5_n46, npu_inst_pe_1_6_5_n45, npu_inst_pe_1_6_5_n44,
         npu_inst_pe_1_6_5_n43, npu_inst_pe_1_6_5_n42, npu_inst_pe_1_6_5_n41,
         npu_inst_pe_1_6_5_n40, npu_inst_pe_1_6_5_n39, npu_inst_pe_1_6_5_n38,
         npu_inst_pe_1_6_5_n37, npu_inst_pe_1_6_5_n27, npu_inst_pe_1_6_5_n26,
         npu_inst_pe_1_6_5_net3265, npu_inst_pe_1_6_5_net3259,
         npu_inst_pe_1_6_5_N94, npu_inst_pe_1_6_5_N93, npu_inst_pe_1_6_5_N84,
         npu_inst_pe_1_6_5_N80, npu_inst_pe_1_6_5_N79, npu_inst_pe_1_6_5_N78,
         npu_inst_pe_1_6_5_N77, npu_inst_pe_1_6_5_N76, npu_inst_pe_1_6_5_N75,
         npu_inst_pe_1_6_5_N74, npu_inst_pe_1_6_5_N73, npu_inst_pe_1_6_5_N72,
         npu_inst_pe_1_6_5_N71, npu_inst_pe_1_6_5_N70, npu_inst_pe_1_6_5_N69,
         npu_inst_pe_1_6_5_N68, npu_inst_pe_1_6_5_N67, npu_inst_pe_1_6_5_N66,
         npu_inst_pe_1_6_5_N65, npu_inst_pe_1_6_5_int_data_0_,
         npu_inst_pe_1_6_5_int_data_1_, npu_inst_pe_1_6_5_int_q_weight_0_,
         npu_inst_pe_1_6_5_int_q_weight_1_,
         npu_inst_pe_1_6_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_5_int_q_reg_h_0__1_, npu_inst_pe_1_6_6_n118,
         npu_inst_pe_1_6_6_n117, npu_inst_pe_1_6_6_n116,
         npu_inst_pe_1_6_6_n115, npu_inst_pe_1_6_6_n114,
         npu_inst_pe_1_6_6_n113, npu_inst_pe_1_6_6_n112,
         npu_inst_pe_1_6_6_n111, npu_inst_pe_1_6_6_n110,
         npu_inst_pe_1_6_6_n109, npu_inst_pe_1_6_6_n108,
         npu_inst_pe_1_6_6_n107, npu_inst_pe_1_6_6_n106,
         npu_inst_pe_1_6_6_n105, npu_inst_pe_1_6_6_n104,
         npu_inst_pe_1_6_6_n103, npu_inst_pe_1_6_6_n102,
         npu_inst_pe_1_6_6_n101, npu_inst_pe_1_6_6_n100, npu_inst_pe_1_6_6_n99,
         npu_inst_pe_1_6_6_n98, npu_inst_pe_1_6_6_n36, npu_inst_pe_1_6_6_n35,
         npu_inst_pe_1_6_6_n34, npu_inst_pe_1_6_6_n33, npu_inst_pe_1_6_6_n32,
         npu_inst_pe_1_6_6_n31, npu_inst_pe_1_6_6_n30, npu_inst_pe_1_6_6_n29,
         npu_inst_pe_1_6_6_n28, npu_inst_pe_1_6_6_n25, npu_inst_pe_1_6_6_n24,
         npu_inst_pe_1_6_6_n23, npu_inst_pe_1_6_6_n22, npu_inst_pe_1_6_6_n21,
         npu_inst_pe_1_6_6_n20, npu_inst_pe_1_6_6_n19, npu_inst_pe_1_6_6_n18,
         npu_inst_pe_1_6_6_n17, npu_inst_pe_1_6_6_n16, npu_inst_pe_1_6_6_n15,
         npu_inst_pe_1_6_6_n14, npu_inst_pe_1_6_6_n13, npu_inst_pe_1_6_6_n12,
         npu_inst_pe_1_6_6_n11, npu_inst_pe_1_6_6_n10, npu_inst_pe_1_6_6_n9,
         npu_inst_pe_1_6_6_n8, npu_inst_pe_1_6_6_n7, npu_inst_pe_1_6_6_n6,
         npu_inst_pe_1_6_6_n5, npu_inst_pe_1_6_6_n4, npu_inst_pe_1_6_6_n3,
         npu_inst_pe_1_6_6_n2, npu_inst_pe_1_6_6_n1,
         npu_inst_pe_1_6_6_sub_77_carry_7_, npu_inst_pe_1_6_6_sub_77_carry_6_,
         npu_inst_pe_1_6_6_sub_77_carry_5_, npu_inst_pe_1_6_6_sub_77_carry_4_,
         npu_inst_pe_1_6_6_sub_77_carry_3_, npu_inst_pe_1_6_6_sub_77_carry_2_,
         npu_inst_pe_1_6_6_sub_77_carry_1_, npu_inst_pe_1_6_6_add_79_carry_7_,
         npu_inst_pe_1_6_6_add_79_carry_6_, npu_inst_pe_1_6_6_add_79_carry_5_,
         npu_inst_pe_1_6_6_add_79_carry_4_, npu_inst_pe_1_6_6_add_79_carry_3_,
         npu_inst_pe_1_6_6_add_79_carry_2_, npu_inst_pe_1_6_6_add_79_carry_1_,
         npu_inst_pe_1_6_6_n97, npu_inst_pe_1_6_6_n96, npu_inst_pe_1_6_6_n95,
         npu_inst_pe_1_6_6_n94, npu_inst_pe_1_6_6_n93, npu_inst_pe_1_6_6_n92,
         npu_inst_pe_1_6_6_n91, npu_inst_pe_1_6_6_n90, npu_inst_pe_1_6_6_n89,
         npu_inst_pe_1_6_6_n88, npu_inst_pe_1_6_6_n87, npu_inst_pe_1_6_6_n86,
         npu_inst_pe_1_6_6_n85, npu_inst_pe_1_6_6_n84, npu_inst_pe_1_6_6_n83,
         npu_inst_pe_1_6_6_n82, npu_inst_pe_1_6_6_n81, npu_inst_pe_1_6_6_n80,
         npu_inst_pe_1_6_6_n79, npu_inst_pe_1_6_6_n78, npu_inst_pe_1_6_6_n77,
         npu_inst_pe_1_6_6_n76, npu_inst_pe_1_6_6_n75, npu_inst_pe_1_6_6_n74,
         npu_inst_pe_1_6_6_n73, npu_inst_pe_1_6_6_n72, npu_inst_pe_1_6_6_n71,
         npu_inst_pe_1_6_6_n70, npu_inst_pe_1_6_6_n69, npu_inst_pe_1_6_6_n68,
         npu_inst_pe_1_6_6_n67, npu_inst_pe_1_6_6_n66, npu_inst_pe_1_6_6_n65,
         npu_inst_pe_1_6_6_n64, npu_inst_pe_1_6_6_n63, npu_inst_pe_1_6_6_n62,
         npu_inst_pe_1_6_6_n61, npu_inst_pe_1_6_6_n60, npu_inst_pe_1_6_6_n59,
         npu_inst_pe_1_6_6_n58, npu_inst_pe_1_6_6_n57, npu_inst_pe_1_6_6_n56,
         npu_inst_pe_1_6_6_n55, npu_inst_pe_1_6_6_n54, npu_inst_pe_1_6_6_n53,
         npu_inst_pe_1_6_6_n52, npu_inst_pe_1_6_6_n51, npu_inst_pe_1_6_6_n50,
         npu_inst_pe_1_6_6_n49, npu_inst_pe_1_6_6_n48, npu_inst_pe_1_6_6_n47,
         npu_inst_pe_1_6_6_n46, npu_inst_pe_1_6_6_n45, npu_inst_pe_1_6_6_n44,
         npu_inst_pe_1_6_6_n43, npu_inst_pe_1_6_6_n42, npu_inst_pe_1_6_6_n41,
         npu_inst_pe_1_6_6_n40, npu_inst_pe_1_6_6_n39, npu_inst_pe_1_6_6_n38,
         npu_inst_pe_1_6_6_n37, npu_inst_pe_1_6_6_n27, npu_inst_pe_1_6_6_n26,
         npu_inst_pe_1_6_6_net3242, npu_inst_pe_1_6_6_net3236,
         npu_inst_pe_1_6_6_N94, npu_inst_pe_1_6_6_N93, npu_inst_pe_1_6_6_N84,
         npu_inst_pe_1_6_6_N80, npu_inst_pe_1_6_6_N79, npu_inst_pe_1_6_6_N78,
         npu_inst_pe_1_6_6_N77, npu_inst_pe_1_6_6_N76, npu_inst_pe_1_6_6_N75,
         npu_inst_pe_1_6_6_N74, npu_inst_pe_1_6_6_N73, npu_inst_pe_1_6_6_N72,
         npu_inst_pe_1_6_6_N71, npu_inst_pe_1_6_6_N70, npu_inst_pe_1_6_6_N69,
         npu_inst_pe_1_6_6_N68, npu_inst_pe_1_6_6_N67, npu_inst_pe_1_6_6_N66,
         npu_inst_pe_1_6_6_N65, npu_inst_pe_1_6_6_int_data_0_,
         npu_inst_pe_1_6_6_int_data_1_, npu_inst_pe_1_6_6_int_q_weight_0_,
         npu_inst_pe_1_6_6_int_q_weight_1_,
         npu_inst_pe_1_6_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_6_int_q_reg_h_0__1_, npu_inst_pe_1_6_7_n118,
         npu_inst_pe_1_6_7_n117, npu_inst_pe_1_6_7_n116,
         npu_inst_pe_1_6_7_n115, npu_inst_pe_1_6_7_n114,
         npu_inst_pe_1_6_7_n113, npu_inst_pe_1_6_7_n112,
         npu_inst_pe_1_6_7_n111, npu_inst_pe_1_6_7_n110,
         npu_inst_pe_1_6_7_n109, npu_inst_pe_1_6_7_n108,
         npu_inst_pe_1_6_7_n107, npu_inst_pe_1_6_7_n106,
         npu_inst_pe_1_6_7_n105, npu_inst_pe_1_6_7_n104,
         npu_inst_pe_1_6_7_n103, npu_inst_pe_1_6_7_n102,
         npu_inst_pe_1_6_7_n101, npu_inst_pe_1_6_7_n100, npu_inst_pe_1_6_7_n99,
         npu_inst_pe_1_6_7_n98, npu_inst_pe_1_6_7_n36, npu_inst_pe_1_6_7_n35,
         npu_inst_pe_1_6_7_n34, npu_inst_pe_1_6_7_n33, npu_inst_pe_1_6_7_n32,
         npu_inst_pe_1_6_7_n31, npu_inst_pe_1_6_7_n30, npu_inst_pe_1_6_7_n29,
         npu_inst_pe_1_6_7_n28, npu_inst_pe_1_6_7_n25, npu_inst_pe_1_6_7_n24,
         npu_inst_pe_1_6_7_n23, npu_inst_pe_1_6_7_n22, npu_inst_pe_1_6_7_n21,
         npu_inst_pe_1_6_7_n20, npu_inst_pe_1_6_7_n19, npu_inst_pe_1_6_7_n18,
         npu_inst_pe_1_6_7_n17, npu_inst_pe_1_6_7_n16, npu_inst_pe_1_6_7_n15,
         npu_inst_pe_1_6_7_n14, npu_inst_pe_1_6_7_n13, npu_inst_pe_1_6_7_n12,
         npu_inst_pe_1_6_7_n11, npu_inst_pe_1_6_7_n10, npu_inst_pe_1_6_7_n9,
         npu_inst_pe_1_6_7_n8, npu_inst_pe_1_6_7_n7, npu_inst_pe_1_6_7_n6,
         npu_inst_pe_1_6_7_n5, npu_inst_pe_1_6_7_n4, npu_inst_pe_1_6_7_n3,
         npu_inst_pe_1_6_7_n2, npu_inst_pe_1_6_7_n1,
         npu_inst_pe_1_6_7_sub_77_carry_7_, npu_inst_pe_1_6_7_sub_77_carry_6_,
         npu_inst_pe_1_6_7_sub_77_carry_5_, npu_inst_pe_1_6_7_sub_77_carry_4_,
         npu_inst_pe_1_6_7_sub_77_carry_3_, npu_inst_pe_1_6_7_sub_77_carry_2_,
         npu_inst_pe_1_6_7_sub_77_carry_1_, npu_inst_pe_1_6_7_add_79_carry_7_,
         npu_inst_pe_1_6_7_add_79_carry_6_, npu_inst_pe_1_6_7_add_79_carry_5_,
         npu_inst_pe_1_6_7_add_79_carry_4_, npu_inst_pe_1_6_7_add_79_carry_3_,
         npu_inst_pe_1_6_7_add_79_carry_2_, npu_inst_pe_1_6_7_add_79_carry_1_,
         npu_inst_pe_1_6_7_n97, npu_inst_pe_1_6_7_n96, npu_inst_pe_1_6_7_n95,
         npu_inst_pe_1_6_7_n94, npu_inst_pe_1_6_7_n93, npu_inst_pe_1_6_7_n92,
         npu_inst_pe_1_6_7_n91, npu_inst_pe_1_6_7_n90, npu_inst_pe_1_6_7_n89,
         npu_inst_pe_1_6_7_n88, npu_inst_pe_1_6_7_n87, npu_inst_pe_1_6_7_n86,
         npu_inst_pe_1_6_7_n85, npu_inst_pe_1_6_7_n84, npu_inst_pe_1_6_7_n83,
         npu_inst_pe_1_6_7_n82, npu_inst_pe_1_6_7_n81, npu_inst_pe_1_6_7_n80,
         npu_inst_pe_1_6_7_n79, npu_inst_pe_1_6_7_n78, npu_inst_pe_1_6_7_n77,
         npu_inst_pe_1_6_7_n76, npu_inst_pe_1_6_7_n75, npu_inst_pe_1_6_7_n74,
         npu_inst_pe_1_6_7_n73, npu_inst_pe_1_6_7_n72, npu_inst_pe_1_6_7_n71,
         npu_inst_pe_1_6_7_n70, npu_inst_pe_1_6_7_n69, npu_inst_pe_1_6_7_n68,
         npu_inst_pe_1_6_7_n67, npu_inst_pe_1_6_7_n66, npu_inst_pe_1_6_7_n65,
         npu_inst_pe_1_6_7_n64, npu_inst_pe_1_6_7_n63, npu_inst_pe_1_6_7_n62,
         npu_inst_pe_1_6_7_n61, npu_inst_pe_1_6_7_n60, npu_inst_pe_1_6_7_n59,
         npu_inst_pe_1_6_7_n58, npu_inst_pe_1_6_7_n57, npu_inst_pe_1_6_7_n56,
         npu_inst_pe_1_6_7_n55, npu_inst_pe_1_6_7_n54, npu_inst_pe_1_6_7_n53,
         npu_inst_pe_1_6_7_n52, npu_inst_pe_1_6_7_n51, npu_inst_pe_1_6_7_n50,
         npu_inst_pe_1_6_7_n49, npu_inst_pe_1_6_7_n48, npu_inst_pe_1_6_7_n47,
         npu_inst_pe_1_6_7_n46, npu_inst_pe_1_6_7_n45, npu_inst_pe_1_6_7_n44,
         npu_inst_pe_1_6_7_n43, npu_inst_pe_1_6_7_n42, npu_inst_pe_1_6_7_n41,
         npu_inst_pe_1_6_7_n40, npu_inst_pe_1_6_7_n39, npu_inst_pe_1_6_7_n38,
         npu_inst_pe_1_6_7_n37, npu_inst_pe_1_6_7_n27, npu_inst_pe_1_6_7_n26,
         npu_inst_pe_1_6_7_net3219, npu_inst_pe_1_6_7_net3213,
         npu_inst_pe_1_6_7_N94, npu_inst_pe_1_6_7_N93, npu_inst_pe_1_6_7_N84,
         npu_inst_pe_1_6_7_N80, npu_inst_pe_1_6_7_N79, npu_inst_pe_1_6_7_N78,
         npu_inst_pe_1_6_7_N77, npu_inst_pe_1_6_7_N76, npu_inst_pe_1_6_7_N75,
         npu_inst_pe_1_6_7_N74, npu_inst_pe_1_6_7_N73, npu_inst_pe_1_6_7_N72,
         npu_inst_pe_1_6_7_N71, npu_inst_pe_1_6_7_N70, npu_inst_pe_1_6_7_N69,
         npu_inst_pe_1_6_7_N68, npu_inst_pe_1_6_7_N67, npu_inst_pe_1_6_7_N66,
         npu_inst_pe_1_6_7_N65, npu_inst_pe_1_6_7_int_data_0_,
         npu_inst_pe_1_6_7_int_data_1_, npu_inst_pe_1_6_7_int_q_weight_0_,
         npu_inst_pe_1_6_7_int_q_weight_1_,
         npu_inst_pe_1_6_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_6_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_6_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_6_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_6_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_6_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_6_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_6_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_6_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_6_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_6_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_6_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_6_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_6_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_6_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_6_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_6_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_6_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_6_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_6_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_6_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_6_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_6_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_6_7_int_q_reg_h_0__1_, npu_inst_pe_1_7_0_n118,
         npu_inst_pe_1_7_0_n117, npu_inst_pe_1_7_0_n116,
         npu_inst_pe_1_7_0_n115, npu_inst_pe_1_7_0_n114,
         npu_inst_pe_1_7_0_n113, npu_inst_pe_1_7_0_n112,
         npu_inst_pe_1_7_0_n111, npu_inst_pe_1_7_0_n110,
         npu_inst_pe_1_7_0_n109, npu_inst_pe_1_7_0_n108,
         npu_inst_pe_1_7_0_n107, npu_inst_pe_1_7_0_n106,
         npu_inst_pe_1_7_0_n105, npu_inst_pe_1_7_0_n104,
         npu_inst_pe_1_7_0_n103, npu_inst_pe_1_7_0_n102,
         npu_inst_pe_1_7_0_n101, npu_inst_pe_1_7_0_n100, npu_inst_pe_1_7_0_n99,
         npu_inst_pe_1_7_0_n98, npu_inst_pe_1_7_0_n36, npu_inst_pe_1_7_0_n35,
         npu_inst_pe_1_7_0_n34, npu_inst_pe_1_7_0_n33, npu_inst_pe_1_7_0_n32,
         npu_inst_pe_1_7_0_n31, npu_inst_pe_1_7_0_n30, npu_inst_pe_1_7_0_n29,
         npu_inst_pe_1_7_0_n28, npu_inst_pe_1_7_0_n25, npu_inst_pe_1_7_0_n24,
         npu_inst_pe_1_7_0_n23, npu_inst_pe_1_7_0_n22, npu_inst_pe_1_7_0_n21,
         npu_inst_pe_1_7_0_n20, npu_inst_pe_1_7_0_n19, npu_inst_pe_1_7_0_n18,
         npu_inst_pe_1_7_0_n17, npu_inst_pe_1_7_0_n16, npu_inst_pe_1_7_0_n15,
         npu_inst_pe_1_7_0_n14, npu_inst_pe_1_7_0_n13, npu_inst_pe_1_7_0_n12,
         npu_inst_pe_1_7_0_n11, npu_inst_pe_1_7_0_n10, npu_inst_pe_1_7_0_n9,
         npu_inst_pe_1_7_0_n8, npu_inst_pe_1_7_0_n7, npu_inst_pe_1_7_0_n6,
         npu_inst_pe_1_7_0_n5, npu_inst_pe_1_7_0_n4, npu_inst_pe_1_7_0_n3,
         npu_inst_pe_1_7_0_n2, npu_inst_pe_1_7_0_n1,
         npu_inst_pe_1_7_0_sub_77_carry_7_, npu_inst_pe_1_7_0_sub_77_carry_6_,
         npu_inst_pe_1_7_0_sub_77_carry_5_, npu_inst_pe_1_7_0_sub_77_carry_4_,
         npu_inst_pe_1_7_0_sub_77_carry_3_, npu_inst_pe_1_7_0_sub_77_carry_2_,
         npu_inst_pe_1_7_0_sub_77_carry_1_, npu_inst_pe_1_7_0_add_79_carry_7_,
         npu_inst_pe_1_7_0_add_79_carry_6_, npu_inst_pe_1_7_0_add_79_carry_5_,
         npu_inst_pe_1_7_0_add_79_carry_4_, npu_inst_pe_1_7_0_add_79_carry_3_,
         npu_inst_pe_1_7_0_add_79_carry_2_, npu_inst_pe_1_7_0_add_79_carry_1_,
         npu_inst_pe_1_7_0_n97, npu_inst_pe_1_7_0_n96, npu_inst_pe_1_7_0_n95,
         npu_inst_pe_1_7_0_n94, npu_inst_pe_1_7_0_n93, npu_inst_pe_1_7_0_n92,
         npu_inst_pe_1_7_0_n91, npu_inst_pe_1_7_0_n90, npu_inst_pe_1_7_0_n89,
         npu_inst_pe_1_7_0_n88, npu_inst_pe_1_7_0_n87, npu_inst_pe_1_7_0_n86,
         npu_inst_pe_1_7_0_n85, npu_inst_pe_1_7_0_n84, npu_inst_pe_1_7_0_n83,
         npu_inst_pe_1_7_0_n82, npu_inst_pe_1_7_0_n81, npu_inst_pe_1_7_0_n80,
         npu_inst_pe_1_7_0_n79, npu_inst_pe_1_7_0_n78, npu_inst_pe_1_7_0_n77,
         npu_inst_pe_1_7_0_n76, npu_inst_pe_1_7_0_n75, npu_inst_pe_1_7_0_n74,
         npu_inst_pe_1_7_0_n73, npu_inst_pe_1_7_0_n72, npu_inst_pe_1_7_0_n71,
         npu_inst_pe_1_7_0_n70, npu_inst_pe_1_7_0_n69, npu_inst_pe_1_7_0_n68,
         npu_inst_pe_1_7_0_n67, npu_inst_pe_1_7_0_n66, npu_inst_pe_1_7_0_n65,
         npu_inst_pe_1_7_0_n64, npu_inst_pe_1_7_0_n63, npu_inst_pe_1_7_0_n62,
         npu_inst_pe_1_7_0_n61, npu_inst_pe_1_7_0_n60, npu_inst_pe_1_7_0_n59,
         npu_inst_pe_1_7_0_n58, npu_inst_pe_1_7_0_n57, npu_inst_pe_1_7_0_n56,
         npu_inst_pe_1_7_0_n55, npu_inst_pe_1_7_0_n54, npu_inst_pe_1_7_0_n53,
         npu_inst_pe_1_7_0_n52, npu_inst_pe_1_7_0_n51, npu_inst_pe_1_7_0_n50,
         npu_inst_pe_1_7_0_n49, npu_inst_pe_1_7_0_n48, npu_inst_pe_1_7_0_n47,
         npu_inst_pe_1_7_0_n46, npu_inst_pe_1_7_0_n45, npu_inst_pe_1_7_0_n44,
         npu_inst_pe_1_7_0_n43, npu_inst_pe_1_7_0_n42, npu_inst_pe_1_7_0_n41,
         npu_inst_pe_1_7_0_n40, npu_inst_pe_1_7_0_n39, npu_inst_pe_1_7_0_n38,
         npu_inst_pe_1_7_0_n37, npu_inst_pe_1_7_0_n27, npu_inst_pe_1_7_0_n26,
         npu_inst_pe_1_7_0_net3196, npu_inst_pe_1_7_0_net3190,
         npu_inst_pe_1_7_0_N94, npu_inst_pe_1_7_0_N93, npu_inst_pe_1_7_0_N84,
         npu_inst_pe_1_7_0_N80, npu_inst_pe_1_7_0_N79, npu_inst_pe_1_7_0_N78,
         npu_inst_pe_1_7_0_N77, npu_inst_pe_1_7_0_N76, npu_inst_pe_1_7_0_N75,
         npu_inst_pe_1_7_0_N74, npu_inst_pe_1_7_0_N73, npu_inst_pe_1_7_0_N72,
         npu_inst_pe_1_7_0_N71, npu_inst_pe_1_7_0_N70, npu_inst_pe_1_7_0_N69,
         npu_inst_pe_1_7_0_N68, npu_inst_pe_1_7_0_N67, npu_inst_pe_1_7_0_N66,
         npu_inst_pe_1_7_0_N65, npu_inst_pe_1_7_0_int_data_0_,
         npu_inst_pe_1_7_0_int_data_1_, npu_inst_pe_1_7_0_int_q_weight_0_,
         npu_inst_pe_1_7_0_int_q_weight_1_,
         npu_inst_pe_1_7_0_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_0_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_0_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_0_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_0_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_0_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_0_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_0_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_0_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_0_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_0_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_0_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_0_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_0_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_0_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_0_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_0_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_0_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_0_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_0_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_0_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_0_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_0_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_0_int_q_reg_h_0__1_, npu_inst_pe_1_7_0_o_data_h_0_,
         npu_inst_pe_1_7_0_o_data_h_1_, npu_inst_pe_1_7_1_n118,
         npu_inst_pe_1_7_1_n117, npu_inst_pe_1_7_1_n116,
         npu_inst_pe_1_7_1_n115, npu_inst_pe_1_7_1_n114,
         npu_inst_pe_1_7_1_n113, npu_inst_pe_1_7_1_n112,
         npu_inst_pe_1_7_1_n111, npu_inst_pe_1_7_1_n110,
         npu_inst_pe_1_7_1_n109, npu_inst_pe_1_7_1_n108,
         npu_inst_pe_1_7_1_n107, npu_inst_pe_1_7_1_n106,
         npu_inst_pe_1_7_1_n105, npu_inst_pe_1_7_1_n104,
         npu_inst_pe_1_7_1_n103, npu_inst_pe_1_7_1_n102,
         npu_inst_pe_1_7_1_n101, npu_inst_pe_1_7_1_n100, npu_inst_pe_1_7_1_n99,
         npu_inst_pe_1_7_1_n98, npu_inst_pe_1_7_1_n36, npu_inst_pe_1_7_1_n35,
         npu_inst_pe_1_7_1_n34, npu_inst_pe_1_7_1_n33, npu_inst_pe_1_7_1_n32,
         npu_inst_pe_1_7_1_n31, npu_inst_pe_1_7_1_n30, npu_inst_pe_1_7_1_n29,
         npu_inst_pe_1_7_1_n28, npu_inst_pe_1_7_1_n25, npu_inst_pe_1_7_1_n24,
         npu_inst_pe_1_7_1_n23, npu_inst_pe_1_7_1_n22, npu_inst_pe_1_7_1_n21,
         npu_inst_pe_1_7_1_n20, npu_inst_pe_1_7_1_n19, npu_inst_pe_1_7_1_n18,
         npu_inst_pe_1_7_1_n17, npu_inst_pe_1_7_1_n16, npu_inst_pe_1_7_1_n15,
         npu_inst_pe_1_7_1_n14, npu_inst_pe_1_7_1_n13, npu_inst_pe_1_7_1_n12,
         npu_inst_pe_1_7_1_n11, npu_inst_pe_1_7_1_n10, npu_inst_pe_1_7_1_n9,
         npu_inst_pe_1_7_1_n8, npu_inst_pe_1_7_1_n7, npu_inst_pe_1_7_1_n6,
         npu_inst_pe_1_7_1_n5, npu_inst_pe_1_7_1_n4, npu_inst_pe_1_7_1_n3,
         npu_inst_pe_1_7_1_n2, npu_inst_pe_1_7_1_n1,
         npu_inst_pe_1_7_1_sub_77_carry_7_, npu_inst_pe_1_7_1_sub_77_carry_6_,
         npu_inst_pe_1_7_1_sub_77_carry_5_, npu_inst_pe_1_7_1_sub_77_carry_4_,
         npu_inst_pe_1_7_1_sub_77_carry_3_, npu_inst_pe_1_7_1_sub_77_carry_2_,
         npu_inst_pe_1_7_1_sub_77_carry_1_, npu_inst_pe_1_7_1_add_79_carry_7_,
         npu_inst_pe_1_7_1_add_79_carry_6_, npu_inst_pe_1_7_1_add_79_carry_5_,
         npu_inst_pe_1_7_1_add_79_carry_4_, npu_inst_pe_1_7_1_add_79_carry_3_,
         npu_inst_pe_1_7_1_add_79_carry_2_, npu_inst_pe_1_7_1_add_79_carry_1_,
         npu_inst_pe_1_7_1_n97, npu_inst_pe_1_7_1_n96, npu_inst_pe_1_7_1_n95,
         npu_inst_pe_1_7_1_n94, npu_inst_pe_1_7_1_n93, npu_inst_pe_1_7_1_n92,
         npu_inst_pe_1_7_1_n91, npu_inst_pe_1_7_1_n90, npu_inst_pe_1_7_1_n89,
         npu_inst_pe_1_7_1_n88, npu_inst_pe_1_7_1_n87, npu_inst_pe_1_7_1_n86,
         npu_inst_pe_1_7_1_n85, npu_inst_pe_1_7_1_n84, npu_inst_pe_1_7_1_n83,
         npu_inst_pe_1_7_1_n82, npu_inst_pe_1_7_1_n81, npu_inst_pe_1_7_1_n80,
         npu_inst_pe_1_7_1_n79, npu_inst_pe_1_7_1_n78, npu_inst_pe_1_7_1_n77,
         npu_inst_pe_1_7_1_n76, npu_inst_pe_1_7_1_n75, npu_inst_pe_1_7_1_n74,
         npu_inst_pe_1_7_1_n73, npu_inst_pe_1_7_1_n72, npu_inst_pe_1_7_1_n71,
         npu_inst_pe_1_7_1_n70, npu_inst_pe_1_7_1_n69, npu_inst_pe_1_7_1_n68,
         npu_inst_pe_1_7_1_n67, npu_inst_pe_1_7_1_n66, npu_inst_pe_1_7_1_n65,
         npu_inst_pe_1_7_1_n64, npu_inst_pe_1_7_1_n63, npu_inst_pe_1_7_1_n62,
         npu_inst_pe_1_7_1_n61, npu_inst_pe_1_7_1_n60, npu_inst_pe_1_7_1_n59,
         npu_inst_pe_1_7_1_n58, npu_inst_pe_1_7_1_n57, npu_inst_pe_1_7_1_n56,
         npu_inst_pe_1_7_1_n55, npu_inst_pe_1_7_1_n54, npu_inst_pe_1_7_1_n53,
         npu_inst_pe_1_7_1_n52, npu_inst_pe_1_7_1_n51, npu_inst_pe_1_7_1_n50,
         npu_inst_pe_1_7_1_n49, npu_inst_pe_1_7_1_n48, npu_inst_pe_1_7_1_n47,
         npu_inst_pe_1_7_1_n46, npu_inst_pe_1_7_1_n45, npu_inst_pe_1_7_1_n44,
         npu_inst_pe_1_7_1_n43, npu_inst_pe_1_7_1_n42, npu_inst_pe_1_7_1_n41,
         npu_inst_pe_1_7_1_n40, npu_inst_pe_1_7_1_n39, npu_inst_pe_1_7_1_n38,
         npu_inst_pe_1_7_1_n37, npu_inst_pe_1_7_1_n27, npu_inst_pe_1_7_1_n26,
         npu_inst_pe_1_7_1_net3173, npu_inst_pe_1_7_1_net3167,
         npu_inst_pe_1_7_1_N94, npu_inst_pe_1_7_1_N93, npu_inst_pe_1_7_1_N84,
         npu_inst_pe_1_7_1_N80, npu_inst_pe_1_7_1_N79, npu_inst_pe_1_7_1_N78,
         npu_inst_pe_1_7_1_N77, npu_inst_pe_1_7_1_N76, npu_inst_pe_1_7_1_N75,
         npu_inst_pe_1_7_1_N74, npu_inst_pe_1_7_1_N73, npu_inst_pe_1_7_1_N72,
         npu_inst_pe_1_7_1_N71, npu_inst_pe_1_7_1_N70, npu_inst_pe_1_7_1_N69,
         npu_inst_pe_1_7_1_N68, npu_inst_pe_1_7_1_N67, npu_inst_pe_1_7_1_N66,
         npu_inst_pe_1_7_1_N65, npu_inst_pe_1_7_1_int_data_0_,
         npu_inst_pe_1_7_1_int_data_1_, npu_inst_pe_1_7_1_int_q_weight_0_,
         npu_inst_pe_1_7_1_int_q_weight_1_,
         npu_inst_pe_1_7_1_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_1_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_1_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_1_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_1_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_1_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_1_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_1_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_1_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_1_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_1_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_1_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_1_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_1_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_1_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_1_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_1_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_1_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_1_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_1_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_1_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_1_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_1_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_1_int_q_reg_h_0__1_, npu_inst_pe_1_7_2_n118,
         npu_inst_pe_1_7_2_n117, npu_inst_pe_1_7_2_n116,
         npu_inst_pe_1_7_2_n115, npu_inst_pe_1_7_2_n114,
         npu_inst_pe_1_7_2_n113, npu_inst_pe_1_7_2_n112,
         npu_inst_pe_1_7_2_n111, npu_inst_pe_1_7_2_n110,
         npu_inst_pe_1_7_2_n109, npu_inst_pe_1_7_2_n108,
         npu_inst_pe_1_7_2_n107, npu_inst_pe_1_7_2_n106,
         npu_inst_pe_1_7_2_n105, npu_inst_pe_1_7_2_n104,
         npu_inst_pe_1_7_2_n103, npu_inst_pe_1_7_2_n102,
         npu_inst_pe_1_7_2_n101, npu_inst_pe_1_7_2_n100, npu_inst_pe_1_7_2_n99,
         npu_inst_pe_1_7_2_n98, npu_inst_pe_1_7_2_n36, npu_inst_pe_1_7_2_n35,
         npu_inst_pe_1_7_2_n34, npu_inst_pe_1_7_2_n33, npu_inst_pe_1_7_2_n32,
         npu_inst_pe_1_7_2_n31, npu_inst_pe_1_7_2_n30, npu_inst_pe_1_7_2_n29,
         npu_inst_pe_1_7_2_n28, npu_inst_pe_1_7_2_n25, npu_inst_pe_1_7_2_n24,
         npu_inst_pe_1_7_2_n23, npu_inst_pe_1_7_2_n22, npu_inst_pe_1_7_2_n21,
         npu_inst_pe_1_7_2_n20, npu_inst_pe_1_7_2_n19, npu_inst_pe_1_7_2_n18,
         npu_inst_pe_1_7_2_n17, npu_inst_pe_1_7_2_n16, npu_inst_pe_1_7_2_n15,
         npu_inst_pe_1_7_2_n14, npu_inst_pe_1_7_2_n13, npu_inst_pe_1_7_2_n12,
         npu_inst_pe_1_7_2_n11, npu_inst_pe_1_7_2_n10, npu_inst_pe_1_7_2_n9,
         npu_inst_pe_1_7_2_n8, npu_inst_pe_1_7_2_n7, npu_inst_pe_1_7_2_n6,
         npu_inst_pe_1_7_2_n5, npu_inst_pe_1_7_2_n4, npu_inst_pe_1_7_2_n3,
         npu_inst_pe_1_7_2_n2, npu_inst_pe_1_7_2_n1,
         npu_inst_pe_1_7_2_sub_77_carry_7_, npu_inst_pe_1_7_2_sub_77_carry_6_,
         npu_inst_pe_1_7_2_sub_77_carry_5_, npu_inst_pe_1_7_2_sub_77_carry_4_,
         npu_inst_pe_1_7_2_sub_77_carry_3_, npu_inst_pe_1_7_2_sub_77_carry_2_,
         npu_inst_pe_1_7_2_sub_77_carry_1_, npu_inst_pe_1_7_2_add_79_carry_7_,
         npu_inst_pe_1_7_2_add_79_carry_6_, npu_inst_pe_1_7_2_add_79_carry_5_,
         npu_inst_pe_1_7_2_add_79_carry_4_, npu_inst_pe_1_7_2_add_79_carry_3_,
         npu_inst_pe_1_7_2_add_79_carry_2_, npu_inst_pe_1_7_2_add_79_carry_1_,
         npu_inst_pe_1_7_2_n97, npu_inst_pe_1_7_2_n96, npu_inst_pe_1_7_2_n95,
         npu_inst_pe_1_7_2_n94, npu_inst_pe_1_7_2_n93, npu_inst_pe_1_7_2_n92,
         npu_inst_pe_1_7_2_n91, npu_inst_pe_1_7_2_n90, npu_inst_pe_1_7_2_n89,
         npu_inst_pe_1_7_2_n88, npu_inst_pe_1_7_2_n87, npu_inst_pe_1_7_2_n86,
         npu_inst_pe_1_7_2_n85, npu_inst_pe_1_7_2_n84, npu_inst_pe_1_7_2_n83,
         npu_inst_pe_1_7_2_n82, npu_inst_pe_1_7_2_n81, npu_inst_pe_1_7_2_n80,
         npu_inst_pe_1_7_2_n79, npu_inst_pe_1_7_2_n78, npu_inst_pe_1_7_2_n77,
         npu_inst_pe_1_7_2_n76, npu_inst_pe_1_7_2_n75, npu_inst_pe_1_7_2_n74,
         npu_inst_pe_1_7_2_n73, npu_inst_pe_1_7_2_n72, npu_inst_pe_1_7_2_n71,
         npu_inst_pe_1_7_2_n70, npu_inst_pe_1_7_2_n69, npu_inst_pe_1_7_2_n68,
         npu_inst_pe_1_7_2_n67, npu_inst_pe_1_7_2_n66, npu_inst_pe_1_7_2_n65,
         npu_inst_pe_1_7_2_n64, npu_inst_pe_1_7_2_n63, npu_inst_pe_1_7_2_n62,
         npu_inst_pe_1_7_2_n61, npu_inst_pe_1_7_2_n60, npu_inst_pe_1_7_2_n59,
         npu_inst_pe_1_7_2_n58, npu_inst_pe_1_7_2_n57, npu_inst_pe_1_7_2_n56,
         npu_inst_pe_1_7_2_n55, npu_inst_pe_1_7_2_n54, npu_inst_pe_1_7_2_n53,
         npu_inst_pe_1_7_2_n52, npu_inst_pe_1_7_2_n51, npu_inst_pe_1_7_2_n50,
         npu_inst_pe_1_7_2_n49, npu_inst_pe_1_7_2_n48, npu_inst_pe_1_7_2_n47,
         npu_inst_pe_1_7_2_n46, npu_inst_pe_1_7_2_n45, npu_inst_pe_1_7_2_n44,
         npu_inst_pe_1_7_2_n43, npu_inst_pe_1_7_2_n42, npu_inst_pe_1_7_2_n41,
         npu_inst_pe_1_7_2_n40, npu_inst_pe_1_7_2_n39, npu_inst_pe_1_7_2_n38,
         npu_inst_pe_1_7_2_n37, npu_inst_pe_1_7_2_n27, npu_inst_pe_1_7_2_n26,
         npu_inst_pe_1_7_2_net3150, npu_inst_pe_1_7_2_net3144,
         npu_inst_pe_1_7_2_N94, npu_inst_pe_1_7_2_N93, npu_inst_pe_1_7_2_N84,
         npu_inst_pe_1_7_2_N80, npu_inst_pe_1_7_2_N79, npu_inst_pe_1_7_2_N78,
         npu_inst_pe_1_7_2_N77, npu_inst_pe_1_7_2_N76, npu_inst_pe_1_7_2_N75,
         npu_inst_pe_1_7_2_N74, npu_inst_pe_1_7_2_N73, npu_inst_pe_1_7_2_N72,
         npu_inst_pe_1_7_2_N71, npu_inst_pe_1_7_2_N70, npu_inst_pe_1_7_2_N69,
         npu_inst_pe_1_7_2_N68, npu_inst_pe_1_7_2_N67, npu_inst_pe_1_7_2_N66,
         npu_inst_pe_1_7_2_N65, npu_inst_pe_1_7_2_int_data_0_,
         npu_inst_pe_1_7_2_int_data_1_, npu_inst_pe_1_7_2_int_q_weight_0_,
         npu_inst_pe_1_7_2_int_q_weight_1_,
         npu_inst_pe_1_7_2_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_2_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_2_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_2_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_2_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_2_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_2_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_2_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_2_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_2_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_2_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_2_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_2_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_2_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_2_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_2_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_2_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_2_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_2_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_2_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_2_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_2_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_2_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_2_int_q_reg_h_0__1_, npu_inst_pe_1_7_3_n118,
         npu_inst_pe_1_7_3_n117, npu_inst_pe_1_7_3_n116,
         npu_inst_pe_1_7_3_n115, npu_inst_pe_1_7_3_n114,
         npu_inst_pe_1_7_3_n113, npu_inst_pe_1_7_3_n112,
         npu_inst_pe_1_7_3_n111, npu_inst_pe_1_7_3_n110,
         npu_inst_pe_1_7_3_n109, npu_inst_pe_1_7_3_n108,
         npu_inst_pe_1_7_3_n107, npu_inst_pe_1_7_3_n106,
         npu_inst_pe_1_7_3_n105, npu_inst_pe_1_7_3_n104,
         npu_inst_pe_1_7_3_n103, npu_inst_pe_1_7_3_n102,
         npu_inst_pe_1_7_3_n101, npu_inst_pe_1_7_3_n100, npu_inst_pe_1_7_3_n99,
         npu_inst_pe_1_7_3_n98, npu_inst_pe_1_7_3_n36, npu_inst_pe_1_7_3_n35,
         npu_inst_pe_1_7_3_n34, npu_inst_pe_1_7_3_n33, npu_inst_pe_1_7_3_n32,
         npu_inst_pe_1_7_3_n31, npu_inst_pe_1_7_3_n30, npu_inst_pe_1_7_3_n29,
         npu_inst_pe_1_7_3_n28, npu_inst_pe_1_7_3_n25, npu_inst_pe_1_7_3_n24,
         npu_inst_pe_1_7_3_n23, npu_inst_pe_1_7_3_n22, npu_inst_pe_1_7_3_n21,
         npu_inst_pe_1_7_3_n20, npu_inst_pe_1_7_3_n19, npu_inst_pe_1_7_3_n18,
         npu_inst_pe_1_7_3_n17, npu_inst_pe_1_7_3_n16, npu_inst_pe_1_7_3_n15,
         npu_inst_pe_1_7_3_n14, npu_inst_pe_1_7_3_n13, npu_inst_pe_1_7_3_n12,
         npu_inst_pe_1_7_3_n11, npu_inst_pe_1_7_3_n10, npu_inst_pe_1_7_3_n9,
         npu_inst_pe_1_7_3_n8, npu_inst_pe_1_7_3_n7, npu_inst_pe_1_7_3_n6,
         npu_inst_pe_1_7_3_n5, npu_inst_pe_1_7_3_n4, npu_inst_pe_1_7_3_n3,
         npu_inst_pe_1_7_3_n2, npu_inst_pe_1_7_3_n1,
         npu_inst_pe_1_7_3_sub_77_carry_7_, npu_inst_pe_1_7_3_sub_77_carry_6_,
         npu_inst_pe_1_7_3_sub_77_carry_5_, npu_inst_pe_1_7_3_sub_77_carry_4_,
         npu_inst_pe_1_7_3_sub_77_carry_3_, npu_inst_pe_1_7_3_sub_77_carry_2_,
         npu_inst_pe_1_7_3_sub_77_carry_1_, npu_inst_pe_1_7_3_add_79_carry_7_,
         npu_inst_pe_1_7_3_add_79_carry_6_, npu_inst_pe_1_7_3_add_79_carry_5_,
         npu_inst_pe_1_7_3_add_79_carry_4_, npu_inst_pe_1_7_3_add_79_carry_3_,
         npu_inst_pe_1_7_3_add_79_carry_2_, npu_inst_pe_1_7_3_add_79_carry_1_,
         npu_inst_pe_1_7_3_n97, npu_inst_pe_1_7_3_n96, npu_inst_pe_1_7_3_n95,
         npu_inst_pe_1_7_3_n94, npu_inst_pe_1_7_3_n93, npu_inst_pe_1_7_3_n92,
         npu_inst_pe_1_7_3_n91, npu_inst_pe_1_7_3_n90, npu_inst_pe_1_7_3_n89,
         npu_inst_pe_1_7_3_n88, npu_inst_pe_1_7_3_n87, npu_inst_pe_1_7_3_n86,
         npu_inst_pe_1_7_3_n85, npu_inst_pe_1_7_3_n84, npu_inst_pe_1_7_3_n83,
         npu_inst_pe_1_7_3_n82, npu_inst_pe_1_7_3_n81, npu_inst_pe_1_7_3_n80,
         npu_inst_pe_1_7_3_n79, npu_inst_pe_1_7_3_n78, npu_inst_pe_1_7_3_n77,
         npu_inst_pe_1_7_3_n76, npu_inst_pe_1_7_3_n75, npu_inst_pe_1_7_3_n74,
         npu_inst_pe_1_7_3_n73, npu_inst_pe_1_7_3_n72, npu_inst_pe_1_7_3_n71,
         npu_inst_pe_1_7_3_n70, npu_inst_pe_1_7_3_n69, npu_inst_pe_1_7_3_n68,
         npu_inst_pe_1_7_3_n67, npu_inst_pe_1_7_3_n66, npu_inst_pe_1_7_3_n65,
         npu_inst_pe_1_7_3_n64, npu_inst_pe_1_7_3_n63, npu_inst_pe_1_7_3_n62,
         npu_inst_pe_1_7_3_n61, npu_inst_pe_1_7_3_n60, npu_inst_pe_1_7_3_n59,
         npu_inst_pe_1_7_3_n58, npu_inst_pe_1_7_3_n57, npu_inst_pe_1_7_3_n56,
         npu_inst_pe_1_7_3_n55, npu_inst_pe_1_7_3_n54, npu_inst_pe_1_7_3_n53,
         npu_inst_pe_1_7_3_n52, npu_inst_pe_1_7_3_n51, npu_inst_pe_1_7_3_n50,
         npu_inst_pe_1_7_3_n49, npu_inst_pe_1_7_3_n48, npu_inst_pe_1_7_3_n47,
         npu_inst_pe_1_7_3_n46, npu_inst_pe_1_7_3_n45, npu_inst_pe_1_7_3_n44,
         npu_inst_pe_1_7_3_n43, npu_inst_pe_1_7_3_n42, npu_inst_pe_1_7_3_n41,
         npu_inst_pe_1_7_3_n40, npu_inst_pe_1_7_3_n39, npu_inst_pe_1_7_3_n38,
         npu_inst_pe_1_7_3_n37, npu_inst_pe_1_7_3_n27, npu_inst_pe_1_7_3_n26,
         npu_inst_pe_1_7_3_net3127, npu_inst_pe_1_7_3_net3121,
         npu_inst_pe_1_7_3_N94, npu_inst_pe_1_7_3_N93, npu_inst_pe_1_7_3_N84,
         npu_inst_pe_1_7_3_N80, npu_inst_pe_1_7_3_N79, npu_inst_pe_1_7_3_N78,
         npu_inst_pe_1_7_3_N77, npu_inst_pe_1_7_3_N76, npu_inst_pe_1_7_3_N75,
         npu_inst_pe_1_7_3_N74, npu_inst_pe_1_7_3_N73, npu_inst_pe_1_7_3_N72,
         npu_inst_pe_1_7_3_N71, npu_inst_pe_1_7_3_N70, npu_inst_pe_1_7_3_N69,
         npu_inst_pe_1_7_3_N68, npu_inst_pe_1_7_3_N67, npu_inst_pe_1_7_3_N66,
         npu_inst_pe_1_7_3_N65, npu_inst_pe_1_7_3_int_data_0_,
         npu_inst_pe_1_7_3_int_data_1_, npu_inst_pe_1_7_3_int_q_weight_0_,
         npu_inst_pe_1_7_3_int_q_weight_1_,
         npu_inst_pe_1_7_3_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_3_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_3_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_3_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_3_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_3_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_3_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_3_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_3_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_3_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_3_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_3_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_3_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_3_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_3_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_3_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_3_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_3_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_3_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_3_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_3_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_3_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_3_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_3_int_q_reg_h_0__1_, npu_inst_pe_1_7_4_n118,
         npu_inst_pe_1_7_4_n117, npu_inst_pe_1_7_4_n116,
         npu_inst_pe_1_7_4_n115, npu_inst_pe_1_7_4_n114,
         npu_inst_pe_1_7_4_n113, npu_inst_pe_1_7_4_n112,
         npu_inst_pe_1_7_4_n111, npu_inst_pe_1_7_4_n110,
         npu_inst_pe_1_7_4_n109, npu_inst_pe_1_7_4_n108,
         npu_inst_pe_1_7_4_n107, npu_inst_pe_1_7_4_n106,
         npu_inst_pe_1_7_4_n105, npu_inst_pe_1_7_4_n104,
         npu_inst_pe_1_7_4_n103, npu_inst_pe_1_7_4_n102,
         npu_inst_pe_1_7_4_n101, npu_inst_pe_1_7_4_n100, npu_inst_pe_1_7_4_n99,
         npu_inst_pe_1_7_4_n98, npu_inst_pe_1_7_4_n36, npu_inst_pe_1_7_4_n35,
         npu_inst_pe_1_7_4_n34, npu_inst_pe_1_7_4_n33, npu_inst_pe_1_7_4_n32,
         npu_inst_pe_1_7_4_n31, npu_inst_pe_1_7_4_n30, npu_inst_pe_1_7_4_n29,
         npu_inst_pe_1_7_4_n28, npu_inst_pe_1_7_4_n25, npu_inst_pe_1_7_4_n24,
         npu_inst_pe_1_7_4_n23, npu_inst_pe_1_7_4_n22, npu_inst_pe_1_7_4_n21,
         npu_inst_pe_1_7_4_n20, npu_inst_pe_1_7_4_n19, npu_inst_pe_1_7_4_n18,
         npu_inst_pe_1_7_4_n17, npu_inst_pe_1_7_4_n16, npu_inst_pe_1_7_4_n15,
         npu_inst_pe_1_7_4_n14, npu_inst_pe_1_7_4_n13, npu_inst_pe_1_7_4_n12,
         npu_inst_pe_1_7_4_n11, npu_inst_pe_1_7_4_n10, npu_inst_pe_1_7_4_n9,
         npu_inst_pe_1_7_4_n8, npu_inst_pe_1_7_4_n7, npu_inst_pe_1_7_4_n6,
         npu_inst_pe_1_7_4_n5, npu_inst_pe_1_7_4_n4, npu_inst_pe_1_7_4_n3,
         npu_inst_pe_1_7_4_n2, npu_inst_pe_1_7_4_n1,
         npu_inst_pe_1_7_4_sub_77_carry_7_, npu_inst_pe_1_7_4_sub_77_carry_6_,
         npu_inst_pe_1_7_4_sub_77_carry_5_, npu_inst_pe_1_7_4_sub_77_carry_4_,
         npu_inst_pe_1_7_4_sub_77_carry_3_, npu_inst_pe_1_7_4_sub_77_carry_2_,
         npu_inst_pe_1_7_4_sub_77_carry_1_, npu_inst_pe_1_7_4_add_79_carry_7_,
         npu_inst_pe_1_7_4_add_79_carry_6_, npu_inst_pe_1_7_4_add_79_carry_5_,
         npu_inst_pe_1_7_4_add_79_carry_4_, npu_inst_pe_1_7_4_add_79_carry_3_,
         npu_inst_pe_1_7_4_add_79_carry_2_, npu_inst_pe_1_7_4_add_79_carry_1_,
         npu_inst_pe_1_7_4_n97, npu_inst_pe_1_7_4_n96, npu_inst_pe_1_7_4_n95,
         npu_inst_pe_1_7_4_n94, npu_inst_pe_1_7_4_n93, npu_inst_pe_1_7_4_n92,
         npu_inst_pe_1_7_4_n91, npu_inst_pe_1_7_4_n90, npu_inst_pe_1_7_4_n89,
         npu_inst_pe_1_7_4_n88, npu_inst_pe_1_7_4_n87, npu_inst_pe_1_7_4_n86,
         npu_inst_pe_1_7_4_n85, npu_inst_pe_1_7_4_n84, npu_inst_pe_1_7_4_n83,
         npu_inst_pe_1_7_4_n82, npu_inst_pe_1_7_4_n81, npu_inst_pe_1_7_4_n80,
         npu_inst_pe_1_7_4_n79, npu_inst_pe_1_7_4_n78, npu_inst_pe_1_7_4_n77,
         npu_inst_pe_1_7_4_n76, npu_inst_pe_1_7_4_n75, npu_inst_pe_1_7_4_n74,
         npu_inst_pe_1_7_4_n73, npu_inst_pe_1_7_4_n72, npu_inst_pe_1_7_4_n71,
         npu_inst_pe_1_7_4_n70, npu_inst_pe_1_7_4_n69, npu_inst_pe_1_7_4_n68,
         npu_inst_pe_1_7_4_n67, npu_inst_pe_1_7_4_n66, npu_inst_pe_1_7_4_n65,
         npu_inst_pe_1_7_4_n64, npu_inst_pe_1_7_4_n63, npu_inst_pe_1_7_4_n62,
         npu_inst_pe_1_7_4_n61, npu_inst_pe_1_7_4_n60, npu_inst_pe_1_7_4_n59,
         npu_inst_pe_1_7_4_n58, npu_inst_pe_1_7_4_n57, npu_inst_pe_1_7_4_n56,
         npu_inst_pe_1_7_4_n55, npu_inst_pe_1_7_4_n54, npu_inst_pe_1_7_4_n53,
         npu_inst_pe_1_7_4_n52, npu_inst_pe_1_7_4_n51, npu_inst_pe_1_7_4_n50,
         npu_inst_pe_1_7_4_n49, npu_inst_pe_1_7_4_n48, npu_inst_pe_1_7_4_n47,
         npu_inst_pe_1_7_4_n46, npu_inst_pe_1_7_4_n45, npu_inst_pe_1_7_4_n44,
         npu_inst_pe_1_7_4_n43, npu_inst_pe_1_7_4_n42, npu_inst_pe_1_7_4_n41,
         npu_inst_pe_1_7_4_n40, npu_inst_pe_1_7_4_n39, npu_inst_pe_1_7_4_n38,
         npu_inst_pe_1_7_4_n37, npu_inst_pe_1_7_4_n27, npu_inst_pe_1_7_4_n26,
         npu_inst_pe_1_7_4_net3104, npu_inst_pe_1_7_4_net3098,
         npu_inst_pe_1_7_4_N94, npu_inst_pe_1_7_4_N93, npu_inst_pe_1_7_4_N84,
         npu_inst_pe_1_7_4_N80, npu_inst_pe_1_7_4_N79, npu_inst_pe_1_7_4_N78,
         npu_inst_pe_1_7_4_N77, npu_inst_pe_1_7_4_N76, npu_inst_pe_1_7_4_N75,
         npu_inst_pe_1_7_4_N74, npu_inst_pe_1_7_4_N73, npu_inst_pe_1_7_4_N72,
         npu_inst_pe_1_7_4_N71, npu_inst_pe_1_7_4_N70, npu_inst_pe_1_7_4_N69,
         npu_inst_pe_1_7_4_N68, npu_inst_pe_1_7_4_N67, npu_inst_pe_1_7_4_N66,
         npu_inst_pe_1_7_4_N65, npu_inst_pe_1_7_4_int_data_0_,
         npu_inst_pe_1_7_4_int_data_1_, npu_inst_pe_1_7_4_int_q_weight_0_,
         npu_inst_pe_1_7_4_int_q_weight_1_,
         npu_inst_pe_1_7_4_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_4_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_4_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_4_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_4_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_4_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_4_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_4_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_4_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_4_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_4_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_4_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_4_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_4_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_4_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_4_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_4_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_4_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_4_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_4_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_4_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_4_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_4_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_4_int_q_reg_h_0__1_, npu_inst_pe_1_7_5_n118,
         npu_inst_pe_1_7_5_n117, npu_inst_pe_1_7_5_n116,
         npu_inst_pe_1_7_5_n115, npu_inst_pe_1_7_5_n114,
         npu_inst_pe_1_7_5_n113, npu_inst_pe_1_7_5_n112,
         npu_inst_pe_1_7_5_n111, npu_inst_pe_1_7_5_n110,
         npu_inst_pe_1_7_5_n109, npu_inst_pe_1_7_5_n108,
         npu_inst_pe_1_7_5_n107, npu_inst_pe_1_7_5_n106,
         npu_inst_pe_1_7_5_n105, npu_inst_pe_1_7_5_n104,
         npu_inst_pe_1_7_5_n103, npu_inst_pe_1_7_5_n102,
         npu_inst_pe_1_7_5_n101, npu_inst_pe_1_7_5_n100, npu_inst_pe_1_7_5_n99,
         npu_inst_pe_1_7_5_n98, npu_inst_pe_1_7_5_n36, npu_inst_pe_1_7_5_n35,
         npu_inst_pe_1_7_5_n34, npu_inst_pe_1_7_5_n33, npu_inst_pe_1_7_5_n32,
         npu_inst_pe_1_7_5_n31, npu_inst_pe_1_7_5_n30, npu_inst_pe_1_7_5_n29,
         npu_inst_pe_1_7_5_n28, npu_inst_pe_1_7_5_n25, npu_inst_pe_1_7_5_n24,
         npu_inst_pe_1_7_5_n23, npu_inst_pe_1_7_5_n22, npu_inst_pe_1_7_5_n21,
         npu_inst_pe_1_7_5_n20, npu_inst_pe_1_7_5_n19, npu_inst_pe_1_7_5_n18,
         npu_inst_pe_1_7_5_n17, npu_inst_pe_1_7_5_n16, npu_inst_pe_1_7_5_n15,
         npu_inst_pe_1_7_5_n14, npu_inst_pe_1_7_5_n13, npu_inst_pe_1_7_5_n12,
         npu_inst_pe_1_7_5_n11, npu_inst_pe_1_7_5_n10, npu_inst_pe_1_7_5_n9,
         npu_inst_pe_1_7_5_n8, npu_inst_pe_1_7_5_n7, npu_inst_pe_1_7_5_n6,
         npu_inst_pe_1_7_5_n5, npu_inst_pe_1_7_5_n4, npu_inst_pe_1_7_5_n3,
         npu_inst_pe_1_7_5_n2, npu_inst_pe_1_7_5_n1,
         npu_inst_pe_1_7_5_sub_77_carry_7_, npu_inst_pe_1_7_5_sub_77_carry_6_,
         npu_inst_pe_1_7_5_sub_77_carry_5_, npu_inst_pe_1_7_5_sub_77_carry_4_,
         npu_inst_pe_1_7_5_sub_77_carry_3_, npu_inst_pe_1_7_5_sub_77_carry_2_,
         npu_inst_pe_1_7_5_sub_77_carry_1_, npu_inst_pe_1_7_5_add_79_carry_7_,
         npu_inst_pe_1_7_5_add_79_carry_6_, npu_inst_pe_1_7_5_add_79_carry_5_,
         npu_inst_pe_1_7_5_add_79_carry_4_, npu_inst_pe_1_7_5_add_79_carry_3_,
         npu_inst_pe_1_7_5_add_79_carry_2_, npu_inst_pe_1_7_5_add_79_carry_1_,
         npu_inst_pe_1_7_5_n97, npu_inst_pe_1_7_5_n96, npu_inst_pe_1_7_5_n95,
         npu_inst_pe_1_7_5_n94, npu_inst_pe_1_7_5_n93, npu_inst_pe_1_7_5_n92,
         npu_inst_pe_1_7_5_n91, npu_inst_pe_1_7_5_n90, npu_inst_pe_1_7_5_n89,
         npu_inst_pe_1_7_5_n88, npu_inst_pe_1_7_5_n87, npu_inst_pe_1_7_5_n86,
         npu_inst_pe_1_7_5_n85, npu_inst_pe_1_7_5_n84, npu_inst_pe_1_7_5_n83,
         npu_inst_pe_1_7_5_n82, npu_inst_pe_1_7_5_n81, npu_inst_pe_1_7_5_n80,
         npu_inst_pe_1_7_5_n79, npu_inst_pe_1_7_5_n78, npu_inst_pe_1_7_5_n77,
         npu_inst_pe_1_7_5_n76, npu_inst_pe_1_7_5_n75, npu_inst_pe_1_7_5_n74,
         npu_inst_pe_1_7_5_n73, npu_inst_pe_1_7_5_n72, npu_inst_pe_1_7_5_n71,
         npu_inst_pe_1_7_5_n70, npu_inst_pe_1_7_5_n69, npu_inst_pe_1_7_5_n68,
         npu_inst_pe_1_7_5_n67, npu_inst_pe_1_7_5_n66, npu_inst_pe_1_7_5_n65,
         npu_inst_pe_1_7_5_n64, npu_inst_pe_1_7_5_n63, npu_inst_pe_1_7_5_n62,
         npu_inst_pe_1_7_5_n61, npu_inst_pe_1_7_5_n60, npu_inst_pe_1_7_5_n59,
         npu_inst_pe_1_7_5_n58, npu_inst_pe_1_7_5_n57, npu_inst_pe_1_7_5_n56,
         npu_inst_pe_1_7_5_n55, npu_inst_pe_1_7_5_n54, npu_inst_pe_1_7_5_n53,
         npu_inst_pe_1_7_5_n52, npu_inst_pe_1_7_5_n51, npu_inst_pe_1_7_5_n50,
         npu_inst_pe_1_7_5_n49, npu_inst_pe_1_7_5_n48, npu_inst_pe_1_7_5_n47,
         npu_inst_pe_1_7_5_n46, npu_inst_pe_1_7_5_n45, npu_inst_pe_1_7_5_n44,
         npu_inst_pe_1_7_5_n43, npu_inst_pe_1_7_5_n42, npu_inst_pe_1_7_5_n41,
         npu_inst_pe_1_7_5_n40, npu_inst_pe_1_7_5_n39, npu_inst_pe_1_7_5_n38,
         npu_inst_pe_1_7_5_n37, npu_inst_pe_1_7_5_n27, npu_inst_pe_1_7_5_n26,
         npu_inst_pe_1_7_5_net3081, npu_inst_pe_1_7_5_net3075,
         npu_inst_pe_1_7_5_N94, npu_inst_pe_1_7_5_N93, npu_inst_pe_1_7_5_N84,
         npu_inst_pe_1_7_5_N80, npu_inst_pe_1_7_5_N79, npu_inst_pe_1_7_5_N78,
         npu_inst_pe_1_7_5_N77, npu_inst_pe_1_7_5_N76, npu_inst_pe_1_7_5_N75,
         npu_inst_pe_1_7_5_N74, npu_inst_pe_1_7_5_N73, npu_inst_pe_1_7_5_N72,
         npu_inst_pe_1_7_5_N71, npu_inst_pe_1_7_5_N70, npu_inst_pe_1_7_5_N69,
         npu_inst_pe_1_7_5_N68, npu_inst_pe_1_7_5_N67, npu_inst_pe_1_7_5_N66,
         npu_inst_pe_1_7_5_N65, npu_inst_pe_1_7_5_int_data_0_,
         npu_inst_pe_1_7_5_int_data_1_, npu_inst_pe_1_7_5_int_q_weight_0_,
         npu_inst_pe_1_7_5_int_q_weight_1_,
         npu_inst_pe_1_7_5_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_5_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_5_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_5_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_5_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_5_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_5_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_5_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_5_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_5_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_5_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_5_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_5_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_5_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_5_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_5_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_5_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_5_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_5_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_5_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_5_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_5_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_5_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_5_int_q_reg_h_0__1_, npu_inst_pe_1_7_6_n118,
         npu_inst_pe_1_7_6_n117, npu_inst_pe_1_7_6_n116,
         npu_inst_pe_1_7_6_n115, npu_inst_pe_1_7_6_n114,
         npu_inst_pe_1_7_6_n113, npu_inst_pe_1_7_6_n112,
         npu_inst_pe_1_7_6_n111, npu_inst_pe_1_7_6_n110,
         npu_inst_pe_1_7_6_n109, npu_inst_pe_1_7_6_n108,
         npu_inst_pe_1_7_6_n107, npu_inst_pe_1_7_6_n106,
         npu_inst_pe_1_7_6_n105, npu_inst_pe_1_7_6_n104,
         npu_inst_pe_1_7_6_n103, npu_inst_pe_1_7_6_n102,
         npu_inst_pe_1_7_6_n101, npu_inst_pe_1_7_6_n100, npu_inst_pe_1_7_6_n99,
         npu_inst_pe_1_7_6_n98, npu_inst_pe_1_7_6_n36, npu_inst_pe_1_7_6_n35,
         npu_inst_pe_1_7_6_n34, npu_inst_pe_1_7_6_n33, npu_inst_pe_1_7_6_n32,
         npu_inst_pe_1_7_6_n31, npu_inst_pe_1_7_6_n30, npu_inst_pe_1_7_6_n29,
         npu_inst_pe_1_7_6_n28, npu_inst_pe_1_7_6_n25, npu_inst_pe_1_7_6_n24,
         npu_inst_pe_1_7_6_n23, npu_inst_pe_1_7_6_n22, npu_inst_pe_1_7_6_n21,
         npu_inst_pe_1_7_6_n20, npu_inst_pe_1_7_6_n19, npu_inst_pe_1_7_6_n18,
         npu_inst_pe_1_7_6_n17, npu_inst_pe_1_7_6_n16, npu_inst_pe_1_7_6_n15,
         npu_inst_pe_1_7_6_n14, npu_inst_pe_1_7_6_n13, npu_inst_pe_1_7_6_n12,
         npu_inst_pe_1_7_6_n11, npu_inst_pe_1_7_6_n10, npu_inst_pe_1_7_6_n9,
         npu_inst_pe_1_7_6_n8, npu_inst_pe_1_7_6_n7, npu_inst_pe_1_7_6_n6,
         npu_inst_pe_1_7_6_n5, npu_inst_pe_1_7_6_n4, npu_inst_pe_1_7_6_n3,
         npu_inst_pe_1_7_6_n2, npu_inst_pe_1_7_6_n1,
         npu_inst_pe_1_7_6_sub_77_carry_7_, npu_inst_pe_1_7_6_sub_77_carry_6_,
         npu_inst_pe_1_7_6_sub_77_carry_5_, npu_inst_pe_1_7_6_sub_77_carry_4_,
         npu_inst_pe_1_7_6_sub_77_carry_3_, npu_inst_pe_1_7_6_sub_77_carry_2_,
         npu_inst_pe_1_7_6_sub_77_carry_1_, npu_inst_pe_1_7_6_add_79_carry_7_,
         npu_inst_pe_1_7_6_add_79_carry_6_, npu_inst_pe_1_7_6_add_79_carry_5_,
         npu_inst_pe_1_7_6_add_79_carry_4_, npu_inst_pe_1_7_6_add_79_carry_3_,
         npu_inst_pe_1_7_6_add_79_carry_2_, npu_inst_pe_1_7_6_add_79_carry_1_,
         npu_inst_pe_1_7_6_n97, npu_inst_pe_1_7_6_n96, npu_inst_pe_1_7_6_n95,
         npu_inst_pe_1_7_6_n94, npu_inst_pe_1_7_6_n93, npu_inst_pe_1_7_6_n92,
         npu_inst_pe_1_7_6_n91, npu_inst_pe_1_7_6_n90, npu_inst_pe_1_7_6_n89,
         npu_inst_pe_1_7_6_n88, npu_inst_pe_1_7_6_n87, npu_inst_pe_1_7_6_n86,
         npu_inst_pe_1_7_6_n85, npu_inst_pe_1_7_6_n84, npu_inst_pe_1_7_6_n83,
         npu_inst_pe_1_7_6_n82, npu_inst_pe_1_7_6_n81, npu_inst_pe_1_7_6_n80,
         npu_inst_pe_1_7_6_n79, npu_inst_pe_1_7_6_n78, npu_inst_pe_1_7_6_n77,
         npu_inst_pe_1_7_6_n76, npu_inst_pe_1_7_6_n75, npu_inst_pe_1_7_6_n74,
         npu_inst_pe_1_7_6_n73, npu_inst_pe_1_7_6_n72, npu_inst_pe_1_7_6_n71,
         npu_inst_pe_1_7_6_n70, npu_inst_pe_1_7_6_n69, npu_inst_pe_1_7_6_n68,
         npu_inst_pe_1_7_6_n67, npu_inst_pe_1_7_6_n66, npu_inst_pe_1_7_6_n65,
         npu_inst_pe_1_7_6_n64, npu_inst_pe_1_7_6_n63, npu_inst_pe_1_7_6_n62,
         npu_inst_pe_1_7_6_n61, npu_inst_pe_1_7_6_n60, npu_inst_pe_1_7_6_n59,
         npu_inst_pe_1_7_6_n58, npu_inst_pe_1_7_6_n57, npu_inst_pe_1_7_6_n56,
         npu_inst_pe_1_7_6_n55, npu_inst_pe_1_7_6_n54, npu_inst_pe_1_7_6_n53,
         npu_inst_pe_1_7_6_n52, npu_inst_pe_1_7_6_n51, npu_inst_pe_1_7_6_n50,
         npu_inst_pe_1_7_6_n49, npu_inst_pe_1_7_6_n48, npu_inst_pe_1_7_6_n47,
         npu_inst_pe_1_7_6_n46, npu_inst_pe_1_7_6_n45, npu_inst_pe_1_7_6_n44,
         npu_inst_pe_1_7_6_n43, npu_inst_pe_1_7_6_n42, npu_inst_pe_1_7_6_n41,
         npu_inst_pe_1_7_6_n40, npu_inst_pe_1_7_6_n39, npu_inst_pe_1_7_6_n38,
         npu_inst_pe_1_7_6_n37, npu_inst_pe_1_7_6_n27, npu_inst_pe_1_7_6_n26,
         npu_inst_pe_1_7_6_net3058, npu_inst_pe_1_7_6_net3052,
         npu_inst_pe_1_7_6_N94, npu_inst_pe_1_7_6_N93, npu_inst_pe_1_7_6_N84,
         npu_inst_pe_1_7_6_N80, npu_inst_pe_1_7_6_N79, npu_inst_pe_1_7_6_N78,
         npu_inst_pe_1_7_6_N77, npu_inst_pe_1_7_6_N76, npu_inst_pe_1_7_6_N75,
         npu_inst_pe_1_7_6_N74, npu_inst_pe_1_7_6_N73, npu_inst_pe_1_7_6_N72,
         npu_inst_pe_1_7_6_N71, npu_inst_pe_1_7_6_N70, npu_inst_pe_1_7_6_N69,
         npu_inst_pe_1_7_6_N68, npu_inst_pe_1_7_6_N67, npu_inst_pe_1_7_6_N66,
         npu_inst_pe_1_7_6_N65, npu_inst_pe_1_7_6_int_data_0_,
         npu_inst_pe_1_7_6_int_data_1_, npu_inst_pe_1_7_6_int_q_weight_0_,
         npu_inst_pe_1_7_6_int_q_weight_1_,
         npu_inst_pe_1_7_6_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_6_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_6_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_6_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_6_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_6_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_6_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_6_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_6_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_6_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_6_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_6_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_6_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_6_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_6_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_6_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_6_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_6_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_6_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_6_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_6_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_6_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_6_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_6_int_q_reg_h_0__1_, npu_inst_pe_1_7_7_n118,
         npu_inst_pe_1_7_7_n117, npu_inst_pe_1_7_7_n116,
         npu_inst_pe_1_7_7_n115, npu_inst_pe_1_7_7_n114,
         npu_inst_pe_1_7_7_n113, npu_inst_pe_1_7_7_n112,
         npu_inst_pe_1_7_7_n111, npu_inst_pe_1_7_7_n110,
         npu_inst_pe_1_7_7_n109, npu_inst_pe_1_7_7_n108,
         npu_inst_pe_1_7_7_n107, npu_inst_pe_1_7_7_n106,
         npu_inst_pe_1_7_7_n105, npu_inst_pe_1_7_7_n104,
         npu_inst_pe_1_7_7_n103, npu_inst_pe_1_7_7_n102,
         npu_inst_pe_1_7_7_n101, npu_inst_pe_1_7_7_n100, npu_inst_pe_1_7_7_n99,
         npu_inst_pe_1_7_7_n98, npu_inst_pe_1_7_7_n36, npu_inst_pe_1_7_7_n35,
         npu_inst_pe_1_7_7_n34, npu_inst_pe_1_7_7_n33, npu_inst_pe_1_7_7_n32,
         npu_inst_pe_1_7_7_n31, npu_inst_pe_1_7_7_n30, npu_inst_pe_1_7_7_n29,
         npu_inst_pe_1_7_7_n28, npu_inst_pe_1_7_7_n25, npu_inst_pe_1_7_7_n24,
         npu_inst_pe_1_7_7_n23, npu_inst_pe_1_7_7_n22, npu_inst_pe_1_7_7_n21,
         npu_inst_pe_1_7_7_n20, npu_inst_pe_1_7_7_n19, npu_inst_pe_1_7_7_n18,
         npu_inst_pe_1_7_7_n17, npu_inst_pe_1_7_7_n16, npu_inst_pe_1_7_7_n15,
         npu_inst_pe_1_7_7_n14, npu_inst_pe_1_7_7_n13, npu_inst_pe_1_7_7_n12,
         npu_inst_pe_1_7_7_n11, npu_inst_pe_1_7_7_n10, npu_inst_pe_1_7_7_n9,
         npu_inst_pe_1_7_7_n8, npu_inst_pe_1_7_7_n7, npu_inst_pe_1_7_7_n6,
         npu_inst_pe_1_7_7_n5, npu_inst_pe_1_7_7_n4, npu_inst_pe_1_7_7_n3,
         npu_inst_pe_1_7_7_n2, npu_inst_pe_1_7_7_n1,
         npu_inst_pe_1_7_7_sub_77_carry_7_, npu_inst_pe_1_7_7_sub_77_carry_6_,
         npu_inst_pe_1_7_7_sub_77_carry_5_, npu_inst_pe_1_7_7_sub_77_carry_4_,
         npu_inst_pe_1_7_7_sub_77_carry_3_, npu_inst_pe_1_7_7_sub_77_carry_2_,
         npu_inst_pe_1_7_7_sub_77_carry_1_, npu_inst_pe_1_7_7_add_79_carry_7_,
         npu_inst_pe_1_7_7_add_79_carry_6_, npu_inst_pe_1_7_7_add_79_carry_5_,
         npu_inst_pe_1_7_7_add_79_carry_4_, npu_inst_pe_1_7_7_add_79_carry_3_,
         npu_inst_pe_1_7_7_add_79_carry_2_, npu_inst_pe_1_7_7_add_79_carry_1_,
         npu_inst_pe_1_7_7_n97, npu_inst_pe_1_7_7_n96, npu_inst_pe_1_7_7_n95,
         npu_inst_pe_1_7_7_n94, npu_inst_pe_1_7_7_n93, npu_inst_pe_1_7_7_n92,
         npu_inst_pe_1_7_7_n91, npu_inst_pe_1_7_7_n90, npu_inst_pe_1_7_7_n89,
         npu_inst_pe_1_7_7_n88, npu_inst_pe_1_7_7_n87, npu_inst_pe_1_7_7_n86,
         npu_inst_pe_1_7_7_n85, npu_inst_pe_1_7_7_n84, npu_inst_pe_1_7_7_n83,
         npu_inst_pe_1_7_7_n82, npu_inst_pe_1_7_7_n81, npu_inst_pe_1_7_7_n80,
         npu_inst_pe_1_7_7_n79, npu_inst_pe_1_7_7_n78, npu_inst_pe_1_7_7_n77,
         npu_inst_pe_1_7_7_n76, npu_inst_pe_1_7_7_n75, npu_inst_pe_1_7_7_n74,
         npu_inst_pe_1_7_7_n73, npu_inst_pe_1_7_7_n72, npu_inst_pe_1_7_7_n71,
         npu_inst_pe_1_7_7_n70, npu_inst_pe_1_7_7_n69, npu_inst_pe_1_7_7_n68,
         npu_inst_pe_1_7_7_n67, npu_inst_pe_1_7_7_n66, npu_inst_pe_1_7_7_n65,
         npu_inst_pe_1_7_7_n64, npu_inst_pe_1_7_7_n63, npu_inst_pe_1_7_7_n62,
         npu_inst_pe_1_7_7_n61, npu_inst_pe_1_7_7_n60, npu_inst_pe_1_7_7_n59,
         npu_inst_pe_1_7_7_n58, npu_inst_pe_1_7_7_n57, npu_inst_pe_1_7_7_n56,
         npu_inst_pe_1_7_7_n55, npu_inst_pe_1_7_7_n54, npu_inst_pe_1_7_7_n53,
         npu_inst_pe_1_7_7_n52, npu_inst_pe_1_7_7_n51, npu_inst_pe_1_7_7_n50,
         npu_inst_pe_1_7_7_n49, npu_inst_pe_1_7_7_n48, npu_inst_pe_1_7_7_n47,
         npu_inst_pe_1_7_7_n46, npu_inst_pe_1_7_7_n45, npu_inst_pe_1_7_7_n44,
         npu_inst_pe_1_7_7_n43, npu_inst_pe_1_7_7_n42, npu_inst_pe_1_7_7_n41,
         npu_inst_pe_1_7_7_n40, npu_inst_pe_1_7_7_n39, npu_inst_pe_1_7_7_n38,
         npu_inst_pe_1_7_7_n37, npu_inst_pe_1_7_7_n27, npu_inst_pe_1_7_7_n26,
         npu_inst_pe_1_7_7_net3035, npu_inst_pe_1_7_7_net3029,
         npu_inst_pe_1_7_7_N94, npu_inst_pe_1_7_7_N93, npu_inst_pe_1_7_7_N84,
         npu_inst_pe_1_7_7_N80, npu_inst_pe_1_7_7_N79, npu_inst_pe_1_7_7_N78,
         npu_inst_pe_1_7_7_N77, npu_inst_pe_1_7_7_N76, npu_inst_pe_1_7_7_N75,
         npu_inst_pe_1_7_7_N74, npu_inst_pe_1_7_7_N73, npu_inst_pe_1_7_7_N72,
         npu_inst_pe_1_7_7_N71, npu_inst_pe_1_7_7_N70, npu_inst_pe_1_7_7_N69,
         npu_inst_pe_1_7_7_N68, npu_inst_pe_1_7_7_N67, npu_inst_pe_1_7_7_N66,
         npu_inst_pe_1_7_7_N65, npu_inst_pe_1_7_7_int_data_0_,
         npu_inst_pe_1_7_7_int_data_1_, npu_inst_pe_1_7_7_int_q_weight_0_,
         npu_inst_pe_1_7_7_int_q_weight_1_,
         npu_inst_pe_1_7_7_int_q_reg_v_5__0_,
         npu_inst_pe_1_7_7_int_q_reg_v_5__1_,
         npu_inst_pe_1_7_7_int_q_reg_v_4__0_,
         npu_inst_pe_1_7_7_int_q_reg_v_4__1_,
         npu_inst_pe_1_7_7_int_q_reg_v_3__0_,
         npu_inst_pe_1_7_7_int_q_reg_v_3__1_,
         npu_inst_pe_1_7_7_int_q_reg_v_2__0_,
         npu_inst_pe_1_7_7_int_q_reg_v_2__1_,
         npu_inst_pe_1_7_7_int_q_reg_v_1__0_,
         npu_inst_pe_1_7_7_int_q_reg_v_1__1_,
         npu_inst_pe_1_7_7_int_q_reg_v_0__0_,
         npu_inst_pe_1_7_7_int_q_reg_v_0__1_,
         npu_inst_pe_1_7_7_int_q_reg_h_5__0_,
         npu_inst_pe_1_7_7_int_q_reg_h_5__1_,
         npu_inst_pe_1_7_7_int_q_reg_h_4__0_,
         npu_inst_pe_1_7_7_int_q_reg_h_4__1_,
         npu_inst_pe_1_7_7_int_q_reg_h_3__0_,
         npu_inst_pe_1_7_7_int_q_reg_h_3__1_,
         npu_inst_pe_1_7_7_int_q_reg_h_2__0_,
         npu_inst_pe_1_7_7_int_q_reg_h_2__1_,
         npu_inst_pe_1_7_7_int_q_reg_h_1__0_,
         npu_inst_pe_1_7_7_int_q_reg_h_1__1_,
         npu_inst_pe_1_7_7_int_q_reg_h_0__0_,
         npu_inst_pe_1_7_7_int_q_reg_h_0__1_, qrelu_i_0_n3, qrelu_i_0_n2,
         qrelu_i_0_n1, qrelu_i_0_n6, qrelu_i_0_n5, qrelu_i_0_n4, qrelu_i_1_n9,
         qrelu_i_1_n8, qrelu_i_1_n7, qrelu_i_1_n3, qrelu_i_1_n2, qrelu_i_1_n1,
         qrelu_i_2_n9, qrelu_i_2_n8, qrelu_i_2_n7, qrelu_i_2_n3, qrelu_i_2_n2,
         qrelu_i_2_n1, qrelu_i_3_n9, qrelu_i_3_n8, qrelu_i_3_n7, qrelu_i_3_n3,
         qrelu_i_3_n2, qrelu_i_3_n1, qrelu_i_4_n9, qrelu_i_4_n8, qrelu_i_4_n7,
         qrelu_i_4_n3, qrelu_i_4_n2, qrelu_i_4_n1, qrelu_i_5_n9, qrelu_i_5_n8,
         qrelu_i_5_n7, qrelu_i_5_n3, qrelu_i_5_n2, qrelu_i_5_n1, qrelu_i_6_n9,
         qrelu_i_6_n8, qrelu_i_6_n7, qrelu_i_6_n3, qrelu_i_6_n2, qrelu_i_6_n1,
         qrelu_i_7_n9, qrelu_i_7_n8, qrelu_i_7_n7, qrelu_i_7_n3, qrelu_i_7_n2,
         qrelu_i_7_n1, p_unit_i_0_n17, p_unit_i_0_n16, p_unit_i_0_n12,
         p_unit_i_0_n11, p_unit_i_0_n7, p_unit_i_0_n6, p_unit_i_0_n5,
         p_unit_i_0_n4, p_unit_i_0_n3, p_unit_i_0_n2, p_unit_i_0_n1,
         p_unit_i_0_n15, p_unit_i_0_n14, p_unit_i_0_n13, p_unit_i_0_n10,
         p_unit_i_0_n9, p_unit_i_0_n8, p_unit_i_0_net3011, p_unit_i_0_N7,
         p_unit_i_0_N6, p_unit_i_0_N5, p_unit_i_0_N3, p_unit_i_0_N2,
         p_unit_i_0_int_ps1_0_, p_unit_i_0_int_ps1_1_, p_unit_i_0_int_ps1_2_,
         p_unit_i_0_int_ps0_0_, p_unit_i_0_int_ps0_1_, p_unit_i_0_int_ps0_2_,
         p_unit_i_1_n17, p_unit_i_1_n16, p_unit_i_1_n12, p_unit_i_1_n11,
         p_unit_i_1_n7, p_unit_i_1_n6, p_unit_i_1_n5, p_unit_i_1_n4,
         p_unit_i_1_n3, p_unit_i_1_n2, p_unit_i_1_n1, p_unit_i_1_n15,
         p_unit_i_1_n14, p_unit_i_1_n13, p_unit_i_1_n10, p_unit_i_1_n9,
         p_unit_i_1_n8, p_unit_i_1_net2993, p_unit_i_1_N7, p_unit_i_1_N6,
         p_unit_i_1_N5, p_unit_i_1_N3, p_unit_i_1_N2, p_unit_i_1_int_ps1_0_,
         p_unit_i_1_int_ps1_1_, p_unit_i_1_int_ps1_2_, p_unit_i_1_int_ps0_0_,
         p_unit_i_1_int_ps0_1_, p_unit_i_1_int_ps0_2_, p_unit_i_2_n17,
         p_unit_i_2_n16, p_unit_i_2_n12, p_unit_i_2_n11, p_unit_i_2_n7,
         p_unit_i_2_n6, p_unit_i_2_n5, p_unit_i_2_n4, p_unit_i_2_n3,
         p_unit_i_2_n2, p_unit_i_2_n1, p_unit_i_2_n15, p_unit_i_2_n14,
         p_unit_i_2_n13, p_unit_i_2_n10, p_unit_i_2_n9, p_unit_i_2_n8,
         p_unit_i_2_net2975, p_unit_i_2_N7, p_unit_i_2_N6, p_unit_i_2_N5,
         p_unit_i_2_N3, p_unit_i_2_N2, p_unit_i_2_int_ps1_0_,
         p_unit_i_2_int_ps1_1_, p_unit_i_2_int_ps1_2_, p_unit_i_2_int_ps0_0_,
         p_unit_i_2_int_ps0_1_, p_unit_i_2_int_ps0_2_, p_unit_i_3_n17,
         p_unit_i_3_n16, p_unit_i_3_n12, p_unit_i_3_n11, p_unit_i_3_n7,
         p_unit_i_3_n6, p_unit_i_3_n5, p_unit_i_3_n4, p_unit_i_3_n3,
         p_unit_i_3_n2, p_unit_i_3_n1, p_unit_i_3_n15, p_unit_i_3_n14,
         p_unit_i_3_n13, p_unit_i_3_n10, p_unit_i_3_n9, p_unit_i_3_n8,
         p_unit_i_3_net2957, p_unit_i_3_N7, p_unit_i_3_N6, p_unit_i_3_N5,
         p_unit_i_3_N3, p_unit_i_3_N2, p_unit_i_3_int_ps1_0_,
         p_unit_i_3_int_ps1_1_, p_unit_i_3_int_ps1_2_, p_unit_i_3_int_ps0_0_,
         p_unit_i_3_int_ps0_1_, p_unit_i_3_int_ps0_2_, round_i_0_n2,
         round_i_0_n1, round_i_0_n3, round_i_1_n4, round_i_1_n2, round_i_1_n1,
         round_i_2_n4, round_i_2_n2, round_i_2_n1, round_i_3_n4, round_i_3_n2,
         round_i_3_n1, hmode_cnt_inst_n12, hmode_cnt_inst_n6,
         hmode_cnt_inst_n4, hmode_cnt_inst_n2, hmode_cnt_inst_n1,
         hmode_cnt_inst_n11, hmode_cnt_inst_n10, hmode_cnt_inst_n9,
         hmode_cnt_inst_n8, hmode_cnt_inst_n7, hmode_cnt_inst_n5,
         hmode_cnt_inst_net2939, hmode_cnt_inst_N12, hmode_cnt_inst_N10,
         vmode_cnt_inst_n12, vmode_cnt_inst_n6, vmode_cnt_inst_n4,
         vmode_cnt_inst_n2, vmode_cnt_inst_n1, vmode_cnt_inst_n11,
         vmode_cnt_inst_n10, vmode_cnt_inst_n9, vmode_cnt_inst_n8,
         vmode_cnt_inst_n7, vmode_cnt_inst_n5, vmode_cnt_inst_net2921,
         vmode_cnt_inst_N12, vmode_cnt_inst_N10, vmode_cnt_inst_q_0_,
         vmode_cnt_inst_q_1_, vmode_cnt_inst_q_2_, res_cnt_inst_n2,
         res_cnt_inst_n1, res_cnt_inst_n14, res_cnt_inst_n13, res_cnt_inst_n12,
         res_cnt_inst_n11, res_cnt_inst_n10, res_cnt_inst_n9, res_cnt_inst_n8,
         res_cnt_inst_n7, res_cnt_inst_n5, res_cnt_inst_net2903,
         res_cnt_inst_N12, res_cnt_inst_N10, res_cnt_inst_q_0_,
         res_cnt_inst_q_1_, res_cnt_inst_q_2_, i_data_npu_cnt_inst_n12,
         i_data_npu_cnt_inst_n6, i_data_npu_cnt_inst_n4,
         i_data_npu_cnt_inst_n2, i_data_npu_cnt_inst_n1,
         i_data_npu_cnt_inst_n11, i_data_npu_cnt_inst_n10,
         i_data_npu_cnt_inst_n9, i_data_npu_cnt_inst_n8,
         i_data_npu_cnt_inst_n7, i_data_npu_cnt_inst_n5,
         i_data_npu_cnt_inst_net2885, i_data_npu_cnt_inst_N12,
         i_data_npu_cnt_inst_N10, i_data_tilev_cnt_inst_n8,
         i_data_tilev_cnt_inst_n6, i_data_tilev_cnt_inst_n3,
         i_data_tilev_cnt_inst_n2, i_data_tilev_cnt_inst_n1,
         i_data_tilev_cnt_inst_n17, i_data_tilev_cnt_inst_n15,
         i_data_tilev_cnt_inst_n14, i_data_tilev_cnt_inst_n13,
         i_data_tilev_cnt_inst_n12, i_data_tilev_cnt_inst_n11,
         i_data_tilev_cnt_inst_n9, i_data_tilev_cnt_inst_n7,
         i_data_tilev_cnt_inst_n5, i_data_tilev_cnt_inst_n4,
         i_data_tilev_cnt_inst_q_0_, i_data_tilev_cnt_inst_q_1_,
         i_data_tileh_cnt_inst_n24, i_data_tileh_cnt_inst_n23,
         i_data_tileh_cnt_inst_n22, i_data_tileh_cnt_inst_n21,
         i_data_tileh_cnt_inst_n20, i_data_tileh_cnt_inst_n19,
         i_data_tileh_cnt_inst_n18, i_data_tileh_cnt_inst_n17,
         i_data_tileh_cnt_inst_n16, i_data_tileh_cnt_inst_n10,
         i_data_tileh_cnt_inst_n8, i_data_tileh_cnt_inst_n6,
         i_data_tileh_cnt_inst_n3, i_data_tileh_cnt_inst_n2,
         i_data_tileh_cnt_inst_n1, ifmaps_cnt_inst_n12, ifmaps_cnt_inst_n6,
         ifmaps_cnt_inst_n4, ifmaps_cnt_inst_n2, ifmaps_cnt_inst_n1,
         ifmaps_cnt_inst_n11, ifmaps_cnt_inst_n10, ifmaps_cnt_inst_n9,
         ifmaps_cnt_inst_n8, ifmaps_cnt_inst_n7, ifmaps_cnt_inst_n5,
         ifmaps_cnt_inst_net2867, ifmaps_cnt_inst_N12, ifmaps_cnt_inst_N10,
         ofmaps_cnt_inst_n4, ofmaps_cnt_inst_n2, ofmaps_cnt_inst_n1,
         ofmaps_cnt_inst_n19, ofmaps_cnt_inst_n18, ofmaps_cnt_inst_n17,
         ofmaps_cnt_inst_n16, ofmaps_cnt_inst_n15, ofmaps_cnt_inst_n14,
         ofmaps_cnt_inst_n13, ofmaps_cnt_inst_n12, ofmaps_cnt_inst_n11,
         ofmaps_cnt_inst_n10, ofmaps_cnt_inst_n9, ofmaps_cnt_inst_n8,
         ofmaps_cnt_inst_n5, ofmaps_cnt_inst_net2849, ofmaps_cnt_inst_N14,
         ofmaps_cnt_inst_N13, ofmaps_cnt_inst_N11, ofmaps_cnt_inst_q_0_,
         ofmaps_cnt_inst_q_1_, ofmaps_cnt_inst_q_2_, ofmaps_cnt_inst_q_3_,
         i_weight_addr_gen_inst_n64, i_weight_addr_gen_inst_n63,
         i_weight_addr_gen_inst_n62, i_weight_addr_gen_inst_n43,
         i_weight_addr_gen_inst_n42, i_weight_addr_gen_inst_n41,
         i_weight_addr_gen_inst_n40, i_weight_addr_gen_inst_n39,
         i_weight_addr_gen_inst_n38, i_weight_addr_gen_inst_n37,
         i_weight_addr_gen_inst_n36, i_weight_addr_gen_inst_n35,
         i_weight_addr_gen_inst_n34, i_weight_addr_gen_inst_n33,
         i_weight_addr_gen_inst_n32, i_weight_addr_gen_inst_n31,
         i_weight_addr_gen_inst_n30, i_weight_addr_gen_inst_n29,
         i_weight_addr_gen_inst_n28, i_weight_addr_gen_inst_n27,
         i_weight_addr_gen_inst_n26, i_weight_addr_gen_inst_n24,
         i_weight_addr_gen_inst_n8, i_weight_addr_gen_inst_n7,
         i_weight_addr_gen_inst_n6, i_weight_addr_gen_inst_n5,
         i_weight_addr_gen_inst_n61, i_weight_addr_gen_inst_n60,
         i_weight_addr_gen_inst_n59, i_weight_addr_gen_inst_n58,
         i_weight_addr_gen_inst_n57, i_weight_addr_gen_inst_n56,
         i_weight_addr_gen_inst_n55, i_weight_addr_gen_inst_n54,
         i_weight_addr_gen_inst_n53, i_weight_addr_gen_inst_n52,
         i_weight_addr_gen_inst_n51, i_weight_addr_gen_inst_n50,
         i_weight_addr_gen_inst_n49, i_weight_addr_gen_inst_n48,
         i_weight_addr_gen_inst_n47, i_weight_addr_gen_inst_n46,
         i_weight_addr_gen_inst_n45, i_weight_addr_gen_inst_n44,
         i_weight_addr_gen_inst_net2832, i_weight_addr_gen_inst_net2826,
         i_weight_addr_gen_inst_N95, i_weight_addr_gen_inst_N94,
         i_weight_addr_gen_inst_N93, i_weight_addr_gen_inst_N92,
         i_weight_addr_gen_inst_N91, i_weight_addr_gen_inst_N90,
         i_weight_addr_gen_inst_N89, i_weight_addr_gen_inst_N88,
         i_weight_addr_gen_inst_N87, i_weight_addr_gen_inst_N86,
         i_weight_addr_gen_inst_N85, i_weight_addr_gen_inst_N84,
         i_weight_addr_gen_inst_N83, i_weight_addr_gen_inst_N82,
         i_weight_addr_gen_inst_N81, i_weight_addr_gen_inst_N80,
         i_weight_addr_gen_inst_N79, i_weight_addr_gen_inst_N58,
         i_weight_addr_gen_inst_N41, i_weight_addr_gen_inst_N40,
         i_weight_addr_gen_inst_N39, i_weight_addr_gen_inst_N38,
         i_weight_addr_gen_inst_N37, i_weight_addr_gen_inst_N36,
         i_weight_addr_gen_inst_N35, i_weight_addr_gen_inst_N34,
         i_weight_addr_gen_inst_N33, i_weight_addr_gen_inst_N32,
         i_weight_addr_gen_inst_N31, i_weight_addr_gen_inst_N30,
         i_weight_addr_gen_inst_N29, i_weight_addr_gen_inst_N28,
         i_weight_addr_gen_inst_N27, i_weight_addr_gen_inst_N26,
         i_weight_addr_gen_inst_N25, i_weight_addr_gen_inst_N24,
         i_weight_addr_gen_inst_N23, i_weight_addr_gen_inst_N22,
         i_weight_addr_gen_inst_N21, i_weight_addr_gen_inst_N20,
         i_weight_addr_gen_inst_N19, i_weight_addr_gen_inst_N18,
         i_weight_addr_gen_inst_N17, i_weight_addr_gen_inst_N16,
         i_weight_addr_gen_inst_N15, i_weight_addr_gen_inst_N14,
         i_weight_addr_gen_inst_N13, i_weight_addr_gen_inst_N12,
         i_weight_addr_gen_inst_N11, i_weight_addr_gen_inst_N10,
         i_weight_addr_gen_inst_int_offs_addr_1_,
         i_weight_addr_gen_inst_int_offs_addr_2_,
         i_weight_addr_gen_inst_int_offs_addr_3_,
         i_weight_addr_gen_inst_int_offs_addr_4_,
         i_weight_addr_gen_inst_int_offs_addr_5_,
         i_weight_addr_gen_inst_int_offs_addr_6_,
         i_weight_addr_gen_inst_int_offs_addr_7_,
         i_weight_addr_gen_inst_int_offs_addr_8_,
         i_weight_addr_gen_inst_int_offs_addr_9_,
         i_weight_addr_gen_inst_int_offs_addr_10_,
         i_weight_addr_gen_inst_int_offs_addr_11_,
         i_weight_addr_gen_inst_int_offs_addr_12_,
         i_weight_addr_gen_inst_int_offs_addr_13_,
         i_weight_addr_gen_inst_int_offs_addr_14_,
         i_weight_addr_gen_inst_int_offs_addr_15_,
         i_weight_addr_gen_inst_int_base_addr_0_,
         i_weight_addr_gen_inst_int_base_addr_1_,
         i_weight_addr_gen_inst_int_base_addr_2_,
         i_weight_addr_gen_inst_int_base_addr_3_,
         i_weight_addr_gen_inst_int_base_addr_4_,
         i_weight_addr_gen_inst_int_base_addr_5_,
         i_weight_addr_gen_inst_int_base_addr_6_,
         i_weight_addr_gen_inst_int_base_addr_7_,
         i_weight_addr_gen_inst_int_base_addr_8_,
         i_weight_addr_gen_inst_int_base_addr_9_,
         i_weight_addr_gen_inst_int_base_addr_10_,
         i_weight_addr_gen_inst_int_base_addr_11_,
         i_weight_addr_gen_inst_int_base_addr_12_,
         i_weight_addr_gen_inst_int_base_addr_13_,
         i_weight_addr_gen_inst_int_base_addr_14_,
         i_weight_addr_gen_inst_int_base_addr_15_,
         i_weight_addr_gen_inst_add_61_n1, i_weight_addr_gen_inst_add_46_n2,
         i_weight_addr_gen_inst_add_44_n2, i_weight_addr_gen_inst_add_32_n33,
         i_weight_addr_gen_inst_add_32_n32, i_weight_addr_gen_inst_add_32_n31,
         i_weight_addr_gen_inst_add_32_n30, i_weight_addr_gen_inst_add_32_n29,
         i_weight_addr_gen_inst_add_32_n28, i_weight_addr_gen_inst_add_32_n27,
         i_weight_addr_gen_inst_add_32_n26, i_weight_addr_gen_inst_add_32_n25,
         i_weight_addr_gen_inst_add_32_n24, i_weight_addr_gen_inst_add_32_n23,
         i_weight_addr_gen_inst_add_32_n22, i_weight_addr_gen_inst_add_32_n21,
         i_weight_addr_gen_inst_add_32_n20, i_weight_addr_gen_inst_add_32_n19,
         i_weight_addr_gen_inst_add_32_n18, i_weight_addr_gen_inst_add_32_n17,
         i_weight_addr_gen_inst_add_32_n16, i_weight_addr_gen_inst_add_32_n15,
         i_weight_addr_gen_inst_add_32_n14, i_weight_addr_gen_inst_add_32_n13,
         i_weight_addr_gen_inst_add_32_n12, i_weight_addr_gen_inst_add_32_n11,
         i_weight_addr_gen_inst_add_32_n10, i_weight_addr_gen_inst_add_32_n9,
         i_weight_addr_gen_inst_add_32_n8, i_weight_addr_gen_inst_add_32_n7,
         i_weight_addr_gen_inst_add_32_n6, i_weight_addr_gen_inst_add_32_n5,
         i_weight_addr_gen_inst_add_32_n4, i_weight_addr_gen_inst_add_32_n3,
         i_weight_addr_gen_inst_add_32_n2, i_weight_addr_gen_inst_add_32_n1,
         i_weight_addr_gen_inst_add_32_carry_2_,
         i_weight_addr_gen_inst_add_32_carry_3_,
         i_weight_addr_gen_inst_add_32_carry_4_,
         i_weight_addr_gen_inst_add_32_carry_5_,
         i_weight_addr_gen_inst_add_32_carry_6_,
         i_weight_addr_gen_inst_add_32_carry_7_,
         i_weight_addr_gen_inst_add_32_carry_8_,
         i_weight_addr_gen_inst_add_32_carry_9_,
         i_weight_addr_gen_inst_add_32_carry_10_,
         i_weight_addr_gen_inst_add_32_carry_11_,
         i_weight_addr_gen_inst_add_32_carry_12_,
         i_weight_addr_gen_inst_add_32_carry_13_,
         i_weight_addr_gen_inst_add_32_carry_14_,
         i_weight_addr_gen_inst_add_32_carry_15_,
         i_data_even_addr_gen_inst_n28, i_data_even_addr_gen_inst_n27,
         i_data_even_addr_gen_inst_n26, i_data_even_addr_gen_inst_n25,
         i_data_even_addr_gen_inst_n24, i_data_even_addr_gen_inst_n23,
         i_data_even_addr_gen_inst_n22, i_data_even_addr_gen_inst_n21,
         i_data_even_addr_gen_inst_n20, i_data_even_addr_gen_inst_n18,
         i_data_even_addr_gen_inst_n8, i_data_even_addr_gen_inst_n7,
         i_data_even_addr_gen_inst_n6, i_data_even_addr_gen_inst_n5,
         i_data_even_addr_gen_inst_n43, i_data_even_addr_gen_inst_n42,
         i_data_even_addr_gen_inst_n41, i_data_even_addr_gen_inst_n40,
         i_data_even_addr_gen_inst_n39, i_data_even_addr_gen_inst_n38,
         i_data_even_addr_gen_inst_n37, i_data_even_addr_gen_inst_n36,
         i_data_even_addr_gen_inst_n35, i_data_even_addr_gen_inst_n34,
         i_data_even_addr_gen_inst_n33, i_data_even_addr_gen_inst_n32,
         i_data_even_addr_gen_inst_net2809, i_data_even_addr_gen_inst_net2803,
         i_data_even_addr_gen_inst_N65, i_data_even_addr_gen_inst_N64,
         i_data_even_addr_gen_inst_N63, i_data_even_addr_gen_inst_N62,
         i_data_even_addr_gen_inst_N61, i_data_even_addr_gen_inst_N60,
         i_data_even_addr_gen_inst_N59, i_data_even_addr_gen_inst_N58,
         i_data_even_addr_gen_inst_N57, i_data_even_addr_gen_inst_N56,
         i_data_even_addr_gen_inst_N55, i_data_even_addr_gen_inst_N40,
         i_data_even_addr_gen_inst_N29, i_data_even_addr_gen_inst_N28,
         i_data_even_addr_gen_inst_N27, i_data_even_addr_gen_inst_N26,
         i_data_even_addr_gen_inst_N25, i_data_even_addr_gen_inst_N24,
         i_data_even_addr_gen_inst_N23, i_data_even_addr_gen_inst_N22,
         i_data_even_addr_gen_inst_N21, i_data_even_addr_gen_inst_N20,
         i_data_even_addr_gen_inst_N19, i_data_even_addr_gen_inst_N18,
         i_data_even_addr_gen_inst_N17, i_data_even_addr_gen_inst_N16,
         i_data_even_addr_gen_inst_N15, i_data_even_addr_gen_inst_N14,
         i_data_even_addr_gen_inst_N13, i_data_even_addr_gen_inst_N12,
         i_data_even_addr_gen_inst_N11, i_data_even_addr_gen_inst_N10,
         i_data_even_addr_gen_inst_int_offs_addr_0_,
         i_data_even_addr_gen_inst_int_offs_addr_1_,
         i_data_even_addr_gen_inst_int_offs_addr_2_,
         i_data_even_addr_gen_inst_int_offs_addr_3_,
         i_data_even_addr_gen_inst_int_offs_addr_4_,
         i_data_even_addr_gen_inst_int_offs_addr_5_,
         i_data_even_addr_gen_inst_int_offs_addr_6_,
         i_data_even_addr_gen_inst_int_offs_addr_7_,
         i_data_even_addr_gen_inst_int_offs_addr_8_,
         i_data_even_addr_gen_inst_int_offs_addr_9_,
         i_data_even_addr_gen_inst_int_base_addr_0_,
         i_data_even_addr_gen_inst_int_base_addr_1_,
         i_data_even_addr_gen_inst_int_base_addr_2_,
         i_data_even_addr_gen_inst_int_base_addr_3_,
         i_data_even_addr_gen_inst_int_base_addr_4_,
         i_data_even_addr_gen_inst_int_base_addr_5_,
         i_data_even_addr_gen_inst_int_base_addr_6_,
         i_data_even_addr_gen_inst_int_base_addr_7_,
         i_data_even_addr_gen_inst_int_base_addr_8_,
         i_data_even_addr_gen_inst_int_base_addr_9_,
         i_data_even_addr_gen_inst_add_61_n1,
         i_data_even_addr_gen_inst_add_46_n2,
         i_data_even_addr_gen_inst_add_44_n2,
         i_data_even_addr_gen_inst_add_32_n2, i_data_odd_addr_gen_inst_n28,
         i_data_odd_addr_gen_inst_n27, i_data_odd_addr_gen_inst_n26,
         i_data_odd_addr_gen_inst_n25, i_data_odd_addr_gen_inst_n24,
         i_data_odd_addr_gen_inst_n23, i_data_odd_addr_gen_inst_n22,
         i_data_odd_addr_gen_inst_n21, i_data_odd_addr_gen_inst_n20,
         i_data_odd_addr_gen_inst_n18, i_data_odd_addr_gen_inst_n8,
         i_data_odd_addr_gen_inst_n7, i_data_odd_addr_gen_inst_n6,
         i_data_odd_addr_gen_inst_n5, i_data_odd_addr_gen_inst_n43,
         i_data_odd_addr_gen_inst_n42, i_data_odd_addr_gen_inst_n41,
         i_data_odd_addr_gen_inst_n40, i_data_odd_addr_gen_inst_n39,
         i_data_odd_addr_gen_inst_n38, i_data_odd_addr_gen_inst_n37,
         i_data_odd_addr_gen_inst_n36, i_data_odd_addr_gen_inst_n35,
         i_data_odd_addr_gen_inst_n34, i_data_odd_addr_gen_inst_n33,
         i_data_odd_addr_gen_inst_n32, i_data_odd_addr_gen_inst_net2786,
         i_data_odd_addr_gen_inst_net2780, i_data_odd_addr_gen_inst_N65,
         i_data_odd_addr_gen_inst_N64, i_data_odd_addr_gen_inst_N63,
         i_data_odd_addr_gen_inst_N62, i_data_odd_addr_gen_inst_N61,
         i_data_odd_addr_gen_inst_N60, i_data_odd_addr_gen_inst_N59,
         i_data_odd_addr_gen_inst_N58, i_data_odd_addr_gen_inst_N57,
         i_data_odd_addr_gen_inst_N56, i_data_odd_addr_gen_inst_N55,
         i_data_odd_addr_gen_inst_N40, i_data_odd_addr_gen_inst_N29,
         i_data_odd_addr_gen_inst_N28, i_data_odd_addr_gen_inst_N27,
         i_data_odd_addr_gen_inst_N26, i_data_odd_addr_gen_inst_N25,
         i_data_odd_addr_gen_inst_N24, i_data_odd_addr_gen_inst_N23,
         i_data_odd_addr_gen_inst_N22, i_data_odd_addr_gen_inst_N21,
         i_data_odd_addr_gen_inst_N20, i_data_odd_addr_gen_inst_N19,
         i_data_odd_addr_gen_inst_N18, i_data_odd_addr_gen_inst_N17,
         i_data_odd_addr_gen_inst_N16, i_data_odd_addr_gen_inst_N15,
         i_data_odd_addr_gen_inst_N14, i_data_odd_addr_gen_inst_N13,
         i_data_odd_addr_gen_inst_N12, i_data_odd_addr_gen_inst_N11,
         i_data_odd_addr_gen_inst_N10,
         i_data_odd_addr_gen_inst_int_offs_addr_0_,
         i_data_odd_addr_gen_inst_int_offs_addr_1_,
         i_data_odd_addr_gen_inst_int_offs_addr_2_,
         i_data_odd_addr_gen_inst_int_offs_addr_3_,
         i_data_odd_addr_gen_inst_int_offs_addr_4_,
         i_data_odd_addr_gen_inst_int_offs_addr_5_,
         i_data_odd_addr_gen_inst_int_offs_addr_6_,
         i_data_odd_addr_gen_inst_int_offs_addr_7_,
         i_data_odd_addr_gen_inst_int_offs_addr_8_,
         i_data_odd_addr_gen_inst_int_offs_addr_9_,
         i_data_odd_addr_gen_inst_int_base_addr_0_,
         i_data_odd_addr_gen_inst_int_base_addr_1_,
         i_data_odd_addr_gen_inst_int_base_addr_2_,
         i_data_odd_addr_gen_inst_int_base_addr_3_,
         i_data_odd_addr_gen_inst_int_base_addr_4_,
         i_data_odd_addr_gen_inst_int_base_addr_5_,
         i_data_odd_addr_gen_inst_int_base_addr_6_,
         i_data_odd_addr_gen_inst_int_base_addr_7_,
         i_data_odd_addr_gen_inst_int_base_addr_8_,
         i_data_odd_addr_gen_inst_int_base_addr_9_,
         i_data_odd_addr_gen_inst_add_61_n1,
         i_data_odd_addr_gen_inst_add_46_n2,
         i_data_odd_addr_gen_inst_add_44_n2,
         i_data_odd_addr_gen_inst_add_32_n2, add_554_n1, add_553_n1;
  wire   [2:0] int_npu_ptr;
  wire   [2:0] int_ifmaps_ptr;
  wire   [2:0] ps_int_ifmaps_ptr;
  wire   [2:0] ps_int_hmode_cnt;
  wire   [15:0] int_i_data_h_npu;
  wire   [15:0] int_i_data_v_npu;
  wire   [2:0] int_hmode_cnt;
  wire   [1:7] int_ckg_rmask;
  wire   [1:7] int_ckg_cmask;
  wire   [63:0] int_o_data_npu;
  wire   [15:0] int_o_data_p;
  wire   [2:0] int_arv_res;
  wire   [2:0] int_d_tc;
  wire   [9:0] int_o_data_even_base_addr;
  wire   [9:0] int_o_data_odd_base_addr;
  wire   [9:0] int_o_data_even_offs_addr;
  wire   [9:0] int_o_data_odd_offs_addr;
  wire   [9:1] add_1_root_add_546_2_carry;
  wire   [9:1] add_1_root_add_544_2_carry;
  wire   [7:0] wrap_act_buffer_inst_int_i_data_if8;
  wire   [7:0] wrap_act_buffer_inst_int_i_data_if7;
  wire   [7:0] wrap_act_buffer_inst_int_i_data_if6;
  wire   [7:0] wrap_act_buffer_inst_int_i_data_if5;
  wire   [7:0] wrap_act_buffer_inst_int_i_data_if4;
  wire   [7:0] wrap_act_buffer_inst_int_i_data_if3;
  wire   [7:0] wrap_act_buffer_inst_int_i_data_if2;
  wire   [7:0] wrap_act_buffer_inst_int_i_data_if1;
  wire   [47:0] wrap_act_buffer_inst_act_buffer_inst_int_data8;
  wire   [47:0] wrap_act_buffer_inst_act_buffer_inst_int_data7;
  wire   [47:0] wrap_act_buffer_inst_act_buffer_inst_int_data6;
  wire   [47:0] wrap_act_buffer_inst_act_buffer_inst_int_data5;
  wire   [47:0] wrap_act_buffer_inst_act_buffer_inst_int_data4;
  wire   [47:0] wrap_act_buffer_inst_act_buffer_inst_int_data3;
  wire   [47:0] wrap_act_buffer_inst_act_buffer_inst_int_data2;
  wire   [47:0] wrap_act_buffer_inst_act_buffer_inst_int_data1;
  wire   [7:0] wrap_act_buffer_inst_act_if_inst_int_data8;
  wire   [7:0] wrap_act_buffer_inst_act_if_inst_int_data7;
  wire   [7:0] wrap_act_buffer_inst_act_if_inst_int_data6;
  wire   [7:0] wrap_act_buffer_inst_act_if_inst_int_data5;
  wire   [7:0] wrap_act_buffer_inst_act_if_inst_int_data4;
  wire   [7:0] wrap_act_buffer_inst_act_if_inst_int_data3;
  wire   [7:0] wrap_act_buffer_inst_act_if_inst_int_data2;
  wire   [7:0] wrap_act_buffer_inst_act_if_inst_int_data1;
  wire   [63:0] npu_inst_int_ckg;
  wire   [15:2] i_weight_addr_gen_inst_add_61_carry;
  wire   [15:2] i_weight_addr_gen_inst_add_46_carry;
  wire   [15:2] i_weight_addr_gen_inst_add_44_carry;
  wire   [9:2] i_data_even_addr_gen_inst_add_61_carry;
  wire   [9:2] i_data_even_addr_gen_inst_add_46_carry;
  wire   [9:2] i_data_even_addr_gen_inst_add_44_carry;
  wire   [9:2] i_data_even_addr_gen_inst_add_32_carry;
  wire   [9:2] i_data_odd_addr_gen_inst_add_61_carry;
  wire   [9:2] i_data_odd_addr_gen_inst_add_46_carry;
  wire   [9:2] i_data_odd_addr_gen_inst_add_44_carry;
  wire   [9:2] i_data_odd_addr_gen_inst_add_32_carry;
  wire   [9:2] add_554_carry;
  wire   [9:2] add_553_carry;
  wire   [9:2] add_539_carry;
  wire   [9:2] add_538_carry;

  DFFR_X1 ps_ctrl_wr_mem_reg ( .D(ctrl_wr_mem), .CK(ck), .RN(n52), .Q(
        o_data_wr), .QN(n16) );
  DFFR_X1 ps_ctrl_en_npu_reg ( .D(ctrl_en_npu), .CK(ck), .RN(n52), .Q(
        ps_ctrl_en_npu) );
  DFFR_X1 ps_ctrl_ldh_v_n_reg ( .D(ctrl_ldh_v_n), .CK(ck), .RN(n52), .Q(
        ps_ctrl_ldh_v_n) );
  DFFR_X1 ps_ctrl_wr_pipe_reg ( .D(ctrl_wr_pipe), .CK(ck), .RN(n52), .Q(
        ps_ctrl_wr_pipe) );
  DFFR_X1 ps_ctrl_en_p_reg ( .D(ctrl_en_p), .CK(ck), .RN(n52), .Q(ps_ctrl_en_p) );
  DFFR_X1 ps_int_ifmaps_ptr_reg_2_ ( .D(int_ifmaps_ptr[2]), .CK(ck), .RN(n52), 
        .Q(ps_int_ifmaps_ptr[2]) );
  DFFR_X1 ps_int_ifmaps_ptr_reg_1_ ( .D(int_ifmaps_ptr[1]), .CK(ck), .RN(n52), 
        .Q(ps_int_ifmaps_ptr[1]) );
  DFFR_X1 ps_int_ifmaps_ptr_reg_0_ ( .D(int_ifmaps_ptr[0]), .CK(ck), .RN(n52), 
        .Q(ps_int_ifmaps_ptr[0]) );
  DFFR_X1 ps_int_hmode_cnt_reg_2_ ( .D(int_hmode_cnt[2]), .CK(ck), .RN(n52), 
        .Q(ps_int_hmode_cnt[2]) );
  DFFR_X1 ps_int_hmode_cnt_reg_1_ ( .D(int_hmode_cnt[1]), .CK(ck), .RN(n52), 
        .Q(ps_int_hmode_cnt[1]) );
  DFFR_X1 ps_int_hmode_cnt_reg_0_ ( .D(int_hmode_cnt[0]), .CK(ck), .RN(n52), 
        .Q(ps_int_hmode_cnt[0]) );
  DFFR_X1 int_q_tc_reg_2_ ( .D(int_d_tc[2]), .CK(net2747), .RN(n56), .Q(
        s_tc_tilev), .QN(n19) );
  DFFR_X1 int_q_tc_reg_1_ ( .D(int_d_tc[1]), .CK(net2747), .RN(n56), .Q(
        s_tc_tileh), .QN(n21) );
  DFFR_X1 int_q_tc_reg_0_ ( .D(int_d_tc[0]), .CK(net2747), .RN(n56), .Q(
        s_tc_ofmaps) );
  DFFR_X1 ps_int_s_tc_tileh_reg ( .D(s_tc_tileh), .CK(ck), .RN(n52), .Q(
        ps_int_s_tc_tileh) );
  DFFR_X1 ps_int_s_tc_res_reg ( .D(s_tc_res), .CK(ck), .RN(n53), .Q(
        ps_int_s_tc_res) );
  DFFR_X1 ps_int_s_tc_tilev_reg ( .D(s_tc_tilev), .CK(ck), .RN(n53), .Q(
        ps_int_s_tc_tilev) );
  DFFR_X1 int_o_data_even_base_addr_reg_0_ ( .D(N40), .CK(net2758), .RN(n56), 
        .Q(int_o_data_even_base_addr[0]) );
  DFFR_X1 int_o_data_even_base_addr_reg_1_ ( .D(N41), .CK(net2758), .RN(n56), 
        .Q(int_o_data_even_base_addr[1]) );
  DFFR_X1 int_o_data_even_base_addr_reg_2_ ( .D(N42), .CK(net2758), .RN(n56), 
        .Q(int_o_data_even_base_addr[2]) );
  DFFR_X1 int_o_data_even_base_addr_reg_3_ ( .D(N43), .CK(net2758), .RN(n56), 
        .Q(int_o_data_even_base_addr[3]) );
  DFFR_X1 int_o_data_even_base_addr_reg_4_ ( .D(N44), .CK(net2758), .RN(n56), 
        .Q(int_o_data_even_base_addr[4]) );
  DFFR_X1 int_o_data_even_base_addr_reg_5_ ( .D(N45), .CK(net2758), .RN(n56), 
        .Q(int_o_data_even_base_addr[5]) );
  DFFR_X1 int_o_data_even_base_addr_reg_6_ ( .D(N46), .CK(net2758), .RN(n56), 
        .Q(int_o_data_even_base_addr[6]) );
  DFFR_X1 int_o_data_even_base_addr_reg_7_ ( .D(N47), .CK(net2758), .RN(n56), 
        .Q(int_o_data_even_base_addr[7]) );
  DFFR_X1 int_o_data_even_base_addr_reg_8_ ( .D(N48), .CK(net2758), .RN(n55), 
        .Q(int_o_data_even_base_addr[8]) );
  DFFR_X1 int_o_data_even_base_addr_reg_9_ ( .D(N49), .CK(net2758), .RN(n55), 
        .Q(int_o_data_even_base_addr[9]) );
  DFFR_X1 int_o_data_odd_base_addr_reg_0_ ( .D(N50), .CK(net2758), .RN(n55), 
        .Q(int_o_data_odd_base_addr[0]) );
  DFFR_X1 int_o_data_odd_base_addr_reg_1_ ( .D(N51), .CK(net2758), .RN(n55), 
        .Q(int_o_data_odd_base_addr[1]) );
  DFFR_X1 int_o_data_odd_base_addr_reg_2_ ( .D(N52), .CK(net2758), .RN(n55), 
        .Q(int_o_data_odd_base_addr[2]) );
  DFFR_X1 int_o_data_odd_base_addr_reg_3_ ( .D(N53), .CK(net2758), .RN(n55), 
        .Q(int_o_data_odd_base_addr[3]) );
  DFFR_X1 int_o_data_odd_base_addr_reg_4_ ( .D(N54), .CK(net2758), .RN(n55), 
        .Q(int_o_data_odd_base_addr[4]) );
  DFFR_X1 int_o_data_odd_base_addr_reg_5_ ( .D(N55), .CK(net2758), .RN(n55), 
        .Q(int_o_data_odd_base_addr[5]) );
  DFFR_X1 int_o_data_odd_base_addr_reg_6_ ( .D(N56), .CK(net2758), .RN(n55), 
        .Q(int_o_data_odd_base_addr[6]) );
  DFFR_X1 int_o_data_odd_base_addr_reg_7_ ( .D(N57), .CK(net2758), .RN(n55), 
        .Q(int_o_data_odd_base_addr[7]) );
  DFFR_X1 int_o_data_odd_base_addr_reg_8_ ( .D(N58), .CK(net2758), .RN(n55), 
        .Q(int_o_data_odd_base_addr[8]) );
  DFFR_X1 int_o_data_odd_base_addr_reg_9_ ( .D(N59), .CK(net2758), .RN(n55), 
        .Q(int_o_data_odd_base_addr[9]) );
  DFFR_X1 int_o_data_wrh_l_n_reg ( .D(n44), .CK(ck), .RN(n53), .Q(
        o_data_wrh_l_n) );
  DFFR_X1 int_o_data_ev_odd_n_reg ( .D(n58), .CK(ck), .RN(n53), .Q(
        o_data_ev_odd_n), .QN(n26) );
  DFFR_X1 int_o_data_odd_offs_addr_reg_0_ ( .D(N113), .CK(net2753), .RN(n54), 
        .Q(int_o_data_odd_offs_addr[0]) );
  DFFR_X1 int_o_data_odd_offs_addr_reg_1_ ( .D(N114), .CK(net2753), .RN(n54), 
        .Q(int_o_data_odd_offs_addr[1]) );
  DFFR_X1 int_o_data_odd_offs_addr_reg_2_ ( .D(N115), .CK(net2753), .RN(n54), 
        .Q(int_o_data_odd_offs_addr[2]) );
  DFFR_X1 int_o_data_odd_offs_addr_reg_3_ ( .D(N116), .CK(net2753), .RN(n54), 
        .Q(int_o_data_odd_offs_addr[3]) );
  DFFR_X1 int_o_data_odd_offs_addr_reg_4_ ( .D(N117), .CK(net2753), .RN(n54), 
        .Q(int_o_data_odd_offs_addr[4]) );
  DFFR_X1 int_o_data_odd_offs_addr_reg_5_ ( .D(N118), .CK(net2753), .RN(n54), 
        .Q(int_o_data_odd_offs_addr[5]) );
  DFFR_X1 int_o_data_odd_offs_addr_reg_6_ ( .D(N119), .CK(net2753), .RN(n54), 
        .Q(int_o_data_odd_offs_addr[6]) );
  DFFR_X1 int_o_data_odd_offs_addr_reg_7_ ( .D(N120), .CK(net2753), .RN(n54), 
        .Q(int_o_data_odd_offs_addr[7]) );
  DFFR_X1 int_o_data_odd_offs_addr_reg_8_ ( .D(N121), .CK(net2753), .RN(n54), 
        .Q(int_o_data_odd_offs_addr[8]) );
  DFFR_X1 int_o_data_odd_offs_addr_reg_9_ ( .D(N122), .CK(net2753), .RN(n54), 
        .Q(int_o_data_odd_offs_addr[9]) );
  DFFR_X1 int_o_data_even_offs_addr_reg_0_ ( .D(N102), .CK(net2763), .RN(n54), 
        .Q(int_o_data_even_offs_addr[0]) );
  DFFR_X1 int_o_data_even_offs_addr_reg_1_ ( .D(N103), .CK(net2763), .RN(n54), 
        .Q(int_o_data_even_offs_addr[1]) );
  DFFR_X1 int_o_data_even_offs_addr_reg_2_ ( .D(N104), .CK(net2763), .RN(n53), 
        .Q(int_o_data_even_offs_addr[2]) );
  DFFR_X1 int_o_data_even_offs_addr_reg_3_ ( .D(N105), .CK(net2763), .RN(n53), 
        .Q(int_o_data_even_offs_addr[3]) );
  DFFR_X1 int_o_data_even_offs_addr_reg_4_ ( .D(N106), .CK(net2763), .RN(n53), 
        .Q(int_o_data_even_offs_addr[4]) );
  DFFR_X1 int_o_data_even_offs_addr_reg_5_ ( .D(N107), .CK(net2763), .RN(n53), 
        .Q(int_o_data_even_offs_addr[5]) );
  DFFR_X1 int_o_data_even_offs_addr_reg_6_ ( .D(N108), .CK(net2763), .RN(n53), 
        .Q(int_o_data_even_offs_addr[6]) );
  DFFR_X1 int_o_data_even_offs_addr_reg_7_ ( .D(N109), .CK(net2763), .RN(n53), 
        .Q(int_o_data_even_offs_addr[7]) );
  DFFR_X1 int_o_data_even_offs_addr_reg_8_ ( .D(N110), .CK(net2763), .RN(n53), 
        .Q(int_o_data_even_offs_addr[8]) );
  DFFR_X1 int_o_data_even_offs_addr_reg_9_ ( .D(N111), .CK(net2763), .RN(n53), 
        .Q(int_o_data_even_offs_addr[9]) );
  NAND3_X1 U79 ( .A1(n65), .A2(n61), .A3(n66), .ZN(n39) );
  FA_X1 add_1_root_add_546_2_U1_1 ( .A(int_o_data_odd_offs_addr[1]), .B(
        arv_ofmaps[1]), .CI(add_1_root_add_546_2_carry[1]), .CO(
        add_1_root_add_546_2_carry[2]), .S(N92) );
  FA_X1 add_1_root_add_546_2_U1_2 ( .A(int_o_data_odd_offs_addr[2]), .B(
        arv_ofmaps[2]), .CI(add_1_root_add_546_2_carry[2]), .CO(
        add_1_root_add_546_2_carry[3]), .S(N93) );
  FA_X1 add_1_root_add_546_2_U1_3 ( .A(int_o_data_odd_offs_addr[3]), .B(
        arv_ofmaps[3]), .CI(add_1_root_add_546_2_carry[3]), .CO(
        add_1_root_add_546_2_carry[4]), .S(N94) );
  FA_X1 add_1_root_add_544_2_U1_1 ( .A(int_o_data_even_offs_addr[1]), .B(
        arv_ofmaps[1]), .CI(add_1_root_add_544_2_carry[1]), .CO(
        add_1_root_add_544_2_carry[2]), .S(N72) );
  FA_X1 add_1_root_add_544_2_U1_2 ( .A(int_o_data_even_offs_addr[2]), .B(
        arv_ofmaps[2]), .CI(add_1_root_add_544_2_carry[2]), .CO(
        add_1_root_add_544_2_carry[3]), .S(N73) );
  FA_X1 add_1_root_add_544_2_U1_3 ( .A(int_o_data_even_offs_addr[3]), .B(
        arv_ofmaps[3]), .CI(add_1_root_add_544_2_carry[3]), .CO(
        add_1_root_add_544_2_carry[4]), .S(N74) );
  INV_X1 U80 ( .A(n42), .ZN(n59) );
  AND2_X1 U81 ( .A1(int_d_tc[1]), .A2(n59), .ZN(int_en_ofmaps_ptr) );
  NOR3_X1 U82 ( .A1(n66), .A2(n65), .A3(n37), .ZN(n35) );
  NOR2_X1 U83 ( .A1(n57), .A2(n42), .ZN(int_c_i_en_odd) );
  INV_X1 U84 ( .A(n36), .ZN(n64) );
  AOI21_X1 U85 ( .B1(n61), .B2(n66), .A(n41), .ZN(n38) );
  AND2_X1 U86 ( .A1(s_tc_npu_ptr), .A2(int_en_npu_ptr), .ZN(int_en_tilev_ptr)
         );
  NAND2_X1 U87 ( .A1(int_d_tc[2]), .A2(int_en_tilev_ptr), .ZN(n42) );
  INV_X1 U88 ( .A(s_tc_res), .ZN(n60) );
  INV_X1 U89 ( .A(n41), .ZN(n62) );
  NAND2_X1 U90 ( .A1(n36), .A2(int_arv_res[1]), .ZN(int_ckg_rmask[6]) );
  INV_X1 U91 ( .A(n40), .ZN(n63) );
  AND2_X1 U92 ( .A1(N74), .A2(n43), .ZN(N105) );
  AND2_X1 U93 ( .A1(N94), .A2(n43), .ZN(N116) );
  INV_X1 U94 ( .A(n32), .ZN(n68) );
  INV_X1 U95 ( .A(N124), .ZN(n67) );
  AND2_X1 U96 ( .A1(N73), .A2(n45), .ZN(N104) );
  AND2_X1 U97 ( .A1(N93), .A2(n45), .ZN(N115) );
  AND2_X1 U98 ( .A1(N72), .A2(n43), .ZN(N103) );
  AND2_X1 U99 ( .A1(N92), .A2(n43), .ZN(N114) );
  BUF_X1 U100 ( .A(n51), .Z(n46) );
  BUF_X1 U101 ( .A(n50), .Z(n48) );
  BUF_X1 U102 ( .A(n51), .Z(n47) );
  BUF_X1 U103 ( .A(n50), .Z(n49) );
  NOR3_X1 U104 ( .A1(n60), .A2(n19), .A3(n21), .ZN(int_c_i_en_weight_addr) );
  OAI21_X1 U105 ( .B1(arv_ckg[1]), .B2(n21), .A(n40), .ZN(int_ckg_cmask[6]) );
  NOR2_X1 U106 ( .A1(n35), .A2(n21), .ZN(int_ckg_cmask[7]) );
  NOR2_X1 U107 ( .A1(n38), .A2(n21), .ZN(int_ckg_cmask[3]) );
  NOR2_X1 U108 ( .A1(n62), .A2(n21), .ZN(int_ckg_cmask[2]) );
  NOR2_X1 U109 ( .A1(n39), .A2(n21), .ZN(int_ckg_cmask[1]) );
  NOR2_X1 U110 ( .A1(i_data_ev_odd_n), .A2(n42), .ZN(int_c_i_en_even) );
  OAI21_X1 U111 ( .B1(arv_ckg[1]), .B2(arv_ckg[0]), .A(arv_ckg[2]), .ZN(n37)
         );
  NOR2_X1 U112 ( .A1(n35), .A2(n19), .ZN(int_ckg_rmask[7]) );
  NOR2_X1 U113 ( .A1(n38), .A2(n19), .ZN(int_ckg_rmask[3]) );
  NOR2_X1 U114 ( .A1(n19), .A2(n62), .ZN(int_ckg_rmask[2]) );
  NOR2_X1 U115 ( .A1(n19), .A2(n39), .ZN(int_ckg_rmask[1]) );
  NOR2_X1 U116 ( .A1(arv_ckg[1]), .A2(arv_ckg[2]), .ZN(n41) );
  AND2_X1 U117 ( .A1(N77), .A2(n45), .ZN(N108) );
  AND2_X1 U118 ( .A1(N97), .A2(n45), .ZN(N119) );
  NAND2_X1 U119 ( .A1(s_tc_tilev), .A2(n65), .ZN(int_arv_res[1]) );
  INV_X1 U120 ( .A(arv_ckg[0]), .ZN(n66) );
  NAND2_X1 U121 ( .A1(s_tc_tilev), .A2(n37), .ZN(n36) );
  NAND2_X1 U122 ( .A1(s_tc_tilev), .A2(n66), .ZN(int_arv_res[0]) );
  NAND2_X1 U123 ( .A1(s_tc_tilev), .A2(n61), .ZN(int_arv_res[2]) );
  NAND2_X1 U124 ( .A1(s_tc_tileh), .A2(n37), .ZN(n40) );
  INV_X1 U125 ( .A(arv_ckg[1]), .ZN(n65) );
  INV_X1 U126 ( .A(arv_ckg[2]), .ZN(n61) );
  AND2_X1 U127 ( .A1(ctrl_ldh_v_n), .A2(s_tc_ifmaps), .ZN(int_en_npu_ptr) );
  AND2_X1 U128 ( .A1(N79), .A2(n45), .ZN(N110) );
  AND2_X1 U129 ( .A1(N75), .A2(n45), .ZN(N106) );
  AND2_X1 U130 ( .A1(N98), .A2(n45), .ZN(N120) );
  AND2_X1 U131 ( .A1(N95), .A2(n45), .ZN(N117) );
  AND2_X1 U132 ( .A1(N80), .A2(n43), .ZN(N111) );
  AND2_X1 U133 ( .A1(N78), .A2(n43), .ZN(N109) );
  AND2_X1 U134 ( .A1(N76), .A2(n43), .ZN(N107) );
  AND2_X1 U135 ( .A1(N100), .A2(n43), .ZN(N122) );
  AND2_X1 U136 ( .A1(N99), .A2(n43), .ZN(N121) );
  AND2_X1 U137 ( .A1(N96), .A2(n43), .ZN(N118) );
  NOR2_X1 U138 ( .A1(arv_ckg[2]), .A2(n21), .ZN(int_ckg_cmask[4]) );
  NOR2_X1 U139 ( .A1(arv_ckg[2]), .A2(n19), .ZN(int_ckg_rmask[4]) );
  NAND2_X1 U140 ( .A1(ps_int_s_tc_tileh), .A2(n68), .ZN(n45) );
  NAND2_X1 U141 ( .A1(ps_int_s_tc_tileh), .A2(n68), .ZN(n43) );
  NAND2_X1 U142 ( .A1(ps_int_s_tc_tilev), .A2(ps_int_s_tc_res), .ZN(n32) );
  NOR2_X1 U143 ( .A1(n45), .A2(n16), .ZN(N124) );
  INV_X1 U144 ( .A(i_data_ev_odd_n), .ZN(n57) );
  OAI21_X1 U145 ( .B1(n32), .B2(n57), .A(n33), .ZN(n44) );
  NAND2_X1 U146 ( .A1(o_data_wrh_l_n), .A2(n32), .ZN(n33) );
  OAI21_X1 U147 ( .B1(n26), .B2(n16), .A(n67), .ZN(N123) );
  OAI21_X1 U148 ( .B1(o_data_ev_odd_n), .B2(n16), .A(n67), .ZN(N125) );
  NAND2_X1 U149 ( .A1(n60), .A2(n34), .ZN(int_en_vmode) );
  NAND2_X1 U150 ( .A1(s_tc_ifmaps), .A2(ctrl_en_vmode), .ZN(n34) );
  AND2_X1 U151 ( .A1(N71), .A2(n45), .ZN(N102) );
  AND2_X1 U152 ( .A1(N91), .A2(n45), .ZN(N113) );
  INV_X1 U153 ( .A(n31), .ZN(n58) );
  AOI22_X1 U154 ( .A1(n68), .A2(int_tileh_ptr_1_), .B1(n32), .B2(
        o_data_ev_odd_n), .ZN(n31) );
  AND2_X1 U155 ( .A1(ctrl_en_hmode), .A2(s_tc_ifmaps), .ZN(int_en_hmode) );
  BUF_X1 U156 ( .A(rst), .Z(n51) );
  BUF_X1 U157 ( .A(rst), .Z(n50) );
  INV_X1 U158 ( .A(n49), .ZN(n52) );
  INV_X1 U159 ( .A(n48), .ZN(n53) );
  INV_X1 U160 ( .A(n49), .ZN(n54) );
  INV_X1 U161 ( .A(n48), .ZN(n55) );
  INV_X1 U162 ( .A(n48), .ZN(n56) );
  XOR2_X1 U163 ( .A(int_o_data_even_offs_addr[9]), .B(
        add_1_root_add_544_2_carry[9]), .Z(N80) );
  AND2_X1 U164 ( .A1(add_1_root_add_544_2_carry[8]), .A2(
        int_o_data_even_offs_addr[8]), .ZN(add_1_root_add_544_2_carry[9]) );
  XOR2_X1 U165 ( .A(int_o_data_even_offs_addr[8]), .B(
        add_1_root_add_544_2_carry[8]), .Z(N79) );
  AND2_X1 U166 ( .A1(add_1_root_add_544_2_carry[7]), .A2(
        int_o_data_even_offs_addr[7]), .ZN(add_1_root_add_544_2_carry[8]) );
  XOR2_X1 U167 ( .A(int_o_data_even_offs_addr[7]), .B(
        add_1_root_add_544_2_carry[7]), .Z(N78) );
  AND2_X1 U168 ( .A1(add_1_root_add_544_2_carry[6]), .A2(
        int_o_data_even_offs_addr[6]), .ZN(add_1_root_add_544_2_carry[7]) );
  XOR2_X1 U169 ( .A(int_o_data_even_offs_addr[6]), .B(
        add_1_root_add_544_2_carry[6]), .Z(N77) );
  AND2_X1 U170 ( .A1(add_1_root_add_544_2_carry[5]), .A2(
        int_o_data_even_offs_addr[5]), .ZN(add_1_root_add_544_2_carry[6]) );
  XOR2_X1 U171 ( .A(int_o_data_even_offs_addr[5]), .B(
        add_1_root_add_544_2_carry[5]), .Z(N76) );
  AND2_X1 U172 ( .A1(add_1_root_add_544_2_carry[4]), .A2(
        int_o_data_even_offs_addr[4]), .ZN(add_1_root_add_544_2_carry[5]) );
  XOR2_X1 U173 ( .A(int_o_data_even_offs_addr[4]), .B(
        add_1_root_add_544_2_carry[4]), .Z(N75) );
  OR2_X1 U174 ( .A1(arv_ofmaps[0]), .A2(int_o_data_even_offs_addr[0]), .ZN(
        add_1_root_add_544_2_carry[1]) );
  XNOR2_X1 U175 ( .A(int_o_data_even_offs_addr[0]), .B(arv_ofmaps[0]), .ZN(N71) );
  XOR2_X1 U176 ( .A(int_o_data_odd_offs_addr[9]), .B(
        add_1_root_add_546_2_carry[9]), .Z(N100) );
  AND2_X1 U177 ( .A1(add_1_root_add_546_2_carry[8]), .A2(
        int_o_data_odd_offs_addr[8]), .ZN(add_1_root_add_546_2_carry[9]) );
  XOR2_X1 U178 ( .A(int_o_data_odd_offs_addr[8]), .B(
        add_1_root_add_546_2_carry[8]), .Z(N99) );
  AND2_X1 U179 ( .A1(add_1_root_add_546_2_carry[7]), .A2(
        int_o_data_odd_offs_addr[7]), .ZN(add_1_root_add_546_2_carry[8]) );
  XOR2_X1 U180 ( .A(int_o_data_odd_offs_addr[7]), .B(
        add_1_root_add_546_2_carry[7]), .Z(N98) );
  AND2_X1 U181 ( .A1(add_1_root_add_546_2_carry[6]), .A2(
        int_o_data_odd_offs_addr[6]), .ZN(add_1_root_add_546_2_carry[7]) );
  XOR2_X1 U182 ( .A(int_o_data_odd_offs_addr[6]), .B(
        add_1_root_add_546_2_carry[6]), .Z(N97) );
  AND2_X1 U183 ( .A1(add_1_root_add_546_2_carry[5]), .A2(
        int_o_data_odd_offs_addr[5]), .ZN(add_1_root_add_546_2_carry[6]) );
  XOR2_X1 U184 ( .A(int_o_data_odd_offs_addr[5]), .B(
        add_1_root_add_546_2_carry[5]), .Z(N96) );
  AND2_X1 U185 ( .A1(add_1_root_add_546_2_carry[4]), .A2(
        int_o_data_odd_offs_addr[4]), .ZN(add_1_root_add_546_2_carry[5]) );
  XOR2_X1 U186 ( .A(int_o_data_odd_offs_addr[4]), .B(
        add_1_root_add_546_2_carry[4]), .Z(N95) );
  OR2_X1 U187 ( .A1(arv_ofmaps[0]), .A2(int_o_data_odd_offs_addr[0]), .ZN(
        add_1_root_add_546_2_carry[1]) );
  XNOR2_X1 U188 ( .A(int_o_data_odd_offs_addr[0]), .B(arv_ofmaps[0]), .ZN(N91)
         );
  INV_X1 wrap_act_buffer_inst_U3 ( .A(n46), .ZN(wrap_act_buffer_inst_n2) );
  INV_X1 wrap_act_buffer_inst_U2 ( .A(n46), .ZN(wrap_act_buffer_inst_n1) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_0_ ( .D(i_actv[0]), .CK(
        wrap_act_buffer_inst_net4501), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[0]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_1_ ( .D(i_actv[1]), .CK(
        wrap_act_buffer_inst_net4501), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[1]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_2_ ( .D(i_actv[2]), .CK(
        wrap_act_buffer_inst_net4501), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[2]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_3_ ( .D(i_actv[3]), .CK(
        wrap_act_buffer_inst_net4501), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[3]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_4_ ( .D(i_actv[4]), .CK(
        wrap_act_buffer_inst_net4501), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[4]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_5_ ( .D(i_actv[5]), .CK(
        wrap_act_buffer_inst_net4501), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[5]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_6_ ( .D(i_actv[6]), .CK(
        wrap_act_buffer_inst_net4501), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[6]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_7_ ( .D(i_actv[7]), .CK(
        wrap_act_buffer_inst_net4501), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[7]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_8_ ( .D(i_actv[8]), .CK(
        wrap_act_buffer_inst_net4501), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[8]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_9_ ( .D(i_actv[9]), .CK(
        wrap_act_buffer_inst_net4501), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[9]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_10_ ( .D(i_actv[10]), .CK(
        wrap_act_buffer_inst_net4501), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[10]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_11_ ( .D(i_actv[11]), .CK(
        wrap_act_buffer_inst_net4501), .RN(wrap_act_buffer_inst_n1), .Q(
        int_i_data_v_npu[11]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_12_ ( .D(i_actv[12]), .CK(
        wrap_act_buffer_inst_net4501), .RN(wrap_act_buffer_inst_n2), .Q(
        int_i_data_v_npu[12]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_13_ ( .D(i_actv[13]), .CK(
        wrap_act_buffer_inst_net4501), .RN(wrap_act_buffer_inst_n2), .Q(
        int_i_data_v_npu[13]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_14_ ( .D(i_actv[14]), .CK(
        wrap_act_buffer_inst_net4501), .RN(wrap_act_buffer_inst_n2), .Q(
        int_i_data_v_npu[14]) );
  DFFR_X1 wrap_act_buffer_inst_int_i_data_v_npu_reg_15_ ( .D(i_actv[15]), .CK(
        wrap_act_buffer_inst_net4501), .RN(wrap_act_buffer_inst_n2), .Q(
        int_i_data_v_npu[15]) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U380 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n248), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n263) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U379 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n247), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n262) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U378 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n246), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n261) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U377 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n245), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n260) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U376 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n244), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n259) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U375 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n243), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n258) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U374 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n242), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n257) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U373 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n240), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n256) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U372 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n238), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n255) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U371 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n236), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n254) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U370 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n234), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n253) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U369 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n252) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U368 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n251) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U367 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n250) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U366 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n249) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U365 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n248) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U364 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n247) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U363 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n246) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U362 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n245) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U361 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n244) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U360 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n243) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U359 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n242) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U358 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n232), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n241) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U357 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n240) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U356 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n239) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U355 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n238) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U354 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n237) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U353 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n236) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U352 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n235) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U351 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n234) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U350 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n233) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U349 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n264), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n232) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U348 ( .A(i_acth[15]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n230) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U347 ( .A(i_acth[14]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n225) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U346 ( .A(i_acth[13]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n220) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U345 ( .A(i_acth[12]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n215) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U344 ( .A(i_acth[11]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n210) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U343 ( .A(i_acth[10]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n205) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U342 ( .A(i_acth[9]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n200) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U341 ( .A(i_acth[8]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n195) );
  INV_X1 wrap_act_buffer_inst_act_buffer_inst_U340 ( .A(ps_int_ifmaps_ptr[0]), 
        .ZN(wrap_act_buffer_inst_act_buffer_inst_n186) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U339 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n12), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n185) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U338 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n13), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n179) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U337 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n14), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n173) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U336 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n15), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n167) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U335 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n16), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n161) );
  CLKBUF_X1 wrap_act_buffer_inst_act_buffer_inst_U334 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n17), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n6) );
  INV_X1 wrap_act_buffer_inst_act_buffer_inst_U333 ( .A(int_npu_ptr[2]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n190) );
  INV_X1 wrap_act_buffer_inst_act_buffer_inst_U332 ( .A(int_npu_ptr[1]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n189) );
  INV_X1 wrap_act_buffer_inst_act_buffer_inst_U331 ( .A(int_npu_ptr[0]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n188) );
  INV_X1 wrap_act_buffer_inst_act_buffer_inst_U330 ( .A(int_ifmaps_ptr[0]), 
        .ZN(wrap_act_buffer_inst_act_buffer_inst_n265) );
  INV_X1 wrap_act_buffer_inst_act_buffer_inst_U329 ( .A(int_ifmaps_ptr[2]), 
        .ZN(wrap_act_buffer_inst_act_buffer_inst_n267) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U328 ( .A(i_acth[15]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n229) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U327 ( .A(i_acth[14]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n224) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U326 ( .A(i_acth[13]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n219) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U325 ( .A(i_acth[12]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n214) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U324 ( .A(i_acth[11]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n209) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U323 ( .A(i_acth[10]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n204) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U322 ( .A(i_acth[9]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n199) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U321 ( .A(i_acth[8]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n194) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U320 ( .A(i_acth[15]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n228) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U319 ( .A(i_acth[14]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n223) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U318 ( .A(i_acth[13]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n218) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U317 ( .A(i_acth[12]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n213) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U316 ( .A(i_acth[11]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n208) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U315 ( .A(i_acth[10]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n203) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U314 ( .A(i_acth[9]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n198) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U313 ( .A(i_acth[8]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n193) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U312 ( .A(i_acth[15]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n227) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U311 ( .A(i_acth[14]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n222) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U310 ( .A(i_acth[13]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n217) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U309 ( .A(i_acth[12]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n212) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U308 ( .A(i_acth[11]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n207) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U307 ( .A(i_acth[10]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n202) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U306 ( .A(i_acth[9]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n197) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U305 ( .A(i_acth[8]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n192) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U304 ( .A(i_acth[15]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n226) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U303 ( .A(i_acth[14]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n221) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U302 ( .A(i_acth[13]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n216) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U301 ( .A(i_acth[12]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n211) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U300 ( .A(i_acth[11]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n206) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U299 ( .A(i_acth[10]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n201) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U298 ( .A(i_acth[9]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n196) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U297 ( .A(i_acth[8]), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n191) );
  INV_X1 wrap_act_buffer_inst_act_buffer_inst_U296 ( .A(int_ifmaps_ptr[1]), 
        .ZN(wrap_act_buffer_inst_act_buffer_inst_n266) );
  NAND4_X1 wrap_act_buffer_inst_act_buffer_inst_U295 ( .A1(ctrl_ldh_v_n), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n265), .A3(
        wrap_act_buffer_inst_act_buffer_inst_n266), .A4(
        wrap_act_buffer_inst_act_buffer_inst_n267), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n145) );
  NAND4_X1 wrap_act_buffer_inst_act_buffer_inst_U294 ( .A1(int_ifmaps_ptr[2]), 
        .A2(ctrl_ldh_v_n), .A3(wrap_act_buffer_inst_act_buffer_inst_n265), 
        .A4(wrap_act_buffer_inst_act_buffer_inst_n266), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n149) );
  NAND4_X1 wrap_act_buffer_inst_act_buffer_inst_U293 ( .A1(int_ifmaps_ptr[1]), 
        .A2(ctrl_ldh_v_n), .A3(wrap_act_buffer_inst_act_buffer_inst_n265), 
        .A4(wrap_act_buffer_inst_act_buffer_inst_n267), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n147) );
  NAND4_X1 wrap_act_buffer_inst_act_buffer_inst_U292 ( .A1(int_ifmaps_ptr[2]), 
        .A2(int_ifmaps_ptr[0]), .A3(ctrl_ldh_v_n), .A4(
        wrap_act_buffer_inst_act_buffer_inst_n266), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n150) );
  NAND4_X1 wrap_act_buffer_inst_act_buffer_inst_U291 ( .A1(int_ifmaps_ptr[1]), 
        .A2(int_ifmaps_ptr[0]), .A3(ctrl_ldh_v_n), .A4(
        wrap_act_buffer_inst_act_buffer_inst_n267), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n148) );
  NAND4_X1 wrap_act_buffer_inst_act_buffer_inst_U290 ( .A1(int_ifmaps_ptr[0]), 
        .A2(ctrl_ldh_v_n), .A3(wrap_act_buffer_inst_act_buffer_inst_n266), 
        .A4(wrap_act_buffer_inst_act_buffer_inst_n267), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n146) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U289 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[20]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[4]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[12]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n135) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U288 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[44]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[28]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[36]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n1), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n134) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U287 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n134), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n135), .ZN(
        wrap_act_buffer_inst_int_i_data_if1[4]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U286 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[19]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[3]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[11]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n57) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U285 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[43]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[27]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[35]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n56) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U284 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n56), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n57), .ZN(
        wrap_act_buffer_inst_int_i_data_if6[3]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U283 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[19]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[3]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[11]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n41) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U282 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[43]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[27]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[35]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n40) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U281 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n40), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n41), .ZN(
        wrap_act_buffer_inst_int_i_data_if7[3]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U280 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[19]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[3]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[11]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n25) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U279 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[43]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[27]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[35]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n24) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U278 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n24), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n25), .ZN(
        wrap_act_buffer_inst_int_i_data_if8[3]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U277 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[21]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[5]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[13]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n69) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U276 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[45]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[29]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[37]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n68) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U275 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n68), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n69), .ZN(
        wrap_act_buffer_inst_int_i_data_if5[5]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U274 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[21]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[5]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[13]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n53) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U273 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[45]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[29]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[37]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n52) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U272 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n52), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n53), .ZN(
        wrap_act_buffer_inst_int_i_data_if6[5]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U264 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[21]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[5]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[13]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n37) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U263 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[45]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[29]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[37]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n36) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U262 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n36), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n37), .ZN(
        wrap_act_buffer_inst_int_i_data_if7[5]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U261 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[23]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[7]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[15]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n65) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U260 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[47]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[31]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[39]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n64) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U259 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n64), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n65), .ZN(
        wrap_act_buffer_inst_int_i_data_if5[7]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U258 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[23]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[7]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[15]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n49) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U257 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[47]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[31]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[39]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n48) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U256 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n48), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n49), .ZN(
        wrap_act_buffer_inst_int_i_data_if6[7]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U255 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[47]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n167), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[31]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n161), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[39]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n6), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n10) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U254 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[23]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n185), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[7]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n179), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[15]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n173), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n11) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U253 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n10), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n11), .ZN(
        wrap_act_buffer_inst_int_i_data_if8[7]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U252 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[23]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[7]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[15]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n33) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U251 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[47]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[31]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[39]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n32) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U250 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n32), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n33), .ZN(
        wrap_act_buffer_inst_int_i_data_if7[7]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U249 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[17]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[1]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[9]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n61) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U248 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[41]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[25]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[33]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n60) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U247 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n60), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n61), .ZN(
        wrap_act_buffer_inst_int_i_data_if6[1]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U246 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[17]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[1]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[9]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n45) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U245 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[41]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[25]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[33]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n44) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U244 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n44), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n45), .ZN(
        wrap_act_buffer_inst_int_i_data_if7[1]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U243 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[17]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[1]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[9]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n29) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U242 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[41]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[25]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[33]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n28) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U241 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n28), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n29), .ZN(
        wrap_act_buffer_inst_int_i_data_if8[1]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U240 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[18]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[2]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[10]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n59) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U239 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[42]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[26]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[34]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n58) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U238 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n58), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n59), .ZN(
        wrap_act_buffer_inst_int_i_data_if6[2]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U237 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[18]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[2]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[10]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n43) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U236 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[42]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[26]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[34]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n42) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U235 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n42), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n43), .ZN(
        wrap_act_buffer_inst_int_i_data_if7[2]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U234 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[18]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[2]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[10]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n27) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U233 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[42]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[26]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[34]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n26) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U232 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n26), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n27), .ZN(
        wrap_act_buffer_inst_int_i_data_if8[2]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U231 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[20]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[4]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[12]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n55) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U230 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[44]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[28]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[36]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n54) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U229 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n54), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n55), .ZN(
        wrap_act_buffer_inst_int_i_data_if6[4]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U228 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[20]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[4]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[12]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n71) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U227 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[44]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[28]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[36]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n70) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U226 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n70), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n71), .ZN(
        wrap_act_buffer_inst_int_i_data_if5[4]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U225 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[20]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[4]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[12]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n39) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U224 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[44]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[28]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[36]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n38) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U223 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n38), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n39), .ZN(
        wrap_act_buffer_inst_int_i_data_if7[4]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U222 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[22]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[6]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[14]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n67) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U221 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[46]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[30]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[38]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n66) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U220 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n66), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n67), .ZN(
        wrap_act_buffer_inst_int_i_data_if5[6]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U219 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[22]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[6]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[14]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n51) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U218 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[46]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[30]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[38]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n50) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U217 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n50), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n51), .ZN(
        wrap_act_buffer_inst_int_i_data_if6[6]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U216 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[46]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n167), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[30]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n161), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[38]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n6), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n18) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U215 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[22]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n185), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[6]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n179), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[14]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n173), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n19) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U214 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n18), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n19), .ZN(
        wrap_act_buffer_inst_int_i_data_if8[6]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U213 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[22]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[6]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[14]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n35) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U212 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[46]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[30]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[38]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n34) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U211 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n34), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n35), .ZN(
        wrap_act_buffer_inst_int_i_data_if7[6]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U210 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[16]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n183), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[0]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n177), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[8]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n171), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n63) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U209 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[40]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n165), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[24]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n159), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[32]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n4), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n62) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U208 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n62), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n63), .ZN(
        wrap_act_buffer_inst_int_i_data_if6[0]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U207 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[16]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[0]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[8]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n31) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U206 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[40]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[24]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[32]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n30) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U205 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n30), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n31), .ZN(
        wrap_act_buffer_inst_int_i_data_if8[0]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U204 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[16]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n184), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[0]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n178), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[8]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n172), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n47) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U203 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[40]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n166), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[24]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n160), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[32]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n5), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n46) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U202 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n46), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n47), .ZN(
        wrap_act_buffer_inst_int_i_data_if7[0]) );
  INV_X1 wrap_act_buffer_inst_act_buffer_inst_U201 ( .A(ps_int_ifmaps_ptr[1]), 
        .ZN(wrap_act_buffer_inst_act_buffer_inst_n187) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U200 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[43]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[27]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[35]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n1), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n136) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U199 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[19]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[3]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[11]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n137) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U198 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n136), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n137), .ZN(
        wrap_act_buffer_inst_int_i_data_if1[3]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U197 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[43]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[27]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[35]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n1), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n120) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U196 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[19]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[3]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[11]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n121) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U195 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n120), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n121), .ZN(
        wrap_act_buffer_inst_int_i_data_if2[3]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U194 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[45]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[29]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[37]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n1), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n132) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U193 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[21]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[5]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[13]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n133) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U192 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n132), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n133), .ZN(
        wrap_act_buffer_inst_int_i_data_if1[5]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U191 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[47]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[31]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[39]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n1), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n128) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U190 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[23]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[7]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[15]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n129) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U189 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n128), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n129), .ZN(
        wrap_act_buffer_inst_int_i_data_if1[7]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U188 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[41]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[25]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[33]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n1), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n140) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U187 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[17]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[1]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[9]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n141) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U186 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n140), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n141), .ZN(
        wrap_act_buffer_inst_int_i_data_if1[1]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U185 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[41]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[25]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[33]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n1), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n124) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U184 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[17]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[1]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[9]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n125) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U183 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n124), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n125), .ZN(
        wrap_act_buffer_inst_int_i_data_if2[1]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U182 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[42]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[26]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[34]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n1), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n138) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U181 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[18]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[2]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[10]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n139) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U180 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n138), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n139), .ZN(
        wrap_act_buffer_inst_int_i_data_if1[2]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U179 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[42]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[26]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[34]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n1), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n122) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U178 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[18]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[2]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[10]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n123) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U177 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n122), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n123), .ZN(
        wrap_act_buffer_inst_int_i_data_if2[2]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U176 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[46]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[30]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[38]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n1), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n130) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U175 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[22]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[6]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[14]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n131) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U174 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n130), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n131), .ZN(
        wrap_act_buffer_inst_int_i_data_if1[6]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U173 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[40]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[24]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[32]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n1), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n142) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U172 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[16]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[0]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[8]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n143) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U171 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n142), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n143), .ZN(
        wrap_act_buffer_inst_int_i_data_if1[0]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U170 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[40]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n162), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[24]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n7), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[32]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n1), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n126) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U169 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[16]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n180), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[0]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n174), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[8]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n168), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n127) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U168 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n126), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n127), .ZN(
        wrap_act_buffer_inst_int_i_data_if2[0]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U167 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[21]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n185), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[5]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n179), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[13]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n173), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n21) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U166 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[45]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n167), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[29]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n161), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[37]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n6), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n20) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U165 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n20), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n21), .ZN(
        wrap_act_buffer_inst_int_i_data_if8[5]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U164 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[20]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n185), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[4]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n179), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[12]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n173), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n23) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U163 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[44]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n167), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[28]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n161), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[36]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n6), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n22) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U162 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n22), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n23), .ZN(
        wrap_act_buffer_inst_int_i_data_if8[4]) );
  AND2_X1 wrap_act_buffer_inst_act_buffer_inst_U161 ( .A1(ps_int_ifmaps_ptr[2]), .A2(wrap_act_buffer_inst_act_buffer_inst_n186), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n14) );
  AND2_X1 wrap_act_buffer_inst_act_buffer_inst_U160 ( .A1(ps_int_ifmaps_ptr[2]), .A2(ps_int_ifmaps_ptr[0]), .ZN(wrap_act_buffer_inst_act_buffer_inst_n13) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U159 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n187), .A2(ps_int_ifmaps_ptr[0]), 
        .ZN(wrap_act_buffer_inst_act_buffer_inst_n16) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U158 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[19]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n182), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[3]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n176), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[11]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n170), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n73) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U157 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[43]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n164), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[27]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n9), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[35]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n3), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n72) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U156 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n72), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n73), .ZN(
        wrap_act_buffer_inst_int_i_data_if5[3]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U155 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[19]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[3]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[11]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n105) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U154 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[43]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[27]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[35]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n2), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n104) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U153 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n104), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n105), .ZN(
        wrap_act_buffer_inst_int_i_data_if3[3]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U152 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[19]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n182), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[3]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n176), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[11]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n170), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n89) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U151 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[43]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n164), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[27]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n9), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[35]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n3), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n88) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U150 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n88), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n89), .ZN(
        wrap_act_buffer_inst_int_i_data_if4[3]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U149 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[21]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[5]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[13]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n117) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U148 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[45]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[29]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[37]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n2), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n116) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U147 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n116), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n117), .ZN(
        wrap_act_buffer_inst_int_i_data_if2[5]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U146 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[21]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[5]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[13]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n101) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U145 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[45]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[29]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[37]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n2), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n100) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U144 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n100), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n101), .ZN(
        wrap_act_buffer_inst_int_i_data_if3[5]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U143 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[21]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n182), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[5]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n176), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[13]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n170), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n85) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U142 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[45]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n164), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[29]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n9), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[37]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n3), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n84) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U141 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n84), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n85), .ZN(
        wrap_act_buffer_inst_int_i_data_if4[5]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U140 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[23]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[7]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[15]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n113) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U139 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[47]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[31]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[39]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n2), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n112) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U138 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n112), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n113), .ZN(
        wrap_act_buffer_inst_int_i_data_if2[7]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U137 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[23]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[7]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[15]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n97) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U136 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[47]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[31]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[39]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n2), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n96) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U135 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n96), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n97), .ZN(
        wrap_act_buffer_inst_int_i_data_if3[7]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U134 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[23]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n182), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[7]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n176), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[15]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n170), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n81) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U133 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[47]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n164), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[31]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n9), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[39]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n3), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n80) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U132 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n80), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n81), .ZN(
        wrap_act_buffer_inst_int_i_data_if4[7]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U131 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[17]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n182), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[1]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n176), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[9]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n170), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n77) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U130 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[41]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n164), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[25]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n9), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[33]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n3), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n76) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U129 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n76), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n77), .ZN(
        wrap_act_buffer_inst_int_i_data_if5[1]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U128 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[17]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[1]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[9]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n109) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U127 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[41]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[25]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[33]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n2), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n108) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U126 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n108), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n109), .ZN(
        wrap_act_buffer_inst_int_i_data_if3[1]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U125 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[17]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n182), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[1]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n176), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[9]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n170), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n93) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U124 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[41]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n164), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[25]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n9), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[33]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n3), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n92) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U123 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n92), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n93), .ZN(
        wrap_act_buffer_inst_int_i_data_if4[1]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U122 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[18]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n182), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[2]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n176), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[10]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n170), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n75) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U121 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[42]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n164), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[26]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n9), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[34]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n3), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n74) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U120 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n74), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n75), .ZN(
        wrap_act_buffer_inst_int_i_data_if5[2]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U119 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[18]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[2]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[10]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n107) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U118 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[42]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[26]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[34]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n2), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n106) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U117 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n106), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n107), .ZN(
        wrap_act_buffer_inst_int_i_data_if3[2]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U116 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[18]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n182), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[2]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n176), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[10]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n170), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n91) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U115 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[42]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n164), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[26]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n9), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[34]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n3), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n90) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U114 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n90), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n91), .ZN(
        wrap_act_buffer_inst_int_i_data_if4[2]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U113 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[20]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[4]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[12]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n119) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U112 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[44]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[28]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[36]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n2), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n118) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U111 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n118), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n119), .ZN(
        wrap_act_buffer_inst_int_i_data_if2[4]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U110 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[20]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[4]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[12]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n103) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U109 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[44]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[28]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[36]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n2), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n102) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U108 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n102), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n103), .ZN(
        wrap_act_buffer_inst_int_i_data_if3[4]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U107 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[20]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n182), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[4]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n176), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[12]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n170), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n87) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U106 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[44]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n164), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[28]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n9), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[36]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n3), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n86) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U105 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n86), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n87), .ZN(
        wrap_act_buffer_inst_int_i_data_if4[4]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U104 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[22]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[6]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[14]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n115) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U103 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[46]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[30]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[38]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n2), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n114) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U102 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n114), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n115), .ZN(
        wrap_act_buffer_inst_int_i_data_if2[6]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U101 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[22]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[6]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[14]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n99) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U100 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[46]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[30]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[38]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n2), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n98) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U99 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n98), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n99), .ZN(
        wrap_act_buffer_inst_int_i_data_if3[6]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U98 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[22]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n182), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[6]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n176), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[14]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n170), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n83) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U97 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[46]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n164), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[30]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n9), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[38]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n3), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n82) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U96 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n82), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n83), .ZN(
        wrap_act_buffer_inst_int_i_data_if4[6]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U95 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[16]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n182), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[0]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n176), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[8]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n170), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n79) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U94 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[40]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n164), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[24]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n9), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[32]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n3), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n78) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U93 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n78), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n79), .ZN(
        wrap_act_buffer_inst_int_i_data_if5[0]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U92 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[16]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n182), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[0]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n176), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[8]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n170), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n95) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U91 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[40]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n164), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[24]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n9), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[32]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n3), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n94) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U90 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n94), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n95), .ZN(
        wrap_act_buffer_inst_int_i_data_if4[0]) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U89 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[16]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n181), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[0]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n175), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[8]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n169), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n111) );
  AOI222_X1 wrap_act_buffer_inst_act_buffer_inst_U88 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[40]), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n163), .B1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[24]), .B2(
        wrap_act_buffer_inst_act_buffer_inst_n8), .C1(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[32]), .C2(
        wrap_act_buffer_inst_act_buffer_inst_n2), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n110) );
  NAND2_X1 wrap_act_buffer_inst_act_buffer_inst_U87 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n110), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n111), .ZN(
        wrap_act_buffer_inst_int_i_data_if3[0]) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U86 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n145), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n157), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N120) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U85 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n149), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n151), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N152) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U84 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n145), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n151), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N156) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U83 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n149), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n152), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N146) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U82 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n145), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n152), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N150) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U81 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n149), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n153), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N140) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U80 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n145), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n153), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N144) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U79 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n149), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n154), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N134) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U78 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n145), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n154), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N138) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U77 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n149), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n155), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N128) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U76 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n145), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n155), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N132) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U75 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n149), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n156), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N122) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U74 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n145), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n156), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N126) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U73 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n149), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n157), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N116) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U72 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n147), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n151), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N154) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U71 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n147), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n152), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N148) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U70 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n147), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n153), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N142) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U69 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n147), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n154), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N136) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U68 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n147), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n155), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N130) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U67 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n147), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n156), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N124) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U66 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n147), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n157), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N118) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U65 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n150), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n151), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N151) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U64 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n148), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n151), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N153) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U63 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n150), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n152), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N145) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U62 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n148), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n152), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N147) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U61 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n150), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n153), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N139) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U60 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n148), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n153), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N141) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U59 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n150), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n154), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N133) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U58 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n148), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n154), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N135) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U57 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n150), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n155), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N127) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U56 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n148), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n155), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N129) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U55 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n150), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n156), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N121) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U54 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n148), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n156), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N123) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U53 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n150), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n157), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N115) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U52 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n148), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n157), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N117) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U51 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n146), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n151), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N155) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U50 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n146), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n152), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N149) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U49 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n146), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n153), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N143) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U48 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n146), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n154), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N137) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U47 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n146), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n155), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N131) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U46 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n146), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n156), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N125) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U45 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n146), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n157), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N119) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U44 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n144), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n150), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N157) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U43 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n144), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n149), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N158) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U42 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n144), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n148), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N159) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U41 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n144), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n147), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N160) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U40 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n144), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n146), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N161) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U39 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n144), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n145), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_N162) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U38 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n15), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n162) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U37 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n15), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n165) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U36 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n15), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n164) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U35 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n15), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n163) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U34 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n14), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n168) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U33 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n17), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n1) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U32 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n17), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n4) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U31 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n17), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n3) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U30 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n17), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n5) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U29 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n17), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n2) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U28 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n13), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n174) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U27 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n13), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n176) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U26 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n13), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n175) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U25 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n16), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n7) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U24 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n16), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n9) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U23 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n16), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n8) );
  NOR2_X1 wrap_act_buffer_inst_act_buffer_inst_U22 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n187), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n186), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n12) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U21 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n15), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n166) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U20 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n14), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n171) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U19 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n14), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n170) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U18 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n14), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n172) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U17 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n14), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n169) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U16 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n13), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n177) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U15 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n13), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n178) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U14 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n16), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n159) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U13 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n16), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n160) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U12 ( .A(n46), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n231) );
  AND4_X1 wrap_act_buffer_inst_act_buffer_inst_U11 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n144), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n151), .A3(
        wrap_act_buffer_inst_act_buffer_inst_n152), .A4(
        wrap_act_buffer_inst_act_buffer_inst_n153), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n158) );
  NAND4_X1 wrap_act_buffer_inst_act_buffer_inst_U10 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n155), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n154), .A3(
        wrap_act_buffer_inst_act_buffer_inst_n156), .A4(
        wrap_act_buffer_inst_act_buffer_inst_n158), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n157) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U9 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n12), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n180) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U8 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n12), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n183) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U7 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n12), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n182) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U6 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n12), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n184) );
  BUF_X1 wrap_act_buffer_inst_act_buffer_inst_U5 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n12), .Z(
        wrap_act_buffer_inst_act_buffer_inst_n181) );
  INV_X1 wrap_act_buffer_inst_act_buffer_inst_U4 ( .A(
        wrap_act_buffer_inst_act_buffer_inst_n231), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n264) );
  NOR3_X1 wrap_act_buffer_inst_act_buffer_inst_U3 ( .A1(ps_int_ifmaps_ptr[1]), 
        .A2(ps_int_ifmaps_ptr[2]), .A3(ps_int_ifmaps_ptr[0]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n15) );
  NOR3_X1 wrap_act_buffer_inst_act_buffer_inst_U2 ( .A1(ps_int_ifmaps_ptr[1]), 
        .A2(ps_int_ifmaps_ptr[2]), .A3(
        wrap_act_buffer_inst_act_buffer_inst_n186), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n17) );
  NAND3_X1 wrap_act_buffer_inst_act_buffer_inst_U271 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n188), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n190), .A3(int_npu_ptr[1]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n155) );
  NAND3_X1 wrap_act_buffer_inst_act_buffer_inst_U270 ( .A1(int_npu_ptr[0]), 
        .A2(wrap_act_buffer_inst_act_buffer_inst_n190), .A3(int_npu_ptr[1]), 
        .ZN(wrap_act_buffer_inst_act_buffer_inst_n154) );
  NAND3_X1 wrap_act_buffer_inst_act_buffer_inst_U269 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n189), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n190), .A3(int_npu_ptr[0]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n156) );
  NAND3_X1 wrap_act_buffer_inst_act_buffer_inst_U268 ( .A1(int_npu_ptr[1]), 
        .A2(int_npu_ptr[0]), .A3(int_npu_ptr[2]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n144) );
  NAND3_X1 wrap_act_buffer_inst_act_buffer_inst_U267 ( .A1(int_npu_ptr[1]), 
        .A2(wrap_act_buffer_inst_act_buffer_inst_n188), .A3(int_npu_ptr[2]), 
        .ZN(wrap_act_buffer_inst_act_buffer_inst_n151) );
  NAND3_X1 wrap_act_buffer_inst_act_buffer_inst_U266 ( .A1(int_npu_ptr[0]), 
        .A2(wrap_act_buffer_inst_act_buffer_inst_n189), .A3(int_npu_ptr[2]), 
        .ZN(wrap_act_buffer_inst_act_buffer_inst_n152) );
  NAND3_X1 wrap_act_buffer_inst_act_buffer_inst_U265 ( .A1(
        wrap_act_buffer_inst_act_buffer_inst_n188), .A2(
        wrap_act_buffer_inst_act_buffer_inst_n189), .A3(int_npu_ptr[2]), .ZN(
        wrap_act_buffer_inst_act_buffer_inst_n153) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_5__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n191), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4755), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n232), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[0]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_5__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n196), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4755), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n232), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[1]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_5__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n201), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4755), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n232), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[2]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_5__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n206), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4755), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n232), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[3]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_5__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n211), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4755), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n232), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[4]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_5__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n216), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4755), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n232), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[5]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_5__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n221), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4755), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n232), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[6]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_5__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n226), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4755), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n232), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[7]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_4__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n191), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4750), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n232), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[8]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_4__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n196), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4750), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n232), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[9]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_4__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n201), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4750), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n232), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[10]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_4__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n206), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4750), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n232), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[11]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_4__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n211), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4750), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n233), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[12]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_4__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n216), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4750), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n233), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[13]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_4__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n221), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4750), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n233), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[14]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_4__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n226), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4750), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n233), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[15]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_3__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n191), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4745), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n233), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[16]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_3__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n196), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4745), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n233), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[17]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_3__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n201), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4745), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n233), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[18]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_3__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n206), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4745), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n233), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[19]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_3__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n211), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4745), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n233), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[20]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_3__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n216), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4745), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n233), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[21]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_3__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n221), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4745), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n233), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[22]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_3__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n226), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4745), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n233), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[23]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_2__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n191), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4740), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n234), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[24]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_2__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n196), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4740), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n234), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[25]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_2__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n201), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4740), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n234), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[26]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_2__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n206), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4740), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n234), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[27]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_2__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n211), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4740), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n234), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[28]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_2__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n216), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4740), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n234), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[29]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_2__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n221), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4740), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n234), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[30]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_2__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n226), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4740), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n234), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[31]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_1__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n191), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4735), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n234), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[32]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_1__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n196), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4735), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n234), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[33]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_1__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n201), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4735), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n234), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[34]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_1__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n206), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4735), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n234), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[35]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_1__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n211), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4735), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n235), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[36]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_1__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n216), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4735), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n235), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[37]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_1__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n221), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4735), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n235), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[38]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_1__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n226), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4735), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n235), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[39]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_0__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n191), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4730), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n235), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[40]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_0__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n196), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4730), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n235), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[41]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_0__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n201), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4730), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n235), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[42]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_0__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n206), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4730), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n235), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[43]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_0__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n211), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4730), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n235), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[44]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_0__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n216), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4730), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n235), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[45]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_0__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n221), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4730), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n235), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[46]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data8_reg_0__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n226), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4730), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n235), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data8[47]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_5__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n191), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4725), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n236), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[0]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_5__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n196), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4725), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n236), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[1]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_5__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n201), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4725), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n236), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[2]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_5__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n206), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4725), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n236), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[3]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_5__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n211), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4725), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n236), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[4]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_5__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n216), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4725), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n236), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[5]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_5__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n221), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4725), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n236), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[6]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_5__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n226), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4725), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n236), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[7]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_4__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n191), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4720), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n236), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[8]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_4__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n196), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4720), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n236), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[9]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_4__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n201), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4720), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n236), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[10]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_4__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n206), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4720), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n236), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[11]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_4__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n211), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4720), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n237), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[12]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_4__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n216), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4720), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n237), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[13]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_4__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n221), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4720), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n237), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[14]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_4__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n226), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4720), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n237), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[15]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_3__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n191), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4715), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n237), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[16]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_3__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n196), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4715), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n237), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[17]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_3__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n201), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4715), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n237), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[18]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_3__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n206), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4715), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n237), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[19]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_3__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n211), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4715), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n237), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[20]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_3__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n216), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4715), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n237), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[21]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_3__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n221), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4715), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n237), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[22]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_3__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n226), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4715), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n237), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[23]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_2__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n191), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4710), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n238), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[24]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_2__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n196), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4710), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n238), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[25]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_2__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n201), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4710), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n238), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[26]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_2__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n206), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4710), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n238), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[27]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_2__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n211), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4710), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n238), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[28]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_2__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n216), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4710), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n238), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[29]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_2__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n221), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4710), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n238), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[30]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_2__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n226), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4710), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n238), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[31]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_1__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n191), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4705), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n238), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[32]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_1__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n196), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4705), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n238), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[33]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_1__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n201), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4705), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n238), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[34]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_1__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n206), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4705), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n238), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[35]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_1__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n211), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4705), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n239), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[36]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_1__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n216), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4705), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n239), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[37]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_1__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n221), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4705), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n239), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[38]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_1__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n226), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4705), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n239), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[39]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_0__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n192), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4700), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n239), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[40]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_0__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n197), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4700), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n239), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[41]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_0__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n202), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4700), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n239), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[42]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_0__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n207), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4700), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n239), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[43]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_0__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n212), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4700), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n239), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[44]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_0__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n217), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4700), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n239), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[45]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_0__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n222), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4700), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n239), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[46]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data7_reg_0__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n227), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4700), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n239), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data7[47]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_5__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n192), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4695), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n240), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[0]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_5__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n197), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4695), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n240), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[1]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_5__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n202), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4695), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n240), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[2]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_5__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n207), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4695), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n240), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[3]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_5__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n212), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4695), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n240), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[4]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_5__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n217), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4695), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n240), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[5]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_5__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n222), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4695), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n240), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[6]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_5__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n227), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4695), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n240), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[7]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_4__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n192), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4690), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n240), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[8]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_4__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n197), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4690), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n240), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[9]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_4__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n202), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4690), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n240), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[10]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_4__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n207), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4690), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n240), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[11]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_4__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n212), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4690), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n241), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[12]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_4__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n217), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4690), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n241), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[13]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_4__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n222), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4690), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n241), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[14]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_4__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n227), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4690), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n241), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[15]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_3__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n192), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4685), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n241), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[16]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_3__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n197), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4685), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n241), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[17]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_3__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n202), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4685), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n241), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[18]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_3__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n207), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4685), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n241), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[19]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_3__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n212), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4685), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n241), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[20]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_3__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n217), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4685), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n241), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[21]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_3__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n222), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4685), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n241), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[22]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_3__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n227), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4685), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n241), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[23]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_2__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n192), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4680), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n242), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[24]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_2__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n197), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4680), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n242), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[25]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_2__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n202), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4680), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n242), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[26]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_2__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n207), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4680), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n242), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[27]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_2__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n212), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4680), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n242), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[28]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_2__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n217), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4680), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n242), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[29]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_2__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n222), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4680), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n242), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[30]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_2__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n227), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4680), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n242), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[31]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_1__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n192), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4675), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n242), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[32]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_1__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n197), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4675), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n242), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[33]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_1__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n202), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4675), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n242), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[34]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_1__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n207), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4675), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n242), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[35]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_1__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n212), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4675), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n243), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[36]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_1__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n217), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4675), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n243), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[37]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_1__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n222), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4675), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n243), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[38]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_1__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n227), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4675), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n243), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[39]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_0__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n192), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4670), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n243), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[40]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_0__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n197), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4670), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n243), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[41]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_0__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n202), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4670), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n243), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[42]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_0__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n207), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4670), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n243), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[43]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_0__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n212), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4670), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n243), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[44]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_0__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n217), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4670), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n243), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[45]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_0__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n222), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4670), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n243), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[46]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data6_reg_0__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n227), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4670), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n243), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data6[47]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_5__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n192), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4665), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n244), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[0]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_5__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n197), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4665), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n244), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[1]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_5__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n202), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4665), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n244), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[2]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_5__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n207), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4665), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n244), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[3]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_5__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n212), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4665), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n244), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[4]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_5__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n217), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4665), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n244), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[5]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_5__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n222), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4665), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n244), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[6]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_5__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n227), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4665), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n244), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[7]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_4__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n192), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4660), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n244), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[8]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_4__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n197), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4660), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n244), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[9]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_4__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n202), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4660), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n244), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[10]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_4__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n207), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4660), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n244), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[11]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_4__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n212), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4660), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n245), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[12]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_4__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n217), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4660), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n245), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[13]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_4__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n222), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4660), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n245), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[14]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_4__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n227), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4660), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n245), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[15]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_3__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n192), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4655), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n245), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[16]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_3__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n197), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4655), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n245), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[17]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_3__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n202), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4655), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n245), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[18]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_3__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n207), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4655), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n245), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[19]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_3__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n212), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4655), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n245), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[20]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_3__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n217), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4655), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n245), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[21]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_3__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n222), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4655), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n245), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[22]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_3__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n227), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4655), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n245), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[23]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_2__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n192), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4650), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n246), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[24]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_2__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n197), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4650), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n246), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[25]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_2__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n202), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4650), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n246), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[26]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_2__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n207), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4650), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n246), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[27]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_2__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n212), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4650), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n246), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[28]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_2__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n217), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4650), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n246), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[29]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_2__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n222), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4650), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n246), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[30]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_2__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n227), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4650), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n246), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[31]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_1__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n193), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4645), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n246), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[32]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_1__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n198), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4645), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n246), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[33]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_1__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n203), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4645), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n246), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[34]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_1__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n208), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4645), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n246), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[35]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_1__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n213), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4645), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n247), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[36]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_1__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n218), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4645), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n247), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[37]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_1__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n223), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4645), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n247), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[38]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_1__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n228), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4645), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n247), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[39]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_0__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n193), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4640), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n247), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[40]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_0__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n198), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4640), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n247), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[41]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_0__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n203), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4640), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n247), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[42]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_0__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n208), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4640), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n247), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[43]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_0__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n213), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4640), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n247), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[44]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_0__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n218), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4640), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n247), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[45]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_0__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n223), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4640), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n247), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[46]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data5_reg_0__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n228), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4640), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n247), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data5[47]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_5__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n193), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4635), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n248), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[0]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_5__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n198), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4635), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n248), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[1]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_5__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n203), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4635), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n248), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[2]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_5__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n208), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4635), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n248), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[3]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_5__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n213), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4635), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n248), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[4]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_5__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n218), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4635), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n248), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[5]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_5__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n223), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4635), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n248), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[6]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_5__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n228), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4635), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n248), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[7]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_4__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n193), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4630), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n248), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[8]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_4__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n198), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4630), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n248), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[9]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_4__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n203), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4630), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n248), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[10]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_4__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n208), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4630), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n248), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[11]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_4__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n213), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4630), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n249), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[12]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_4__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n218), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4630), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n249), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[13]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_4__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n223), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4630), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n249), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[14]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_4__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n228), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4630), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n249), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[15]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_3__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n193), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4625), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n249), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[16]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_3__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n198), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4625), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n249), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[17]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_3__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n203), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4625), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n249), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[18]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_3__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n208), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4625), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n249), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[19]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_3__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n213), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4625), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n249), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[20]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_3__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n218), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4625), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n249), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[21]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_3__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n223), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4625), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n249), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[22]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_3__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n228), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4625), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n249), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[23]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_2__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n193), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4620), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n250), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[24]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_2__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n198), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4620), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n250), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[25]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_2__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n203), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4620), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n250), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[26]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_2__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n208), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4620), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n250), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[27]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_2__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n213), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4620), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n250), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[28]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_2__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n218), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4620), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n250), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[29]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_2__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n223), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4620), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n250), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[30]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_2__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n228), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4620), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n250), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[31]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_1__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n193), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4615), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n250), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[32]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_1__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n198), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4615), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n250), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[33]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_1__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n203), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4615), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n250), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[34]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_1__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n208), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4615), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n250), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[35]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_1__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n213), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4615), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n251), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[36]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_1__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n218), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4615), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n251), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[37]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_1__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n223), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4615), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n251), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[38]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_1__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n228), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4615), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n251), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[39]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_0__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n193), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4610), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n251), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[40]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_0__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n198), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4610), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n251), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[41]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_0__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n203), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4610), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n251), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[42]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_0__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n208), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4610), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n251), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[43]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_0__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n213), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4610), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n251), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[44]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_0__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n218), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4610), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n251), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[45]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_0__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n223), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4610), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n251), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[46]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data4_reg_0__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n228), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4610), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n251), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data4[47]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_5__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n193), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4605), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n252), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[0]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_5__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n198), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4605), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n252), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[1]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_5__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n203), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4605), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n252), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[2]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_5__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n208), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4605), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n252), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[3]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_5__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n213), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4605), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n252), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[4]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_5__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n218), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4605), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n252), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[5]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_5__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n223), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4605), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n252), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[6]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_5__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n228), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4605), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n252), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[7]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_4__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n193), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4600), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n252), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[8]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_4__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n198), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4600), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n252), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[9]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_4__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n203), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4600), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n252), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[10]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_4__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n208), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4600), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n252), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[11]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_4__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n213), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4600), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n253), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[12]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_4__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n218), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4600), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n253), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[13]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_4__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n223), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4600), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n253), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[14]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_4__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n228), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4600), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n253), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[15]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_3__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n193), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4595), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n253), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[16]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_3__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n198), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4595), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n253), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[17]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_3__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n203), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4595), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n253), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[18]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_3__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n208), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4595), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n253), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[19]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_3__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n213), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4595), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n253), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[20]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_3__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n218), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4595), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n253), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[21]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_3__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n223), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4595), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n253), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[22]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_3__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n228), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4595), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n253), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[23]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_2__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n194), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4590), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n254), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[24]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_2__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n199), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4590), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n254), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[25]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_2__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n204), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4590), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n254), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[26]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_2__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n209), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4590), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n254), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[27]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_2__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n214), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4590), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n254), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[28]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_2__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n219), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4590), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n254), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[29]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_2__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n224), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4590), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n254), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[30]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_2__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n229), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4590), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n254), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[31]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_1__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n194), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4585), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n254), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[32]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_1__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n199), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4585), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n254), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[33]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_1__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n204), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4585), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n254), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[34]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_1__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n209), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4585), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n254), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[35]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_1__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n214), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4585), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n255), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[36]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_1__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n219), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4585), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n255), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[37]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_1__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n224), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4585), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n255), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[38]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_1__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n229), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4585), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n255), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[39]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_0__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n194), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4580), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n255), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[40]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_0__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n199), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4580), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n255), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[41]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_0__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n204), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4580), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n255), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[42]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_0__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n209), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4580), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n255), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[43]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_0__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n214), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4580), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n255), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[44]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_0__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n219), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4580), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n255), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[45]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_0__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n224), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4580), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n255), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[46]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data3_reg_0__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n229), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4580), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n255), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data3[47]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_5__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n194), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4575), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n256), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[0]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_5__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n199), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4575), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n256), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[1]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_5__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n204), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4575), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n256), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[2]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_5__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n209), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4575), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n256), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[3]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_5__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n214), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4575), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n256), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[4]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_5__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n219), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4575), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n256), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[5]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_5__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n224), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4575), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n256), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[6]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_5__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n229), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4575), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n256), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[7]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_4__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n194), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4570), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n256), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[8]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_4__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n199), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4570), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n256), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[9]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_4__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n204), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4570), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n256), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[10]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_4__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n209), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4570), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n256), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[11]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_4__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n214), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4570), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n257), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[12]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_4__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n219), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4570), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n257), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[13]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_4__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n224), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4570), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n257), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[14]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_4__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n229), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4570), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n257), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[15]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_3__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n194), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4565), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n257), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[16]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_3__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n199), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4565), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n257), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[17]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_3__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n204), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4565), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n257), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[18]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_3__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n209), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4565), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n257), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[19]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_3__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n214), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4565), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n257), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[20]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_3__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n219), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4565), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n257), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[21]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_3__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n224), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4565), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n257), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[22]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_3__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n229), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4565), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n257), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[23]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_2__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n194), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4560), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n258), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[24]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_2__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n199), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4560), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n258), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[25]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_2__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n204), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4560), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n258), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[26]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_2__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n209), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4560), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n258), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[27]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_2__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n214), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4560), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n258), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[28]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_2__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n219), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4560), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n258), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[29]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_2__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n224), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4560), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n258), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[30]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_2__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n229), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4560), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n258), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[31]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_1__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n194), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4555), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n258), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[32]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_1__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n199), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4555), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n258), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[33]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_1__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n204), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4555), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n258), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[34]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_1__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n209), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4555), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n258), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[35]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_1__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n214), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4555), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n259), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[36]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_1__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n219), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4555), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n259), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[37]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_1__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n224), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4555), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n259), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[38]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_1__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n229), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4555), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n259), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[39]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_0__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n194), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4550), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n259), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[40]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_0__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n199), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4550), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n259), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[41]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_0__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n204), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4550), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n259), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[42]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_0__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n209), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4550), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n259), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[43]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_0__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n214), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4550), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n259), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[44]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_0__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n219), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4550), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n259), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[45]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_0__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n224), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4550), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n259), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[46]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data2_reg_0__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n229), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4550), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n259), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data2[47]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_5__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n194), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4545), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n260), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[0]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_5__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n199), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4545), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n260), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[1]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_5__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n204), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4545), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n260), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[2]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_5__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n209), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4545), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n260), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[3]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_5__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n214), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4545), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n260), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[4]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_5__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n219), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4545), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n260), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[5]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_5__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n224), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4545), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n260), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[6]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_5__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n229), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4545), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n260), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[7]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_4__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n194), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4540), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n260), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[8]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_4__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n199), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4540), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n260), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[9]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_4__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n204), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4540), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n260), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[10]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_4__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n209), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4540), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n260), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[11]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_4__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n214), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4540), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n261), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[12]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_4__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n219), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4540), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n261), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[13]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_4__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n224), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4540), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n261), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[14]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_4__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n229), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4540), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n261), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[15]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_3__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n195), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4535), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n261), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[16]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_3__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n200), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4535), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n261), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[17]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_3__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n205), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4535), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n261), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[18]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_3__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n210), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4535), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n261), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[19]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_3__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n215), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4535), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n261), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[20]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_3__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n220), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4535), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n261), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[21]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_3__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n225), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4535), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n261), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[22]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_3__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n230), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4535), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n261), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[23]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_2__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n195), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4530), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n262), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[24]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_2__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n200), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4530), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n262), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[25]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_2__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n205), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4530), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n262), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[26]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_2__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n210), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4530), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n262), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[27]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_2__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n215), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4530), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n262), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[28]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_2__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n220), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4530), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n262), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[29]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_2__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n225), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4530), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n262), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[30]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_2__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n230), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4530), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n262), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[31]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_1__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n195), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4525), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n262), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[32]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_1__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n200), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4525), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n262), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[33]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_1__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n205), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4525), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n262), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[34]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_1__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n210), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4525), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n262), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[35]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_1__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n215), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4525), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n263), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[36]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_1__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n220), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4525), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n263), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[37]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_1__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n225), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4525), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n263), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[38]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_1__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n230), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4525), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n263), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[39]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_0__0_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n195), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4519), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n263), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[40]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_0__1_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n200), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4519), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n263), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[41]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_0__2_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n205), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4519), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n263), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[42]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_0__3_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n210), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4519), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n263), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[43]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_0__4_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n215), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4519), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n263), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[44]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_0__5_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n220), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4519), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n263), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[45]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_0__6_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n225), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4519), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n263), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[46]) );
  DFFR_X1 wrap_act_buffer_inst_act_buffer_inst_int_data1_reg_0__7_ ( .D(
        wrap_act_buffer_inst_act_buffer_inst_n230), .CK(
        wrap_act_buffer_inst_act_buffer_inst_net4519), .RN(
        wrap_act_buffer_inst_act_buffer_inst_n263), .Q(
        wrap_act_buffer_inst_act_buffer_inst_int_data1[47]) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data1_reg_0__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N120), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4519) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data1_reg_1__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N119), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4525) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data1_reg_2__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N118), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4530) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data1_reg_3__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N117), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4535) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data1_reg_4__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N116), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4540) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data1_reg_5__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N115), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4545) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data2_reg_0__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N126), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4550) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data2_reg_1__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N125), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4555) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data2_reg_2__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N124), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4560) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data2_reg_3__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N123), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4565) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data2_reg_4__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N122), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4570) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data2_reg_5__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N121), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4575) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data3_reg_0__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N132), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4580) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data3_reg_1__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N131), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4585) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data3_reg_2__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N130), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4590) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data3_reg_3__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N129), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4595) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data3_reg_4__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N128), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4600) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data3_reg_5__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N127), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4605) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data4_reg_0__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N138), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4610) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data4_reg_1__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N137), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4615) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data4_reg_2__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N136), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4620) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data4_reg_3__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N135), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4625) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data4_reg_4__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N134), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4630) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data4_reg_5__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N133), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4635) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data5_reg_0__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N144), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4640) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data5_reg_1__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N143), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4645) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data5_reg_2__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N142), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4650) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data5_reg_3__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N141), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4655) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data5_reg_4__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N140), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4660) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data5_reg_5__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N139), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4665) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data6_reg_0__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N150), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4670) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data6_reg_1__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N149), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4675) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data6_reg_2__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N148), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4680) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data6_reg_3__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N147), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4685) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data6_reg_4__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N146), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4690) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data6_reg_5__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N145), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4695) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data7_reg_0__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N156), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4700) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data7_reg_1__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N155), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4705) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data7_reg_2__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N154), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4710) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data7_reg_3__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N153), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4715) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data7_reg_4__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N152), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4720) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data7_reg_5__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N151), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4725) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data8_reg_0__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N162), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4730) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data8_reg_1__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N161), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4735) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data8_reg_2__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N160), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4740) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data8_reg_3__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N159), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4745) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data8_reg_4__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N158), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4750) );
  CLKGATETST_X1 wrap_act_buffer_inst_act_buffer_inst_clk_gate_int_data8_reg_5__latch ( 
        .CK(ck), .E(wrap_act_buffer_inst_act_buffer_inst_N157), .SE(1'b0), 
        .GCK(wrap_act_buffer_inst_act_buffer_inst_net4755) );
  NOR3_X4 wrap_act_buffer_inst_act_if_inst_U392 ( .A1(ps_int_hmode_cnt[0]), 
        .A2(1'b0), .A3(wrap_act_buffer_inst_act_if_inst_n312), .ZN(
        wrap_act_buffer_inst_act_if_inst_n7) );
  CLKBUF_X1 wrap_act_buffer_inst_act_if_inst_U391 ( .A(int_npu_ptr[0]), .Z(
        wrap_act_buffer_inst_act_if_inst_n305) );
  CLKBUF_X1 wrap_act_buffer_inst_act_if_inst_U390 ( .A(int_npu_ptr[1]), .Z(
        wrap_act_buffer_inst_act_if_inst_n299) );
  CLKBUF_X1 wrap_act_buffer_inst_act_if_inst_U389 ( .A(int_npu_ptr[2]), .Z(
        wrap_act_buffer_inst_act_if_inst_n293) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U388 ( .A(
        wrap_act_buffer_inst_act_if_inst_n130), .B(
        wrap_act_buffer_inst_act_if_inst_n131), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n164) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U387 ( .A(
        wrap_act_buffer_inst_act_if_inst_n124), .B(
        wrap_act_buffer_inst_act_if_inst_n125), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n163) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U386 ( .A(
        wrap_act_buffer_inst_act_if_inst_n118), .B(
        wrap_act_buffer_inst_act_if_inst_n119), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n162) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U385 ( .A(
        wrap_act_buffer_inst_act_if_inst_n112), .B(
        wrap_act_buffer_inst_act_if_inst_n113), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n161) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U384 ( .A(
        wrap_act_buffer_inst_act_if_inst_n106), .B(
        wrap_act_buffer_inst_act_if_inst_n107), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n160) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U383 ( .A(
        wrap_act_buffer_inst_act_if_inst_n100), .B(
        wrap_act_buffer_inst_act_if_inst_n101), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n159) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U382 ( .A(
        wrap_act_buffer_inst_act_if_inst_n94), .B(
        wrap_act_buffer_inst_act_if_inst_n95), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n158) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U381 ( .A(
        wrap_act_buffer_inst_act_if_inst_n88), .B(
        wrap_act_buffer_inst_act_if_inst_n89), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n157) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U380 ( .A(
        wrap_act_buffer_inst_act_if_inst_n82), .B(
        wrap_act_buffer_inst_act_if_inst_n83), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n156) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U379 ( .A(
        wrap_act_buffer_inst_act_if_inst_n76), .B(
        wrap_act_buffer_inst_act_if_inst_n77), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n155) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U378 ( .A(
        wrap_act_buffer_inst_act_if_inst_n70), .B(
        wrap_act_buffer_inst_act_if_inst_n71), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n154) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U377 ( .A(
        wrap_act_buffer_inst_act_if_inst_n64), .B(
        wrap_act_buffer_inst_act_if_inst_n65), .S(
        wrap_act_buffer_inst_act_if_inst_n298), .Z(
        wrap_act_buffer_inst_act_if_inst_n153) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U376 ( .A(
        wrap_act_buffer_inst_act_if_inst_n58), .B(
        wrap_act_buffer_inst_act_if_inst_n59), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n152) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U375 ( .A(
        wrap_act_buffer_inst_act_if_inst_n52), .B(
        wrap_act_buffer_inst_act_if_inst_n53), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n151) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U374 ( .A(
        wrap_act_buffer_inst_act_if_inst_n46), .B(
        wrap_act_buffer_inst_act_if_inst_n47), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n150) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U373 ( .A(
        wrap_act_buffer_inst_act_if_inst_n40), .B(
        wrap_act_buffer_inst_act_if_inst_n41), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n149) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U372 ( .A(
        wrap_act_buffer_inst_act_if_inst_n127), .B(
        wrap_act_buffer_inst_act_if_inst_n128), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n148) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U371 ( .A(
        wrap_act_buffer_inst_act_if_inst_n121), .B(
        wrap_act_buffer_inst_act_if_inst_n122), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n147) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U370 ( .A(
        wrap_act_buffer_inst_act_if_inst_n115), .B(
        wrap_act_buffer_inst_act_if_inst_n116), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n146) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U369 ( .A(
        wrap_act_buffer_inst_act_if_inst_n109), .B(
        wrap_act_buffer_inst_act_if_inst_n110), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n145) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U368 ( .A(
        wrap_act_buffer_inst_act_if_inst_n103), .B(
        wrap_act_buffer_inst_act_if_inst_n104), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n144) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U367 ( .A(
        wrap_act_buffer_inst_act_if_inst_n97), .B(
        wrap_act_buffer_inst_act_if_inst_n98), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n143) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U366 ( .A(
        wrap_act_buffer_inst_act_if_inst_n91), .B(
        wrap_act_buffer_inst_act_if_inst_n92), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n142) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U365 ( .A(
        wrap_act_buffer_inst_act_if_inst_n85), .B(
        wrap_act_buffer_inst_act_if_inst_n86), .S(
        wrap_act_buffer_inst_act_if_inst_n297), .Z(
        wrap_act_buffer_inst_act_if_inst_n141) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U364 ( .A(
        wrap_act_buffer_inst_act_if_inst_n79), .B(
        wrap_act_buffer_inst_act_if_inst_n80), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n140) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U363 ( .A(
        wrap_act_buffer_inst_act_if_inst_n73), .B(
        wrap_act_buffer_inst_act_if_inst_n74), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n139) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U362 ( .A(
        wrap_act_buffer_inst_act_if_inst_n67), .B(
        wrap_act_buffer_inst_act_if_inst_n68), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n138) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U361 ( .A(
        wrap_act_buffer_inst_act_if_inst_n61), .B(
        wrap_act_buffer_inst_act_if_inst_n62), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n137) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U360 ( .A(
        wrap_act_buffer_inst_act_if_inst_n55), .B(
        wrap_act_buffer_inst_act_if_inst_n56), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n136) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U359 ( .A(
        wrap_act_buffer_inst_act_if_inst_n49), .B(
        wrap_act_buffer_inst_act_if_inst_n50), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n135) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U358 ( .A(
        wrap_act_buffer_inst_act_if_inst_n43), .B(
        wrap_act_buffer_inst_act_if_inst_n44), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n134) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U357 ( .A(
        wrap_act_buffer_inst_act_if_inst_n1), .B(
        wrap_act_buffer_inst_act_if_inst_n2), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n133) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U356 ( .A(
        wrap_act_buffer_inst_act_if_inst_n131), .B(
        wrap_act_buffer_inst_act_if_inst_n130), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n132) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U355 ( .A(
        wrap_act_buffer_inst_act_if_inst_n180), .B(
        wrap_act_buffer_inst_act_if_inst_n172), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n131) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U354 ( .A(
        wrap_act_buffer_inst_act_if_inst_n226), .B(
        wrap_act_buffer_inst_act_if_inst_n204), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n130) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U353 ( .A(
        wrap_act_buffer_inst_act_if_inst_n128), .B(
        wrap_act_buffer_inst_act_if_inst_n127), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n129) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U352 ( .A(
        wrap_act_buffer_inst_act_if_inst_n288), .B(
        wrap_act_buffer_inst_act_if_inst_n250), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n128) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U351 ( .A(
        wrap_act_buffer_inst_act_if_inst_n196), .B(
        wrap_act_buffer_inst_act_if_inst_n188), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n127) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U350 ( .A(
        wrap_act_buffer_inst_act_if_inst_n125), .B(
        wrap_act_buffer_inst_act_if_inst_n124), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n126) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U349 ( .A(
        wrap_act_buffer_inst_act_if_inst_n179), .B(
        wrap_act_buffer_inst_act_if_inst_n171), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n125) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U348 ( .A(
        wrap_act_buffer_inst_act_if_inst_n223), .B(
        wrap_act_buffer_inst_act_if_inst_n203), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n124) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U347 ( .A(
        wrap_act_buffer_inst_act_if_inst_n122), .B(
        wrap_act_buffer_inst_act_if_inst_n121), .S(
        wrap_act_buffer_inst_act_if_inst_n296), .Z(
        wrap_act_buffer_inst_act_if_inst_n123) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U346 ( .A(
        wrap_act_buffer_inst_act_if_inst_n283), .B(
        wrap_act_buffer_inst_act_if_inst_n247), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n122) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U345 ( .A(
        wrap_act_buffer_inst_act_if_inst_n195), .B(
        wrap_act_buffer_inst_act_if_inst_n187), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n121) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U344 ( .A(
        wrap_act_buffer_inst_act_if_inst_n119), .B(
        wrap_act_buffer_inst_act_if_inst_n118), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n120) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U343 ( .A(
        wrap_act_buffer_inst_act_if_inst_n178), .B(
        wrap_act_buffer_inst_act_if_inst_n170), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n119) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U342 ( .A(
        wrap_act_buffer_inst_act_if_inst_n220), .B(
        wrap_act_buffer_inst_act_if_inst_n202), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n118) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U341 ( .A(
        wrap_act_buffer_inst_act_if_inst_n116), .B(
        wrap_act_buffer_inst_act_if_inst_n115), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n117) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U340 ( .A(
        wrap_act_buffer_inst_act_if_inst_n278), .B(
        wrap_act_buffer_inst_act_if_inst_n244), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n116) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U339 ( .A(
        wrap_act_buffer_inst_act_if_inst_n194), .B(
        wrap_act_buffer_inst_act_if_inst_n186), .S(
        wrap_act_buffer_inst_act_if_inst_n310), .Z(
        wrap_act_buffer_inst_act_if_inst_n115) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U338 ( .A(
        wrap_act_buffer_inst_act_if_inst_n113), .B(
        wrap_act_buffer_inst_act_if_inst_n112), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n114) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U337 ( .A(
        wrap_act_buffer_inst_act_if_inst_n177), .B(
        wrap_act_buffer_inst_act_if_inst_n169), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n113) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U336 ( .A(
        wrap_act_buffer_inst_act_if_inst_n217), .B(
        wrap_act_buffer_inst_act_if_inst_n201), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n112) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U335 ( .A(
        wrap_act_buffer_inst_act_if_inst_n110), .B(
        wrap_act_buffer_inst_act_if_inst_n109), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n111) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U334 ( .A(
        wrap_act_buffer_inst_act_if_inst_n273), .B(
        wrap_act_buffer_inst_act_if_inst_n241), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n110) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U333 ( .A(
        wrap_act_buffer_inst_act_if_inst_n193), .B(
        wrap_act_buffer_inst_act_if_inst_n185), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n109) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U332 ( .A(
        wrap_act_buffer_inst_act_if_inst_n107), .B(
        wrap_act_buffer_inst_act_if_inst_n106), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n108) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U331 ( .A(
        wrap_act_buffer_inst_act_if_inst_n176), .B(
        wrap_act_buffer_inst_act_if_inst_n168), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n107) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U330 ( .A(
        wrap_act_buffer_inst_act_if_inst_n214), .B(
        wrap_act_buffer_inst_act_if_inst_n200), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n106) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U329 ( .A(
        wrap_act_buffer_inst_act_if_inst_n104), .B(
        wrap_act_buffer_inst_act_if_inst_n103), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n105) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U328 ( .A(
        wrap_act_buffer_inst_act_if_inst_n268), .B(
        wrap_act_buffer_inst_act_if_inst_n238), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n104) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U327 ( .A(
        wrap_act_buffer_inst_act_if_inst_n192), .B(
        wrap_act_buffer_inst_act_if_inst_n184), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n103) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U326 ( .A(
        wrap_act_buffer_inst_act_if_inst_n101), .B(
        wrap_act_buffer_inst_act_if_inst_n100), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n102) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U325 ( .A(
        wrap_act_buffer_inst_act_if_inst_n175), .B(
        wrap_act_buffer_inst_act_if_inst_n167), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n101) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U324 ( .A(
        wrap_act_buffer_inst_act_if_inst_n211), .B(
        wrap_act_buffer_inst_act_if_inst_n199), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n100) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U323 ( .A(
        wrap_act_buffer_inst_act_if_inst_n98), .B(
        wrap_act_buffer_inst_act_if_inst_n97), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n99) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U322 ( .A(
        wrap_act_buffer_inst_act_if_inst_n263), .B(
        wrap_act_buffer_inst_act_if_inst_n235), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n98) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U321 ( .A(
        wrap_act_buffer_inst_act_if_inst_n191), .B(
        wrap_act_buffer_inst_act_if_inst_n183), .S(
        wrap_act_buffer_inst_act_if_inst_n309), .Z(
        wrap_act_buffer_inst_act_if_inst_n97) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U320 ( .A(
        wrap_act_buffer_inst_act_if_inst_n95), .B(
        wrap_act_buffer_inst_act_if_inst_n94), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n96) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U319 ( .A(
        wrap_act_buffer_inst_act_if_inst_n174), .B(
        wrap_act_buffer_inst_act_if_inst_n166), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n95) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U318 ( .A(
        wrap_act_buffer_inst_act_if_inst_n208), .B(
        wrap_act_buffer_inst_act_if_inst_n198), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n94) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U317 ( .A(
        wrap_act_buffer_inst_act_if_inst_n92), .B(
        wrap_act_buffer_inst_act_if_inst_n91), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n93) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U316 ( .A(
        wrap_act_buffer_inst_act_if_inst_n258), .B(
        wrap_act_buffer_inst_act_if_inst_n232), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n92) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U315 ( .A(
        wrap_act_buffer_inst_act_if_inst_n190), .B(
        wrap_act_buffer_inst_act_if_inst_n182), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n91) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U314 ( .A(
        wrap_act_buffer_inst_act_if_inst_n89), .B(
        wrap_act_buffer_inst_act_if_inst_n88), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n90) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U313 ( .A(
        wrap_act_buffer_inst_act_if_inst_n173), .B(
        wrap_act_buffer_inst_act_if_inst_n165), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n89) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U312 ( .A(
        wrap_act_buffer_inst_act_if_inst_n205), .B(
        wrap_act_buffer_inst_act_if_inst_n197), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n88) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U311 ( .A(
        wrap_act_buffer_inst_act_if_inst_n86), .B(
        wrap_act_buffer_inst_act_if_inst_n85), .S(
        wrap_act_buffer_inst_act_if_inst_n295), .Z(
        wrap_act_buffer_inst_act_if_inst_n87) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U310 ( .A(
        wrap_act_buffer_inst_act_if_inst_n253), .B(
        wrap_act_buffer_inst_act_if_inst_n229), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n86) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U309 ( .A(
        wrap_act_buffer_inst_act_if_inst_n189), .B(
        wrap_act_buffer_inst_act_if_inst_n181), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n85) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U308 ( .A(
        wrap_act_buffer_inst_act_if_inst_n83), .B(
        wrap_act_buffer_inst_act_if_inst_n82), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n84) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U307 ( .A(
        wrap_act_buffer_inst_act_if_inst_n172), .B(
        wrap_act_buffer_inst_act_if_inst_n288), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n83) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U306 ( .A(
        wrap_act_buffer_inst_act_if_inst_n204), .B(
        wrap_act_buffer_inst_act_if_inst_n196), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n82) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U305 ( .A(
        wrap_act_buffer_inst_act_if_inst_n80), .B(
        wrap_act_buffer_inst_act_if_inst_n79), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n81) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U304 ( .A(
        wrap_act_buffer_inst_act_if_inst_n250), .B(
        wrap_act_buffer_inst_act_if_inst_n226), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n80) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U303 ( .A(
        wrap_act_buffer_inst_act_if_inst_n188), .B(
        wrap_act_buffer_inst_act_if_inst_n180), .S(
        wrap_act_buffer_inst_act_if_inst_n308), .Z(
        wrap_act_buffer_inst_act_if_inst_n79) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U302 ( .A(
        wrap_act_buffer_inst_act_if_inst_n77), .B(
        wrap_act_buffer_inst_act_if_inst_n76), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n78) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U301 ( .A(
        wrap_act_buffer_inst_act_if_inst_n171), .B(
        wrap_act_buffer_inst_act_if_inst_n283), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n77) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U300 ( .A(
        wrap_act_buffer_inst_act_if_inst_n203), .B(
        wrap_act_buffer_inst_act_if_inst_n195), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n76) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U299 ( .A(
        wrap_act_buffer_inst_act_if_inst_n74), .B(
        wrap_act_buffer_inst_act_if_inst_n73), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n75) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U298 ( .A(
        wrap_act_buffer_inst_act_if_inst_n247), .B(
        wrap_act_buffer_inst_act_if_inst_n223), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n74) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U297 ( .A(
        wrap_act_buffer_inst_act_if_inst_n187), .B(
        wrap_act_buffer_inst_act_if_inst_n179), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n73) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U296 ( .A(
        wrap_act_buffer_inst_act_if_inst_n71), .B(
        wrap_act_buffer_inst_act_if_inst_n70), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n72) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U295 ( .A(
        wrap_act_buffer_inst_act_if_inst_n170), .B(
        wrap_act_buffer_inst_act_if_inst_n278), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n71) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U294 ( .A(
        wrap_act_buffer_inst_act_if_inst_n202), .B(
        wrap_act_buffer_inst_act_if_inst_n194), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n70) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U293 ( .A(
        wrap_act_buffer_inst_act_if_inst_n68), .B(
        wrap_act_buffer_inst_act_if_inst_n67), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n69) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U292 ( .A(
        wrap_act_buffer_inst_act_if_inst_n244), .B(
        wrap_act_buffer_inst_act_if_inst_n220), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n68) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U291 ( .A(
        wrap_act_buffer_inst_act_if_inst_n186), .B(
        wrap_act_buffer_inst_act_if_inst_n178), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n67) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U290 ( .A(
        wrap_act_buffer_inst_act_if_inst_n65), .B(
        wrap_act_buffer_inst_act_if_inst_n64), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n66) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U289 ( .A(
        wrap_act_buffer_inst_act_if_inst_n169), .B(
        wrap_act_buffer_inst_act_if_inst_n273), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n65) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U288 ( .A(
        wrap_act_buffer_inst_act_if_inst_n201), .B(
        wrap_act_buffer_inst_act_if_inst_n193), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n64) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U287 ( .A(
        wrap_act_buffer_inst_act_if_inst_n62), .B(
        wrap_act_buffer_inst_act_if_inst_n61), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n63) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U286 ( .A(
        wrap_act_buffer_inst_act_if_inst_n241), .B(
        wrap_act_buffer_inst_act_if_inst_n217), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n62) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U285 ( .A(
        wrap_act_buffer_inst_act_if_inst_n185), .B(
        wrap_act_buffer_inst_act_if_inst_n177), .S(
        wrap_act_buffer_inst_act_if_inst_n307), .Z(
        wrap_act_buffer_inst_act_if_inst_n61) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U284 ( .A(
        wrap_act_buffer_inst_act_if_inst_n59), .B(
        wrap_act_buffer_inst_act_if_inst_n58), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n60) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U283 ( .A(
        wrap_act_buffer_inst_act_if_inst_n168), .B(
        wrap_act_buffer_inst_act_if_inst_n268), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n59) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U282 ( .A(
        wrap_act_buffer_inst_act_if_inst_n200), .B(
        wrap_act_buffer_inst_act_if_inst_n192), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n58) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U281 ( .A(
        wrap_act_buffer_inst_act_if_inst_n56), .B(
        wrap_act_buffer_inst_act_if_inst_n55), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n57) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U280 ( .A(
        wrap_act_buffer_inst_act_if_inst_n238), .B(
        wrap_act_buffer_inst_act_if_inst_n214), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n56) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U279 ( .A(
        wrap_act_buffer_inst_act_if_inst_n184), .B(
        wrap_act_buffer_inst_act_if_inst_n176), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n55) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U278 ( .A(
        wrap_act_buffer_inst_act_if_inst_n53), .B(
        wrap_act_buffer_inst_act_if_inst_n52), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n54) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U277 ( .A(
        wrap_act_buffer_inst_act_if_inst_n167), .B(
        wrap_act_buffer_inst_act_if_inst_n263), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n53) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U276 ( .A(
        wrap_act_buffer_inst_act_if_inst_n199), .B(
        wrap_act_buffer_inst_act_if_inst_n191), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n52) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U275 ( .A(
        wrap_act_buffer_inst_act_if_inst_n50), .B(
        wrap_act_buffer_inst_act_if_inst_n49), .S(
        wrap_act_buffer_inst_act_if_inst_n294), .Z(
        wrap_act_buffer_inst_act_if_inst_n51) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U274 ( .A(
        wrap_act_buffer_inst_act_if_inst_n235), .B(
        wrap_act_buffer_inst_act_if_inst_n211), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n50) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U273 ( .A(
        wrap_act_buffer_inst_act_if_inst_n183), .B(
        wrap_act_buffer_inst_act_if_inst_n175), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n49) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U272 ( .A(
        wrap_act_buffer_inst_act_if_inst_n47), .B(
        wrap_act_buffer_inst_act_if_inst_n46), .S(
        wrap_act_buffer_inst_act_if_inst_n293), .Z(
        wrap_act_buffer_inst_act_if_inst_n48) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U271 ( .A(
        wrap_act_buffer_inst_act_if_inst_n166), .B(
        wrap_act_buffer_inst_act_if_inst_n258), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n47) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U270 ( .A(
        wrap_act_buffer_inst_act_if_inst_n198), .B(
        wrap_act_buffer_inst_act_if_inst_n190), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n46) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U269 ( .A(
        wrap_act_buffer_inst_act_if_inst_n44), .B(
        wrap_act_buffer_inst_act_if_inst_n43), .S(
        wrap_act_buffer_inst_act_if_inst_n293), .Z(
        wrap_act_buffer_inst_act_if_inst_n45) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U268 ( .A(
        wrap_act_buffer_inst_act_if_inst_n232), .B(
        wrap_act_buffer_inst_act_if_inst_n208), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n44) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U267 ( .A(
        wrap_act_buffer_inst_act_if_inst_n182), .B(
        wrap_act_buffer_inst_act_if_inst_n174), .S(
        wrap_act_buffer_inst_act_if_inst_n306), .Z(
        wrap_act_buffer_inst_act_if_inst_n43) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U266 ( .A(
        wrap_act_buffer_inst_act_if_inst_n41), .B(
        wrap_act_buffer_inst_act_if_inst_n40), .S(
        wrap_act_buffer_inst_act_if_inst_n293), .Z(
        wrap_act_buffer_inst_act_if_inst_n42) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U265 ( .A(
        wrap_act_buffer_inst_act_if_inst_n165), .B(
        wrap_act_buffer_inst_act_if_inst_n253), .S(
        wrap_act_buffer_inst_act_if_inst_n305), .Z(
        wrap_act_buffer_inst_act_if_inst_n41) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U264 ( .A(
        wrap_act_buffer_inst_act_if_inst_n197), .B(
        wrap_act_buffer_inst_act_if_inst_n189), .S(
        wrap_act_buffer_inst_act_if_inst_n305), .Z(
        wrap_act_buffer_inst_act_if_inst_n40) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U263 ( .A(
        wrap_act_buffer_inst_act_if_inst_n2), .B(
        wrap_act_buffer_inst_act_if_inst_n1), .S(
        wrap_act_buffer_inst_act_if_inst_n293), .Z(
        wrap_act_buffer_inst_act_if_inst_n39) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U262 ( .A(
        wrap_act_buffer_inst_act_if_inst_n229), .B(
        wrap_act_buffer_inst_act_if_inst_n205), .S(
        wrap_act_buffer_inst_act_if_inst_n305), .Z(
        wrap_act_buffer_inst_act_if_inst_n2) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U261 ( .A(
        wrap_act_buffer_inst_act_if_inst_n181), .B(
        wrap_act_buffer_inst_act_if_inst_n173), .S(
        wrap_act_buffer_inst_act_if_inst_n305), .Z(
        wrap_act_buffer_inst_act_if_inst_n1) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U260 ( .A(
        wrap_act_buffer_inst_act_if_inst_n289), .B(
        wrap_act_buffer_inst_act_if_inst_n228), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data1[7]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U259 ( .A(
        wrap_act_buffer_inst_act_if_inst_n284), .B(
        wrap_act_buffer_inst_act_if_inst_n225), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data1[6]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U258 ( .A(
        wrap_act_buffer_inst_act_if_inst_n279), .B(
        wrap_act_buffer_inst_act_if_inst_n222), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data1[5]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U257 ( .A(
        wrap_act_buffer_inst_act_if_inst_n274), .B(
        wrap_act_buffer_inst_act_if_inst_n219), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data1[4]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U256 ( .A(
        wrap_act_buffer_inst_act_if_inst_n269), .B(
        wrap_act_buffer_inst_act_if_inst_n216), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data1[3]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U255 ( .A(
        wrap_act_buffer_inst_act_if_inst_n264), .B(
        wrap_act_buffer_inst_act_if_inst_n213), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data1[2]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U254 ( .A(
        wrap_act_buffer_inst_act_if_inst_n259), .B(
        wrap_act_buffer_inst_act_if_inst_n210), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data1[1]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U253 ( .A(
        wrap_act_buffer_inst_act_if_inst_n254), .B(
        wrap_act_buffer_inst_act_if_inst_n207), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data1[0]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U252 ( .A(
        wrap_act_buffer_inst_act_if_inst_n251), .B(
        wrap_act_buffer_inst_act_if_inst_n292), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data2[7]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U251 ( .A(
        wrap_act_buffer_inst_act_if_inst_n248), .B(
        wrap_act_buffer_inst_act_if_inst_n287), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data2[6]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U250 ( .A(
        wrap_act_buffer_inst_act_if_inst_n245), .B(
        wrap_act_buffer_inst_act_if_inst_n282), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data2[5]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U249 ( .A(
        wrap_act_buffer_inst_act_if_inst_n242), .B(
        wrap_act_buffer_inst_act_if_inst_n277), .S(
        wrap_act_buffer_inst_act_if_inst_n304), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data2[4]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U248 ( .A(
        wrap_act_buffer_inst_act_if_inst_n239), .B(
        wrap_act_buffer_inst_act_if_inst_n272), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data2[3]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U247 ( .A(
        wrap_act_buffer_inst_act_if_inst_n236), .B(
        wrap_act_buffer_inst_act_if_inst_n267), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data2[2]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U246 ( .A(
        wrap_act_buffer_inst_act_if_inst_n233), .B(
        wrap_act_buffer_inst_act_if_inst_n262), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data2[1]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U245 ( .A(
        wrap_act_buffer_inst_act_if_inst_n230), .B(
        wrap_act_buffer_inst_act_if_inst_n257), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data2[0]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U244 ( .A(
        wrap_act_buffer_inst_act_if_inst_n228), .B(
        wrap_act_buffer_inst_act_if_inst_n290), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data3[7]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U243 ( .A(
        wrap_act_buffer_inst_act_if_inst_n225), .B(
        wrap_act_buffer_inst_act_if_inst_n285), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data3[6]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U242 ( .A(
        wrap_act_buffer_inst_act_if_inst_n222), .B(
        wrap_act_buffer_inst_act_if_inst_n280), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data3[5]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U241 ( .A(
        wrap_act_buffer_inst_act_if_inst_n219), .B(
        wrap_act_buffer_inst_act_if_inst_n275), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data3[4]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U240 ( .A(
        wrap_act_buffer_inst_act_if_inst_n216), .B(
        wrap_act_buffer_inst_act_if_inst_n270), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data3[3]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U239 ( .A(
        wrap_act_buffer_inst_act_if_inst_n213), .B(
        wrap_act_buffer_inst_act_if_inst_n265), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data3[2]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U238 ( .A(
        wrap_act_buffer_inst_act_if_inst_n210), .B(
        wrap_act_buffer_inst_act_if_inst_n260), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data3[1]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U237 ( .A(
        wrap_act_buffer_inst_act_if_inst_n207), .B(
        wrap_act_buffer_inst_act_if_inst_n255), .S(
        wrap_act_buffer_inst_act_if_inst_n303), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data3[0]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U236 ( .A(
        wrap_act_buffer_inst_act_if_inst_n292), .B(
        wrap_act_buffer_inst_act_if_inst_n252), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data4[7]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U235 ( .A(
        wrap_act_buffer_inst_act_if_inst_n287), .B(
        wrap_act_buffer_inst_act_if_inst_n249), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data4[6]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U234 ( .A(
        wrap_act_buffer_inst_act_if_inst_n282), .B(
        wrap_act_buffer_inst_act_if_inst_n246), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data4[5]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U233 ( .A(
        wrap_act_buffer_inst_act_if_inst_n277), .B(
        wrap_act_buffer_inst_act_if_inst_n243), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data4[4]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U232 ( .A(
        wrap_act_buffer_inst_act_if_inst_n272), .B(
        wrap_act_buffer_inst_act_if_inst_n240), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data4[3]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U231 ( .A(
        wrap_act_buffer_inst_act_if_inst_n267), .B(
        wrap_act_buffer_inst_act_if_inst_n237), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data4[2]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U230 ( .A(
        wrap_act_buffer_inst_act_if_inst_n262), .B(
        wrap_act_buffer_inst_act_if_inst_n234), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data4[1]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U229 ( .A(
        wrap_act_buffer_inst_act_if_inst_n257), .B(
        wrap_act_buffer_inst_act_if_inst_n231), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data4[0]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U228 ( .A(
        wrap_act_buffer_inst_act_if_inst_n290), .B(
        wrap_act_buffer_inst_act_if_inst_n227), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data5[7]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U227 ( .A(
        wrap_act_buffer_inst_act_if_inst_n285), .B(
        wrap_act_buffer_inst_act_if_inst_n224), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data5[6]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U226 ( .A(
        wrap_act_buffer_inst_act_if_inst_n280), .B(
        wrap_act_buffer_inst_act_if_inst_n221), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data5[5]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U225 ( .A(
        wrap_act_buffer_inst_act_if_inst_n275), .B(
        wrap_act_buffer_inst_act_if_inst_n218), .S(
        wrap_act_buffer_inst_act_if_inst_n302), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data5[4]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U224 ( .A(
        wrap_act_buffer_inst_act_if_inst_n270), .B(
        wrap_act_buffer_inst_act_if_inst_n215), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data5[3]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U223 ( .A(
        wrap_act_buffer_inst_act_if_inst_n265), .B(
        wrap_act_buffer_inst_act_if_inst_n212), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data5[2]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U222 ( .A(
        wrap_act_buffer_inst_act_if_inst_n260), .B(
        wrap_act_buffer_inst_act_if_inst_n209), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data5[1]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U221 ( .A(
        wrap_act_buffer_inst_act_if_inst_n255), .B(
        wrap_act_buffer_inst_act_if_inst_n206), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data5[0]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U220 ( .A(
        wrap_act_buffer_inst_act_if_inst_n252), .B(
        wrap_act_buffer_inst_act_if_inst_n291), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data6[7]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U219 ( .A(
        wrap_act_buffer_inst_act_if_inst_n249), .B(
        wrap_act_buffer_inst_act_if_inst_n286), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data6[6]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U218 ( .A(
        wrap_act_buffer_inst_act_if_inst_n246), .B(
        wrap_act_buffer_inst_act_if_inst_n281), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data6[5]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U217 ( .A(
        wrap_act_buffer_inst_act_if_inst_n243), .B(
        wrap_act_buffer_inst_act_if_inst_n276), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data6[4]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U216 ( .A(
        wrap_act_buffer_inst_act_if_inst_n240), .B(
        wrap_act_buffer_inst_act_if_inst_n271), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data6[3]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U215 ( .A(
        wrap_act_buffer_inst_act_if_inst_n237), .B(
        wrap_act_buffer_inst_act_if_inst_n266), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data6[2]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U214 ( .A(
        wrap_act_buffer_inst_act_if_inst_n234), .B(
        wrap_act_buffer_inst_act_if_inst_n261), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data6[1]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U213 ( .A(
        wrap_act_buffer_inst_act_if_inst_n231), .B(
        wrap_act_buffer_inst_act_if_inst_n256), .S(
        wrap_act_buffer_inst_act_if_inst_n301), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data6[0]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U212 ( .A(
        wrap_act_buffer_inst_act_if_inst_n227), .B(
        wrap_act_buffer_inst_act_if_inst_n289), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data7[7]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U211 ( .A(
        wrap_act_buffer_inst_act_if_inst_n224), .B(
        wrap_act_buffer_inst_act_if_inst_n284), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data7[6]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U210 ( .A(
        wrap_act_buffer_inst_act_if_inst_n221), .B(
        wrap_act_buffer_inst_act_if_inst_n279), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data7[5]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U209 ( .A(
        wrap_act_buffer_inst_act_if_inst_n218), .B(
        wrap_act_buffer_inst_act_if_inst_n274), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data7[4]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U208 ( .A(
        wrap_act_buffer_inst_act_if_inst_n215), .B(
        wrap_act_buffer_inst_act_if_inst_n269), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data7[3]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U207 ( .A(
        wrap_act_buffer_inst_act_if_inst_n212), .B(
        wrap_act_buffer_inst_act_if_inst_n264), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data7[2]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U206 ( .A(
        wrap_act_buffer_inst_act_if_inst_n209), .B(
        wrap_act_buffer_inst_act_if_inst_n259), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data7[1]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U205 ( .A(
        wrap_act_buffer_inst_act_if_inst_n206), .B(
        wrap_act_buffer_inst_act_if_inst_n254), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data7[0]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U204 ( .A(
        wrap_act_buffer_inst_act_if_inst_n291), .B(
        wrap_act_buffer_inst_act_if_inst_n251), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data8[7]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U203 ( .A(
        wrap_act_buffer_inst_act_if_inst_n286), .B(
        wrap_act_buffer_inst_act_if_inst_n248), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data8[6]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U202 ( .A(
        wrap_act_buffer_inst_act_if_inst_n281), .B(
        wrap_act_buffer_inst_act_if_inst_n245), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data8[5]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U201 ( .A(
        wrap_act_buffer_inst_act_if_inst_n276), .B(
        wrap_act_buffer_inst_act_if_inst_n242), .S(
        wrap_act_buffer_inst_act_if_inst_n300), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data8[4]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U200 ( .A(
        wrap_act_buffer_inst_act_if_inst_n271), .B(
        wrap_act_buffer_inst_act_if_inst_n239), .S(
        wrap_act_buffer_inst_act_if_inst_n299), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data8[3]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U199 ( .A(
        wrap_act_buffer_inst_act_if_inst_n266), .B(
        wrap_act_buffer_inst_act_if_inst_n236), .S(
        wrap_act_buffer_inst_act_if_inst_n299), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data8[2]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U198 ( .A(
        wrap_act_buffer_inst_act_if_inst_n261), .B(
        wrap_act_buffer_inst_act_if_inst_n233), .S(
        wrap_act_buffer_inst_act_if_inst_n299), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data8[1]) );
  MUX2_X1 wrap_act_buffer_inst_act_if_inst_U197 ( .A(
        wrap_act_buffer_inst_act_if_inst_n256), .B(
        wrap_act_buffer_inst_act_if_inst_n230), .S(
        wrap_act_buffer_inst_act_if_inst_n299), .Z(
        wrap_act_buffer_inst_act_if_inst_int_data8[0]) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U196 ( .A(1'b0), .ZN(
        wrap_act_buffer_inst_act_if_inst_n311) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U195 ( .A(ps_int_hmode_cnt[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n312) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U194 ( .A(int_npu_ptr[0]), .Z(
        wrap_act_buffer_inst_act_if_inst_n310) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U193 ( .A(int_npu_ptr[2]), .Z(
        wrap_act_buffer_inst_act_if_inst_n295) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U192 ( .A(int_npu_ptr[2]), .Z(
        wrap_act_buffer_inst_act_if_inst_n296) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U191 ( .A(int_npu_ptr[2]), .Z(
        wrap_act_buffer_inst_act_if_inst_n294) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U190 ( .A(int_npu_ptr[2]), .Z(
        wrap_act_buffer_inst_act_if_inst_n298) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U189 ( .A(int_npu_ptr[2]), .Z(
        wrap_act_buffer_inst_act_if_inst_n297) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U188 ( .A(int_npu_ptr[1]), .Z(
        wrap_act_buffer_inst_act_if_inst_n304) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U187 ( .A(int_npu_ptr[1]), .Z(
        wrap_act_buffer_inst_act_if_inst_n303) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U186 ( .A(int_npu_ptr[1]), .Z(
        wrap_act_buffer_inst_act_if_inst_n302) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U185 ( .A(int_npu_ptr[1]), .Z(
        wrap_act_buffer_inst_act_if_inst_n301) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U184 ( .A(int_npu_ptr[1]), .Z(
        wrap_act_buffer_inst_act_if_inst_n300) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U183 ( .A(int_npu_ptr[0]), .Z(
        wrap_act_buffer_inst_act_if_inst_n309) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U182 ( .A(int_npu_ptr[0]), .Z(
        wrap_act_buffer_inst_act_if_inst_n308) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U181 ( .A(int_npu_ptr[0]), .Z(
        wrap_act_buffer_inst_act_if_inst_n306) );
  BUF_X1 wrap_act_buffer_inst_act_if_inst_U180 ( .A(int_npu_ptr[0]), .Z(
        wrap_act_buffer_inst_act_if_inst_n307) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U179 ( .A(
        wrap_act_buffer_inst_int_i_data_if1[4]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n273) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U178 ( .A(
        wrap_act_buffer_inst_int_i_data_if6[3]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n184) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U177 ( .A(
        wrap_act_buffer_inst_int_i_data_if7[3]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n176) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U176 ( .A(
        wrap_act_buffer_inst_int_i_data_if8[3]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n168) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U175 ( .A(
        wrap_act_buffer_inst_int_i_data_if5[5]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n194) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U174 ( .A(
        wrap_act_buffer_inst_int_i_data_if6[5]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n186) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U173 ( .A(
        wrap_act_buffer_inst_int_i_data_if7[5]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n178) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U172 ( .A(
        wrap_act_buffer_inst_int_i_data_if5[7]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n196) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U171 ( .A(
        wrap_act_buffer_inst_int_i_data_if6[7]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n188) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U170 ( .A(
        wrap_act_buffer_inst_int_i_data_if8[7]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n172) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U169 ( .A(
        wrap_act_buffer_inst_int_i_data_if7[7]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n180) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U168 ( .A(
        wrap_act_buffer_inst_int_i_data_if6[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n182) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U167 ( .A(
        wrap_act_buffer_inst_int_i_data_if7[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n174) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U166 ( .A(
        wrap_act_buffer_inst_int_i_data_if8[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n166) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U165 ( .A(
        wrap_act_buffer_inst_int_i_data_if6[2]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n183) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U164 ( .A(
        wrap_act_buffer_inst_int_i_data_if7[2]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n175) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U163 ( .A(
        wrap_act_buffer_inst_int_i_data_if8[2]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n167) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U162 ( .A(
        wrap_act_buffer_inst_int_i_data_if6[4]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n185) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U161 ( .A(
        wrap_act_buffer_inst_int_i_data_if5[4]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n193) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U160 ( .A(
        wrap_act_buffer_inst_int_i_data_if7[4]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n177) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U159 ( .A(
        wrap_act_buffer_inst_int_i_data_if5[6]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n195) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U158 ( .A(
        wrap_act_buffer_inst_int_i_data_if6[6]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n187) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U157 ( .A(
        wrap_act_buffer_inst_int_i_data_if8[6]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n171) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U156 ( .A(
        wrap_act_buffer_inst_int_i_data_if7[6]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n179) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U155 ( .A(
        wrap_act_buffer_inst_int_i_data_if6[0]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n181) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U154 ( .A(
        wrap_act_buffer_inst_int_i_data_if8[0]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n165) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U153 ( .A(
        wrap_act_buffer_inst_int_i_data_if7[0]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n173) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U152 ( .A(
        wrap_act_buffer_inst_int_i_data_if1[3]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n268) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U151 ( .A(
        wrap_act_buffer_inst_int_i_data_if2[3]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n238) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U150 ( .A(
        wrap_act_buffer_inst_int_i_data_if1[5]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n278) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U149 ( .A(
        wrap_act_buffer_inst_int_i_data_if1[7]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n288) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U148 ( .A(
        wrap_act_buffer_inst_int_i_data_if1[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n258) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U147 ( .A(
        wrap_act_buffer_inst_int_i_data_if2[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n232) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U146 ( .A(
        wrap_act_buffer_inst_int_i_data_if1[2]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n263) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U145 ( .A(
        wrap_act_buffer_inst_int_i_data_if2[2]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n235) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U144 ( .A(
        wrap_act_buffer_inst_int_i_data_if1[6]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n283) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U143 ( .A(
        wrap_act_buffer_inst_int_i_data_if1[0]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n253) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U142 ( .A(
        wrap_act_buffer_inst_int_i_data_if2[0]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n229) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U141 ( .A(
        wrap_act_buffer_inst_int_i_data_if8[5]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n170) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U140 ( .A(
        wrap_act_buffer_inst_int_i_data_if8[4]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n169) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U139 ( .A(
        wrap_act_buffer_inst_int_i_data_if5[3]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n192) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U138 ( .A(
        wrap_act_buffer_inst_int_i_data_if3[3]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n214) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U137 ( .A(
        wrap_act_buffer_inst_int_i_data_if4[3]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n200) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U136 ( .A(
        wrap_act_buffer_inst_int_i_data_if2[5]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n244) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U135 ( .A(
        wrap_act_buffer_inst_int_i_data_if3[5]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n220) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U134 ( .A(
        wrap_act_buffer_inst_int_i_data_if4[5]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n202) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U133 ( .A(
        wrap_act_buffer_inst_int_i_data_if2[7]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n250) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U132 ( .A(
        wrap_act_buffer_inst_int_i_data_if3[7]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n226) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U131 ( .A(
        wrap_act_buffer_inst_int_i_data_if4[7]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n204) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U130 ( .A(
        wrap_act_buffer_inst_int_i_data_if5[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n190) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U129 ( .A(
        wrap_act_buffer_inst_int_i_data_if3[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n208) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U128 ( .A(
        wrap_act_buffer_inst_int_i_data_if4[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n198) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U127 ( .A(
        wrap_act_buffer_inst_int_i_data_if5[2]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n191) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U126 ( .A(
        wrap_act_buffer_inst_int_i_data_if3[2]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n211) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U125 ( .A(
        wrap_act_buffer_inst_int_i_data_if4[2]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n199) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U124 ( .A(
        wrap_act_buffer_inst_int_i_data_if2[4]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n241) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U123 ( .A(
        wrap_act_buffer_inst_int_i_data_if3[4]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n217) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U122 ( .A(
        wrap_act_buffer_inst_int_i_data_if4[4]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n201) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U121 ( .A(
        wrap_act_buffer_inst_int_i_data_if2[6]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n247) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U120 ( .A(
        wrap_act_buffer_inst_int_i_data_if3[6]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n223) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U119 ( .A(
        wrap_act_buffer_inst_int_i_data_if4[6]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n203) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U118 ( .A(
        wrap_act_buffer_inst_int_i_data_if5[0]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n189) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U117 ( .A(
        wrap_act_buffer_inst_int_i_data_if4[0]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n197) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U116 ( .A(
        wrap_act_buffer_inst_int_i_data_if3[0]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n205) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U115 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data8[7]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data8[1]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n4) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U114 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data8[3]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data8[5]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n3) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U113 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n3), .A2(
        wrap_act_buffer_inst_act_if_inst_n4), .ZN(int_i_data_h_npu[1]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U112 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data8[6]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data8[0]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n10) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U111 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data8[2]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data8[4]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n9) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U110 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n9), .A2(
        wrap_act_buffer_inst_act_if_inst_n10), .ZN(int_i_data_h_npu[0]) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U109 ( .A(
        wrap_act_buffer_inst_act_if_inst_n160), .ZN(
        wrap_act_buffer_inst_act_if_inst_n216) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U108 ( .A(
        wrap_act_buffer_inst_act_if_inst_n162), .ZN(
        wrap_act_buffer_inst_act_if_inst_n222) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U107 ( .A(
        wrap_act_buffer_inst_act_if_inst_n164), .ZN(
        wrap_act_buffer_inst_act_if_inst_n228) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U106 ( .A(
        wrap_act_buffer_inst_act_if_inst_n158), .ZN(
        wrap_act_buffer_inst_act_if_inst_n210) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U105 ( .A(
        wrap_act_buffer_inst_act_if_inst_n159), .ZN(
        wrap_act_buffer_inst_act_if_inst_n213) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U104 ( .A(
        wrap_act_buffer_inst_act_if_inst_n161), .ZN(
        wrap_act_buffer_inst_act_if_inst_n219) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U103 ( .A(
        wrap_act_buffer_inst_act_if_inst_n163), .ZN(
        wrap_act_buffer_inst_act_if_inst_n225) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U102 ( .A(
        wrap_act_buffer_inst_act_if_inst_n157), .ZN(
        wrap_act_buffer_inst_act_if_inst_n207) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U101 ( .A(
        wrap_act_buffer_inst_act_if_inst_n152), .ZN(
        wrap_act_buffer_inst_act_if_inst_n272) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U100 ( .A(
        wrap_act_buffer_inst_act_if_inst_n154), .ZN(
        wrap_act_buffer_inst_act_if_inst_n282) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U99 ( .A(
        wrap_act_buffer_inst_act_if_inst_n156), .ZN(
        wrap_act_buffer_inst_act_if_inst_n292) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U98 ( .A(
        wrap_act_buffer_inst_act_if_inst_n45), .ZN(
        wrap_act_buffer_inst_act_if_inst_n233) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U97 ( .A(
        wrap_act_buffer_inst_act_if_inst_n150), .ZN(
        wrap_act_buffer_inst_act_if_inst_n262) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U96 ( .A(
        wrap_act_buffer_inst_act_if_inst_n151), .ZN(
        wrap_act_buffer_inst_act_if_inst_n267) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U95 ( .A(
        wrap_act_buffer_inst_act_if_inst_n153), .ZN(
        wrap_act_buffer_inst_act_if_inst_n277) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U94 ( .A(
        wrap_act_buffer_inst_act_if_inst_n155), .ZN(
        wrap_act_buffer_inst_act_if_inst_n287) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U93 ( .A(
        wrap_act_buffer_inst_act_if_inst_n39), .ZN(
        wrap_act_buffer_inst_act_if_inst_n230) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U92 ( .A(
        wrap_act_buffer_inst_act_if_inst_n149), .ZN(
        wrap_act_buffer_inst_act_if_inst_n257) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U91 ( .A(
        wrap_act_buffer_inst_act_if_inst_n144), .ZN(
        wrap_act_buffer_inst_act_if_inst_n270) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U90 ( .A(
        wrap_act_buffer_inst_act_if_inst_n146), .ZN(
        wrap_act_buffer_inst_act_if_inst_n280) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U89 ( .A(
        wrap_act_buffer_inst_act_if_inst_n148), .ZN(
        wrap_act_buffer_inst_act_if_inst_n290) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U88 ( .A(
        wrap_act_buffer_inst_act_if_inst_n142), .ZN(
        wrap_act_buffer_inst_act_if_inst_n260) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U87 ( .A(
        wrap_act_buffer_inst_act_if_inst_n143), .ZN(
        wrap_act_buffer_inst_act_if_inst_n265) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U86 ( .A(
        wrap_act_buffer_inst_act_if_inst_n145), .ZN(
        wrap_act_buffer_inst_act_if_inst_n275) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U85 ( .A(
        wrap_act_buffer_inst_act_if_inst_n147), .ZN(
        wrap_act_buffer_inst_act_if_inst_n285) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U84 ( .A(
        wrap_act_buffer_inst_act_if_inst_n141), .ZN(
        wrap_act_buffer_inst_act_if_inst_n255) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U83 ( .A(
        wrap_act_buffer_inst_act_if_inst_n48), .ZN(
        wrap_act_buffer_inst_act_if_inst_n261) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U82 ( .A(
        wrap_act_buffer_inst_act_if_inst_n42), .ZN(
        wrap_act_buffer_inst_act_if_inst_n256) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U81 ( .A(
        wrap_act_buffer_inst_act_if_inst_n105), .ZN(
        wrap_act_buffer_inst_act_if_inst_n269) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U80 ( .A(
        wrap_act_buffer_inst_act_if_inst_n117), .ZN(
        wrap_act_buffer_inst_act_if_inst_n279) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U79 ( .A(
        wrap_act_buffer_inst_act_if_inst_n129), .ZN(
        wrap_act_buffer_inst_act_if_inst_n289) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U78 ( .A(
        wrap_act_buffer_inst_act_if_inst_n93), .ZN(
        wrap_act_buffer_inst_act_if_inst_n259) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U77 ( .A(
        wrap_act_buffer_inst_act_if_inst_n99), .ZN(
        wrap_act_buffer_inst_act_if_inst_n264) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U76 ( .A(
        wrap_act_buffer_inst_act_if_inst_n111), .ZN(
        wrap_act_buffer_inst_act_if_inst_n274) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U75 ( .A(
        wrap_act_buffer_inst_act_if_inst_n123), .ZN(
        wrap_act_buffer_inst_act_if_inst_n284) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U74 ( .A(
        wrap_act_buffer_inst_act_if_inst_n87), .ZN(
        wrap_act_buffer_inst_act_if_inst_n254) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U73 ( .A(
        wrap_act_buffer_inst_act_if_inst_n57), .ZN(
        wrap_act_buffer_inst_act_if_inst_n239) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U72 ( .A(
        wrap_act_buffer_inst_act_if_inst_n69), .ZN(
        wrap_act_buffer_inst_act_if_inst_n245) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U71 ( .A(
        wrap_act_buffer_inst_act_if_inst_n81), .ZN(
        wrap_act_buffer_inst_act_if_inst_n251) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U70 ( .A(
        wrap_act_buffer_inst_act_if_inst_n51), .ZN(
        wrap_act_buffer_inst_act_if_inst_n236) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U69 ( .A(
        wrap_act_buffer_inst_act_if_inst_n63), .ZN(
        wrap_act_buffer_inst_act_if_inst_n242) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U68 ( .A(
        wrap_act_buffer_inst_act_if_inst_n75), .ZN(
        wrap_act_buffer_inst_act_if_inst_n248) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U67 ( .A(
        wrap_act_buffer_inst_act_if_inst_n136), .ZN(
        wrap_act_buffer_inst_act_if_inst_n240) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U66 ( .A(
        wrap_act_buffer_inst_act_if_inst_n138), .ZN(
        wrap_act_buffer_inst_act_if_inst_n246) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U65 ( .A(
        wrap_act_buffer_inst_act_if_inst_n140), .ZN(
        wrap_act_buffer_inst_act_if_inst_n252) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U64 ( .A(
        wrap_act_buffer_inst_act_if_inst_n134), .ZN(
        wrap_act_buffer_inst_act_if_inst_n234) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U63 ( .A(
        wrap_act_buffer_inst_act_if_inst_n135), .ZN(
        wrap_act_buffer_inst_act_if_inst_n237) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U62 ( .A(
        wrap_act_buffer_inst_act_if_inst_n137), .ZN(
        wrap_act_buffer_inst_act_if_inst_n243) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U61 ( .A(
        wrap_act_buffer_inst_act_if_inst_n139), .ZN(
        wrap_act_buffer_inst_act_if_inst_n249) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U60 ( .A(
        wrap_act_buffer_inst_act_if_inst_n133), .ZN(
        wrap_act_buffer_inst_act_if_inst_n231) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U59 ( .A(
        wrap_act_buffer_inst_act_if_inst_n108), .ZN(
        wrap_act_buffer_inst_act_if_inst_n215) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U58 ( .A(
        wrap_act_buffer_inst_act_if_inst_n120), .ZN(
        wrap_act_buffer_inst_act_if_inst_n221) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U57 ( .A(
        wrap_act_buffer_inst_act_if_inst_n132), .ZN(
        wrap_act_buffer_inst_act_if_inst_n227) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U56 ( .A(
        wrap_act_buffer_inst_act_if_inst_n96), .ZN(
        wrap_act_buffer_inst_act_if_inst_n209) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U55 ( .A(
        wrap_act_buffer_inst_act_if_inst_n102), .ZN(
        wrap_act_buffer_inst_act_if_inst_n212) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U54 ( .A(
        wrap_act_buffer_inst_act_if_inst_n114), .ZN(
        wrap_act_buffer_inst_act_if_inst_n218) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U53 ( .A(
        wrap_act_buffer_inst_act_if_inst_n126), .ZN(
        wrap_act_buffer_inst_act_if_inst_n224) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U52 ( .A(
        wrap_act_buffer_inst_act_if_inst_n90), .ZN(
        wrap_act_buffer_inst_act_if_inst_n206) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U51 ( .A(
        wrap_act_buffer_inst_act_if_inst_n60), .ZN(
        wrap_act_buffer_inst_act_if_inst_n271) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U50 ( .A(
        wrap_act_buffer_inst_act_if_inst_n72), .ZN(
        wrap_act_buffer_inst_act_if_inst_n281) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U49 ( .A(
        wrap_act_buffer_inst_act_if_inst_n84), .ZN(
        wrap_act_buffer_inst_act_if_inst_n291) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U48 ( .A(
        wrap_act_buffer_inst_act_if_inst_n54), .ZN(
        wrap_act_buffer_inst_act_if_inst_n266) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U47 ( .A(
        wrap_act_buffer_inst_act_if_inst_n66), .ZN(
        wrap_act_buffer_inst_act_if_inst_n276) );
  INV_X1 wrap_act_buffer_inst_act_if_inst_U46 ( .A(
        wrap_act_buffer_inst_act_if_inst_n78), .ZN(
        wrap_act_buffer_inst_act_if_inst_n286) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U45 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data1[7]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data1[1]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n36) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U44 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data1[3]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data1[5]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n35) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U43 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n35), .A2(
        wrap_act_buffer_inst_act_if_inst_n36), .ZN(int_i_data_h_npu[15]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U42 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data1[6]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data1[0]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n38) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U41 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data1[2]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data1[4]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n37) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U40 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n37), .A2(
        wrap_act_buffer_inst_act_if_inst_n38), .ZN(int_i_data_h_npu[14]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U39 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data2[7]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data2[1]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n32) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U38 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data2[3]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data2[5]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n31) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U37 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n31), .A2(
        wrap_act_buffer_inst_act_if_inst_n32), .ZN(int_i_data_h_npu[13]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U36 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data2[6]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data2[0]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n34) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U35 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data2[2]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data2[4]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n33) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U34 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n33), .A2(
        wrap_act_buffer_inst_act_if_inst_n34), .ZN(int_i_data_h_npu[12]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U33 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data3[7]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data3[1]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n28) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U32 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data3[3]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data3[5]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n27) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U31 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n27), .A2(
        wrap_act_buffer_inst_act_if_inst_n28), .ZN(int_i_data_h_npu[11]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U30 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data3[6]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data3[0]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n30) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U29 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data3[2]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data3[4]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n29) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U28 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n29), .A2(
        wrap_act_buffer_inst_act_if_inst_n30), .ZN(int_i_data_h_npu[10]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U27 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data4[7]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data4[1]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n24) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U26 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data4[3]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data4[5]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n23) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U25 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n23), .A2(
        wrap_act_buffer_inst_act_if_inst_n24), .ZN(int_i_data_h_npu[9]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U24 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data4[6]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data4[0]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n26) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U23 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data4[2]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data4[4]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n25) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U22 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n25), .A2(
        wrap_act_buffer_inst_act_if_inst_n26), .ZN(int_i_data_h_npu[8]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U21 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data5[7]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data5[1]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n20) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U20 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data5[3]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data5[5]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n19) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U19 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n19), .A2(
        wrap_act_buffer_inst_act_if_inst_n20), .ZN(int_i_data_h_npu[7]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U18 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data5[6]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data5[0]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n22) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U17 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data5[2]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data5[4]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n21) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U16 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n21), .A2(
        wrap_act_buffer_inst_act_if_inst_n22), .ZN(int_i_data_h_npu[6]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U15 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data6[7]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data6[1]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n16) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U14 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data6[3]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data6[5]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n15) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U13 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n15), .A2(
        wrap_act_buffer_inst_act_if_inst_n16), .ZN(int_i_data_h_npu[5]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U12 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data6[6]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data6[0]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n18) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U11 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data6[2]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data6[4]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n17) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U10 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n17), .A2(
        wrap_act_buffer_inst_act_if_inst_n18), .ZN(int_i_data_h_npu[4]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U9 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data7[7]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data7[1]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n12) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U8 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data7[3]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data7[5]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n11) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U7 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n11), .A2(
        wrap_act_buffer_inst_act_if_inst_n12), .ZN(int_i_data_h_npu[3]) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U6 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data7[6]), .A2(
        wrap_act_buffer_inst_act_if_inst_n5), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data7[0]), .B2(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n14) );
  AOI22_X1 wrap_act_buffer_inst_act_if_inst_U5 ( .A1(
        wrap_act_buffer_inst_act_if_inst_int_data7[2]), .A2(
        wrap_act_buffer_inst_act_if_inst_n7), .B1(
        wrap_act_buffer_inst_act_if_inst_int_data7[4]), .B2(
        wrap_act_buffer_inst_act_if_inst_n8), .ZN(
        wrap_act_buffer_inst_act_if_inst_n13) );
  NAND2_X1 wrap_act_buffer_inst_act_if_inst_U4 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n13), .A2(
        wrap_act_buffer_inst_act_if_inst_n14), .ZN(int_i_data_h_npu[2]) );
  AND3_X1 wrap_act_buffer_inst_act_if_inst_U3 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n312), .A2(
        wrap_act_buffer_inst_act_if_inst_n311), .A3(ps_int_hmode_cnt[0]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n8) );
  AND3_X1 wrap_act_buffer_inst_act_if_inst_U2 ( .A1(ps_int_hmode_cnt[0]), .A2(
        wrap_act_buffer_inst_act_if_inst_n311), .A3(ps_int_hmode_cnt[1]), .ZN(
        wrap_act_buffer_inst_act_if_inst_n6) );
  NOR3_X4 wrap_act_buffer_inst_act_if_inst_U1 ( .A1(
        wrap_act_buffer_inst_act_if_inst_n7), .A2(
        wrap_act_buffer_inst_act_if_inst_n8), .A3(
        wrap_act_buffer_inst_act_if_inst_n6), .ZN(
        wrap_act_buffer_inst_act_if_inst_n5) );
  CLKGATETST_X1 wrap_act_buffer_inst_clk_gate_int_i_data_v_npu_reg_latch ( 
        .CK(ck), .E(ctrl_ldh_v_n), .SE(1'b0), .GCK(
        wrap_act_buffer_inst_net4501) );
  CLKBUF_X1 npu_inst_U189 ( .A(i_weight[1]), .Z(npu_inst_n101) );
  CLKBUF_X1 npu_inst_U188 ( .A(i_weight[0]), .Z(npu_inst_n95) );
  CLKBUF_X1 npu_inst_U187 ( .A(ps_int_ifmaps_ptr[0]), .Z(npu_inst_n54) );
  INV_X1 npu_inst_U186 ( .A(1'b0), .ZN(npu_inst_n111) );
  INV_X1 npu_inst_U185 ( .A(1'b0), .ZN(npu_inst_n110) );
  NAND2_X1 npu_inst_U184 ( .A1(npu_inst_n111), .A2(npu_inst_n110), .ZN(
        npu_inst_int_ckg[63]) );
  BUF_X1 npu_inst_U183 ( .A(ps_ctrl_wr_pipe), .Z(npu_inst_n10) );
  NAND2_X1 npu_inst_U182 ( .A1(npu_inst_n125), .A2(npu_inst_n118), .ZN(
        npu_inst_int_ckg[27]) );
  BUF_X1 npu_inst_U181 ( .A(ps_ctrl_ldh_v_n), .Z(npu_inst_n33) );
  BUF_X1 npu_inst_U180 ( .A(ps_ctrl_ldh_v_n), .Z(npu_inst_n32) );
  BUF_X1 npu_inst_U179 ( .A(ps_ctrl_wr_pipe), .Z(npu_inst_n8) );
  BUF_X1 npu_inst_U178 ( .A(ps_ctrl_wr_pipe), .Z(npu_inst_n9) );
  NAND2_X1 npu_inst_U177 ( .A1(npu_inst_n111), .A2(npu_inst_n118), .ZN(
        npu_inst_int_ckg[59]) );
  BUF_X1 npu_inst_U176 ( .A(ps_ctrl_en_npu), .Z(npu_inst_n48) );
  BUF_X1 npu_inst_U175 ( .A(ps_ctrl_en_npu), .Z(npu_inst_n43) );
  BUF_X1 npu_inst_U174 ( .A(ps_ctrl_en_npu), .Z(npu_inst_n44) );
  BUF_X1 npu_inst_U173 ( .A(ps_ctrl_en_npu), .Z(npu_inst_n45) );
  BUF_X1 npu_inst_U172 ( .A(ps_ctrl_en_npu), .Z(npu_inst_n46) );
  BUF_X1 npu_inst_U171 ( .A(ps_ctrl_en_npu), .Z(npu_inst_n47) );
  BUF_X1 npu_inst_U170 ( .A(i_weight[1]), .Z(npu_inst_n100) );
  BUF_X1 npu_inst_U169 ( .A(i_weight[0]), .Z(npu_inst_n94) );
  BUF_X1 npu_inst_U168 ( .A(i_weight[1]), .Z(npu_inst_n99) );
  BUF_X1 npu_inst_U167 ( .A(i_weight[0]), .Z(npu_inst_n93) );
  BUF_X1 npu_inst_U166 ( .A(i_weight[1]), .Z(npu_inst_n98) );
  BUF_X1 npu_inst_U165 ( .A(i_weight[0]), .Z(npu_inst_n92) );
  BUF_X1 npu_inst_U164 ( .A(i_weight[1]), .Z(npu_inst_n97) );
  BUF_X1 npu_inst_U163 ( .A(i_weight[0]), .Z(npu_inst_n91) );
  BUF_X1 npu_inst_U162 ( .A(i_weight[1]), .Z(npu_inst_n96) );
  BUF_X1 npu_inst_U161 ( .A(i_weight[0]), .Z(npu_inst_n90) );
  NAND2_X1 npu_inst_U160 ( .A1(npu_inst_n125), .A2(npu_inst_n110), .ZN(
        npu_inst_int_ckg[31]) );
  INV_X1 npu_inst_U159 ( .A(int_ckg_rmask[4]), .ZN(npu_inst_n125) );
  INV_X1 npu_inst_U158 ( .A(int_ckg_cmask[4]), .ZN(npu_inst_n118) );
  BUF_X1 npu_inst_U157 ( .A(ps_int_ifmaps_ptr[2]), .Z(npu_inst_n73) );
  BUF_X1 npu_inst_U156 ( .A(ps_int_ifmaps_ptr[2]), .Z(npu_inst_n71) );
  BUF_X1 npu_inst_U155 ( .A(ps_int_ifmaps_ptr[2]), .Z(npu_inst_n72) );
  NAND2_X1 npu_inst_U154 ( .A1(npu_inst_n111), .A2(npu_inst_n119), .ZN(
        npu_inst_int_ckg[58]) );
  NAND2_X1 npu_inst_U153 ( .A1(npu_inst_n111), .A2(npu_inst_n112), .ZN(
        npu_inst_int_ckg[62]) );
  NAND2_X1 npu_inst_U152 ( .A1(npu_inst_n111), .A2(npu_inst_n117), .ZN(
        npu_inst_int_ckg[61]) );
  NAND2_X1 npu_inst_U151 ( .A1(npu_inst_n111), .A2(npu_inst_n114), .ZN(
        npu_inst_int_ckg[60]) );
  NAND2_X1 npu_inst_U150 ( .A1(npu_inst_n111), .A2(npu_inst_n121), .ZN(
        npu_inst_int_ckg[56]) );
  BUF_X1 npu_inst_U149 ( .A(ps_int_ifmaps_ptr[1]), .Z(npu_inst_n56) );
  NAND2_X1 npu_inst_U148 ( .A1(npu_inst_n123), .A2(npu_inst_n110), .ZN(
        npu_inst_int_ckg[23]) );
  NAND2_X1 npu_inst_U147 ( .A1(npu_inst_n123), .A2(npu_inst_n112), .ZN(
        npu_inst_int_ckg[22]) );
  NAND2_X1 npu_inst_U146 ( .A1(npu_inst_n123), .A2(npu_inst_n117), .ZN(
        npu_inst_int_ckg[21]) );
  NAND2_X1 npu_inst_U145 ( .A1(npu_inst_n123), .A2(npu_inst_n114), .ZN(
        npu_inst_int_ckg[20]) );
  NAND2_X1 npu_inst_U144 ( .A1(npu_inst_n123), .A2(npu_inst_n118), .ZN(
        npu_inst_int_ckg[19]) );
  NAND2_X1 npu_inst_U143 ( .A1(npu_inst_n123), .A2(npu_inst_n119), .ZN(
        npu_inst_int_ckg[18]) );
  NAND2_X1 npu_inst_U142 ( .A1(npu_inst_n123), .A2(npu_inst_n120), .ZN(
        npu_inst_int_ckg[17]) );
  NAND2_X1 npu_inst_U141 ( .A1(npu_inst_n123), .A2(npu_inst_n121), .ZN(
        npu_inst_int_ckg[16]) );
  BUF_X1 npu_inst_U140 ( .A(ps_int_ifmaps_ptr[1]), .Z(npu_inst_n55) );
  BUF_X1 npu_inst_U139 ( .A(ps_int_ifmaps_ptr[0]), .Z(npu_inst_n53) );
  BUF_X1 npu_inst_U138 ( .A(ps_int_ifmaps_ptr[0]), .Z(npu_inst_n52) );
  BUF_X1 npu_inst_U137 ( .A(ps_int_ifmaps_ptr[0]), .Z(npu_inst_n51) );
  BUF_X1 npu_inst_U136 ( .A(ps_int_ifmaps_ptr[0]), .Z(npu_inst_n50) );
  BUF_X1 npu_inst_U135 ( .A(ps_int_ifmaps_ptr[0]), .Z(npu_inst_n49) );
  NAND2_X1 npu_inst_U134 ( .A1(npu_inst_n111), .A2(npu_inst_n120), .ZN(
        npu_inst_int_ckg[57]) );
  NAND2_X1 npu_inst_U133 ( .A1(npu_inst_n113), .A2(npu_inst_n110), .ZN(
        npu_inst_int_ckg[55]) );
  NAND2_X1 npu_inst_U132 ( .A1(npu_inst_n113), .A2(npu_inst_n112), .ZN(
        npu_inst_int_ckg[54]) );
  NAND2_X1 npu_inst_U131 ( .A1(npu_inst_n113), .A2(npu_inst_n117), .ZN(
        npu_inst_int_ckg[53]) );
  NAND2_X1 npu_inst_U130 ( .A1(npu_inst_n113), .A2(npu_inst_n114), .ZN(
        npu_inst_int_ckg[52]) );
  NAND2_X1 npu_inst_U129 ( .A1(npu_inst_n113), .A2(npu_inst_n118), .ZN(
        npu_inst_int_ckg[51]) );
  NAND2_X1 npu_inst_U128 ( .A1(npu_inst_n113), .A2(npu_inst_n119), .ZN(
        npu_inst_int_ckg[50]) );
  NAND2_X1 npu_inst_U127 ( .A1(npu_inst_n113), .A2(npu_inst_n120), .ZN(
        npu_inst_int_ckg[49]) );
  NAND2_X1 npu_inst_U126 ( .A1(npu_inst_n113), .A2(npu_inst_n121), .ZN(
        npu_inst_int_ckg[48]) );
  NAND2_X1 npu_inst_U125 ( .A1(npu_inst_n116), .A2(npu_inst_n110), .ZN(
        npu_inst_int_ckg[47]) );
  NAND2_X1 npu_inst_U124 ( .A1(npu_inst_n116), .A2(npu_inst_n112), .ZN(
        npu_inst_int_ckg[46]) );
  NAND2_X1 npu_inst_U123 ( .A1(npu_inst_n116), .A2(npu_inst_n117), .ZN(
        npu_inst_int_ckg[45]) );
  NAND2_X1 npu_inst_U122 ( .A1(npu_inst_n116), .A2(npu_inst_n114), .ZN(
        npu_inst_int_ckg[44]) );
  NAND2_X1 npu_inst_U121 ( .A1(npu_inst_n116), .A2(npu_inst_n118), .ZN(
        npu_inst_int_ckg[43]) );
  NAND2_X1 npu_inst_U120 ( .A1(npu_inst_n116), .A2(npu_inst_n119), .ZN(
        npu_inst_int_ckg[42]) );
  NAND2_X1 npu_inst_U119 ( .A1(npu_inst_n116), .A2(npu_inst_n120), .ZN(
        npu_inst_int_ckg[41]) );
  NAND2_X1 npu_inst_U118 ( .A1(npu_inst_n116), .A2(npu_inst_n121), .ZN(
        npu_inst_int_ckg[40]) );
  NAND2_X1 npu_inst_U117 ( .A1(npu_inst_n115), .A2(npu_inst_n110), .ZN(
        npu_inst_int_ckg[39]) );
  NAND2_X1 npu_inst_U116 ( .A1(npu_inst_n115), .A2(npu_inst_n112), .ZN(
        npu_inst_int_ckg[38]) );
  NAND2_X1 npu_inst_U115 ( .A1(npu_inst_n115), .A2(npu_inst_n117), .ZN(
        npu_inst_int_ckg[37]) );
  NAND2_X1 npu_inst_U114 ( .A1(npu_inst_n115), .A2(npu_inst_n114), .ZN(
        npu_inst_int_ckg[36]) );
  NAND2_X1 npu_inst_U113 ( .A1(npu_inst_n115), .A2(npu_inst_n118), .ZN(
        npu_inst_int_ckg[35]) );
  NAND2_X1 npu_inst_U112 ( .A1(npu_inst_n115), .A2(npu_inst_n119), .ZN(
        npu_inst_int_ckg[34]) );
  NAND2_X1 npu_inst_U111 ( .A1(npu_inst_n115), .A2(npu_inst_n120), .ZN(
        npu_inst_int_ckg[33]) );
  NAND2_X1 npu_inst_U110 ( .A1(npu_inst_n115), .A2(npu_inst_n121), .ZN(
        npu_inst_int_ckg[32]) );
  NAND2_X1 npu_inst_U109 ( .A1(npu_inst_n125), .A2(npu_inst_n112), .ZN(
        npu_inst_int_ckg[30]) );
  NAND2_X1 npu_inst_U108 ( .A1(npu_inst_n125), .A2(npu_inst_n117), .ZN(
        npu_inst_int_ckg[29]) );
  NAND2_X1 npu_inst_U107 ( .A1(npu_inst_n125), .A2(npu_inst_n114), .ZN(
        npu_inst_int_ckg[28]) );
  NAND2_X1 npu_inst_U106 ( .A1(npu_inst_n125), .A2(npu_inst_n119), .ZN(
        npu_inst_int_ckg[26]) );
  NAND2_X1 npu_inst_U105 ( .A1(npu_inst_n125), .A2(npu_inst_n120), .ZN(
        npu_inst_int_ckg[25]) );
  NAND2_X1 npu_inst_U104 ( .A1(npu_inst_n125), .A2(npu_inst_n121), .ZN(
        npu_inst_int_ckg[24]) );
  NAND2_X1 npu_inst_U103 ( .A1(npu_inst_n124), .A2(npu_inst_n110), .ZN(
        npu_inst_int_ckg[15]) );
  NAND2_X1 npu_inst_U102 ( .A1(npu_inst_n124), .A2(npu_inst_n112), .ZN(
        npu_inst_int_ckg[14]) );
  NAND2_X1 npu_inst_U101 ( .A1(npu_inst_n124), .A2(npu_inst_n117), .ZN(
        npu_inst_int_ckg[13]) );
  NAND2_X1 npu_inst_U100 ( .A1(npu_inst_n124), .A2(npu_inst_n114), .ZN(
        npu_inst_int_ckg[12]) );
  NAND2_X1 npu_inst_U99 ( .A1(npu_inst_n124), .A2(npu_inst_n118), .ZN(
        npu_inst_int_ckg[11]) );
  NAND2_X1 npu_inst_U98 ( .A1(npu_inst_n124), .A2(npu_inst_n119), .ZN(
        npu_inst_int_ckg[10]) );
  NAND2_X1 npu_inst_U97 ( .A1(npu_inst_n124), .A2(npu_inst_n120), .ZN(
        npu_inst_int_ckg[9]) );
  NAND2_X1 npu_inst_U96 ( .A1(npu_inst_n124), .A2(npu_inst_n121), .ZN(
        npu_inst_int_ckg[8]) );
  NAND2_X1 npu_inst_U95 ( .A1(npu_inst_n122), .A2(npu_inst_n110), .ZN(
        npu_inst_int_ckg[7]) );
  NAND2_X1 npu_inst_U94 ( .A1(npu_inst_n122), .A2(npu_inst_n112), .ZN(
        npu_inst_int_ckg[6]) );
  NAND2_X1 npu_inst_U93 ( .A1(npu_inst_n122), .A2(npu_inst_n117), .ZN(
        npu_inst_int_ckg[5]) );
  NAND2_X1 npu_inst_U92 ( .A1(npu_inst_n122), .A2(npu_inst_n114), .ZN(
        npu_inst_int_ckg[4]) );
  NAND2_X1 npu_inst_U91 ( .A1(npu_inst_n122), .A2(npu_inst_n118), .ZN(
        npu_inst_int_ckg[3]) );
  NAND2_X1 npu_inst_U90 ( .A1(npu_inst_n122), .A2(npu_inst_n119), .ZN(
        npu_inst_int_ckg[2]) );
  NAND2_X1 npu_inst_U89 ( .A1(npu_inst_n122), .A2(npu_inst_n120), .ZN(
        npu_inst_int_ckg[1]) );
  NAND2_X1 npu_inst_U88 ( .A1(npu_inst_n122), .A2(npu_inst_n121), .ZN(
        npu_inst_int_ckg[0]) );
  INV_X1 npu_inst_U87 ( .A(int_ckg_rmask[1]), .ZN(npu_inst_n113) );
  INV_X1 npu_inst_U86 ( .A(int_ckg_rmask[2]), .ZN(npu_inst_n116) );
  INV_X1 npu_inst_U85 ( .A(int_ckg_rmask[3]), .ZN(npu_inst_n115) );
  INV_X1 npu_inst_U84 ( .A(int_ckg_rmask[7]), .ZN(npu_inst_n122) );
  INV_X1 npu_inst_U83 ( .A(int_ckg_cmask[1]), .ZN(npu_inst_n112) );
  INV_X1 npu_inst_U82 ( .A(int_ckg_cmask[2]), .ZN(npu_inst_n117) );
  INV_X1 npu_inst_U81 ( .A(int_ckg_cmask[3]), .ZN(npu_inst_n114) );
  INV_X1 npu_inst_U80 ( .A(int_ckg_cmask[7]), .ZN(npu_inst_n121) );
  INV_X1 npu_inst_U79 ( .A(int_ckg_cmask[6]), .ZN(npu_inst_n120) );
  BUF_X1 npu_inst_U78 ( .A(npu_inst_n10), .Z(npu_inst_n2) );
  BUF_X1 npu_inst_U77 ( .A(npu_inst_n10), .Z(npu_inst_n1) );
  BUF_X1 npu_inst_U76 ( .A(npu_inst_n8), .Z(npu_inst_n7) );
  BUF_X1 npu_inst_U75 ( .A(npu_inst_n8), .Z(npu_inst_n6) );
  BUF_X1 npu_inst_U74 ( .A(npu_inst_n9), .Z(npu_inst_n5) );
  BUF_X1 npu_inst_U73 ( .A(npu_inst_n9), .Z(npu_inst_n4) );
  BUF_X1 npu_inst_U72 ( .A(npu_inst_n9), .Z(npu_inst_n3) );
  BUF_X2 npu_inst_U71 ( .A(npu_inst_n33), .Z(npu_inst_n42) );
  BUF_X2 npu_inst_U70 ( .A(npu_inst_n33), .Z(npu_inst_n41) );
  BUF_X2 npu_inst_U69 ( .A(npu_inst_n33), .Z(npu_inst_n40) );
  BUF_X2 npu_inst_U68 ( .A(npu_inst_n33), .Z(npu_inst_n39) );
  BUF_X2 npu_inst_U67 ( .A(npu_inst_n32), .Z(npu_inst_n38) );
  BUF_X2 npu_inst_U66 ( .A(npu_inst_n32), .Z(npu_inst_n37) );
  BUF_X2 npu_inst_U65 ( .A(npu_inst_n32), .Z(npu_inst_n36) );
  BUF_X2 npu_inst_U64 ( .A(npu_inst_n32), .Z(npu_inst_n35) );
  BUF_X2 npu_inst_U63 ( .A(npu_inst_n32), .Z(npu_inst_n34) );
  BUF_X1 npu_inst_U62 ( .A(npu_inst_n73), .Z(npu_inst_n64) );
  BUF_X1 npu_inst_U61 ( .A(npu_inst_n73), .Z(npu_inst_n63) );
  BUF_X1 npu_inst_U60 ( .A(npu_inst_n71), .Z(npu_inst_n70) );
  BUF_X1 npu_inst_U59 ( .A(npu_inst_n71), .Z(npu_inst_n69) );
  BUF_X1 npu_inst_U58 ( .A(npu_inst_n71), .Z(npu_inst_n68) );
  BUF_X1 npu_inst_U57 ( .A(npu_inst_n72), .Z(npu_inst_n67) );
  BUF_X1 npu_inst_U56 ( .A(npu_inst_n72), .Z(npu_inst_n66) );
  BUF_X1 npu_inst_U55 ( .A(npu_inst_n72), .Z(npu_inst_n65) );
  INV_X1 npu_inst_U54 ( .A(n63), .ZN(npu_inst_n119) );
  INV_X1 npu_inst_U53 ( .A(int_ckg_rmask[6]), .ZN(npu_inst_n124) );
  BUF_X1 npu_inst_U52 ( .A(npu_inst_n56), .Z(npu_inst_n62) );
  INV_X1 npu_inst_U51 ( .A(n64), .ZN(npu_inst_n123) );
  BUF_X1 npu_inst_U50 ( .A(npu_inst_n56), .Z(npu_inst_n61) );
  BUF_X1 npu_inst_U49 ( .A(npu_inst_n56), .Z(npu_inst_n60) );
  BUF_X1 npu_inst_U48 ( .A(npu_inst_n55), .Z(npu_inst_n59) );
  BUF_X1 npu_inst_U47 ( .A(npu_inst_n55), .Z(npu_inst_n58) );
  BUF_X1 npu_inst_U46 ( .A(npu_inst_n55), .Z(npu_inst_n57) );
  BUF_X1 npu_inst_U45 ( .A(n47), .Z(npu_inst_n103) );
  BUF_X1 npu_inst_U44 ( .A(n47), .Z(npu_inst_n102) );
  BUF_X1 npu_inst_U43 ( .A(npu_inst_n7), .Z(npu_inst_n31) );
  BUF_X1 npu_inst_U42 ( .A(npu_inst_n7), .Z(npu_inst_n30) );
  BUF_X1 npu_inst_U41 ( .A(npu_inst_n7), .Z(npu_inst_n29) );
  BUF_X1 npu_inst_U40 ( .A(npu_inst_n6), .Z(npu_inst_n28) );
  BUF_X1 npu_inst_U39 ( .A(npu_inst_n6), .Z(npu_inst_n27) );
  BUF_X1 npu_inst_U38 ( .A(npu_inst_n6), .Z(npu_inst_n26) );
  BUF_X1 npu_inst_U37 ( .A(npu_inst_n5), .Z(npu_inst_n25) );
  BUF_X1 npu_inst_U36 ( .A(npu_inst_n5), .Z(npu_inst_n24) );
  BUF_X1 npu_inst_U35 ( .A(npu_inst_n5), .Z(npu_inst_n23) );
  BUF_X1 npu_inst_U34 ( .A(npu_inst_n4), .Z(npu_inst_n22) );
  BUF_X1 npu_inst_U33 ( .A(npu_inst_n4), .Z(npu_inst_n21) );
  BUF_X1 npu_inst_U32 ( .A(npu_inst_n4), .Z(npu_inst_n20) );
  BUF_X1 npu_inst_U31 ( .A(npu_inst_n3), .Z(npu_inst_n19) );
  BUF_X1 npu_inst_U30 ( .A(npu_inst_n3), .Z(npu_inst_n18) );
  BUF_X1 npu_inst_U29 ( .A(npu_inst_n3), .Z(npu_inst_n17) );
  BUF_X1 npu_inst_U28 ( .A(npu_inst_n2), .Z(npu_inst_n16) );
  BUF_X1 npu_inst_U27 ( .A(npu_inst_n2), .Z(npu_inst_n15) );
  BUF_X1 npu_inst_U26 ( .A(npu_inst_n2), .Z(npu_inst_n14) );
  BUF_X1 npu_inst_U25 ( .A(npu_inst_n1), .Z(npu_inst_n13) );
  BUF_X1 npu_inst_U24 ( .A(npu_inst_n1), .Z(npu_inst_n12) );
  BUF_X1 npu_inst_U23 ( .A(npu_inst_n1), .Z(npu_inst_n11) );
  BUF_X1 npu_inst_U22 ( .A(npu_inst_n70), .Z(npu_inst_n89) );
  BUF_X1 npu_inst_U21 ( .A(npu_inst_n70), .Z(npu_inst_n88) );
  BUF_X1 npu_inst_U20 ( .A(npu_inst_n69), .Z(npu_inst_n87) );
  BUF_X1 npu_inst_U19 ( .A(npu_inst_n69), .Z(npu_inst_n86) );
  BUF_X1 npu_inst_U18 ( .A(npu_inst_n68), .Z(npu_inst_n85) );
  BUF_X1 npu_inst_U17 ( .A(npu_inst_n68), .Z(npu_inst_n84) );
  BUF_X1 npu_inst_U16 ( .A(npu_inst_n67), .Z(npu_inst_n83) );
  BUF_X1 npu_inst_U15 ( .A(npu_inst_n67), .Z(npu_inst_n82) );
  BUF_X1 npu_inst_U14 ( .A(npu_inst_n66), .Z(npu_inst_n81) );
  BUF_X1 npu_inst_U13 ( .A(npu_inst_n66), .Z(npu_inst_n80) );
  BUF_X1 npu_inst_U12 ( .A(npu_inst_n65), .Z(npu_inst_n79) );
  BUF_X1 npu_inst_U11 ( .A(npu_inst_n65), .Z(npu_inst_n78) );
  BUF_X1 npu_inst_U10 ( .A(npu_inst_n64), .Z(npu_inst_n77) );
  BUF_X1 npu_inst_U9 ( .A(npu_inst_n64), .Z(npu_inst_n76) );
  BUF_X1 npu_inst_U8 ( .A(npu_inst_n63), .Z(npu_inst_n75) );
  BUF_X1 npu_inst_U7 ( .A(npu_inst_n63), .Z(npu_inst_n74) );
  BUF_X1 npu_inst_U6 ( .A(npu_inst_n103), .Z(npu_inst_n109) );
  BUF_X1 npu_inst_U5 ( .A(npu_inst_n103), .Z(npu_inst_n108) );
  BUF_X1 npu_inst_U4 ( .A(npu_inst_n103), .Z(npu_inst_n107) );
  BUF_X1 npu_inst_U3 ( .A(npu_inst_n102), .Z(npu_inst_n106) );
  BUF_X1 npu_inst_U2 ( .A(npu_inst_n102), .Z(npu_inst_n105) );
  BUF_X1 npu_inst_U1 ( .A(npu_inst_n102), .Z(npu_inst_n104) );
  MUX2_X1 npu_inst_pe_1_0_0_U151 ( .A(npu_inst_pe_1_0_0_n29), .B(
        npu_inst_pe_1_0_0_n24), .S(npu_inst_pe_1_0_0_n5), .Z(
        npu_inst_pe_1_0_0_N93) );
  MUX2_X1 npu_inst_pe_1_0_0_U150 ( .A(npu_inst_pe_1_0_0_n28), .B(
        npu_inst_pe_1_0_0_n25), .S(npu_inst_n62), .Z(npu_inst_pe_1_0_0_n29) );
  MUX2_X1 npu_inst_pe_1_0_0_U149 ( .A(npu_inst_pe_1_0_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_0_n2), .Z(
        npu_inst_pe_1_0_0_n28) );
  MUX2_X1 npu_inst_pe_1_0_0_U148 ( .A(npu_inst_pe_1_0_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_0_n2), .Z(
        npu_inst_pe_1_0_0_n25) );
  MUX2_X1 npu_inst_pe_1_0_0_U147 ( .A(npu_inst_pe_1_0_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_0_n2), .Z(
        npu_inst_pe_1_0_0_n24) );
  MUX2_X1 npu_inst_pe_1_0_0_U146 ( .A(npu_inst_pe_1_0_0_n23), .B(
        npu_inst_pe_1_0_0_n20), .S(npu_inst_pe_1_0_0_n5), .Z(
        npu_inst_pe_1_0_0_N94) );
  MUX2_X1 npu_inst_pe_1_0_0_U145 ( .A(npu_inst_pe_1_0_0_n22), .B(
        npu_inst_pe_1_0_0_n21), .S(npu_inst_n62), .Z(npu_inst_pe_1_0_0_n23) );
  MUX2_X1 npu_inst_pe_1_0_0_U144 ( .A(npu_inst_pe_1_0_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_0_n2), .Z(
        npu_inst_pe_1_0_0_n22) );
  MUX2_X1 npu_inst_pe_1_0_0_U143 ( .A(npu_inst_pe_1_0_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_0_n2), .Z(
        npu_inst_pe_1_0_0_n21) );
  MUX2_X1 npu_inst_pe_1_0_0_U142 ( .A(npu_inst_pe_1_0_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_0_n2), .Z(
        npu_inst_pe_1_0_0_n20) );
  MUX2_X1 npu_inst_pe_1_0_0_U141 ( .A(npu_inst_pe_1_0_0_n19), .B(
        npu_inst_pe_1_0_0_n16), .S(npu_inst_pe_1_0_0_n5), .Z(
        npu_inst_pe_1_0_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_0_0_U140 ( .A(npu_inst_pe_1_0_0_n18), .B(
        npu_inst_pe_1_0_0_n17), .S(npu_inst_n62), .Z(npu_inst_pe_1_0_0_n19) );
  MUX2_X1 npu_inst_pe_1_0_0_U139 ( .A(npu_inst_pe_1_0_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_0_n2), .Z(
        npu_inst_pe_1_0_0_n18) );
  MUX2_X1 npu_inst_pe_1_0_0_U138 ( .A(npu_inst_pe_1_0_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_0_n2), .Z(
        npu_inst_pe_1_0_0_n17) );
  MUX2_X1 npu_inst_pe_1_0_0_U137 ( .A(npu_inst_pe_1_0_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_0_n2), .Z(
        npu_inst_pe_1_0_0_n16) );
  MUX2_X1 npu_inst_pe_1_0_0_U136 ( .A(npu_inst_pe_1_0_0_n15), .B(
        npu_inst_pe_1_0_0_n12), .S(npu_inst_pe_1_0_0_n5), .Z(
        npu_inst_pe_1_0_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_0_0_U135 ( .A(npu_inst_pe_1_0_0_n14), .B(
        npu_inst_pe_1_0_0_n13), .S(npu_inst_n62), .Z(npu_inst_pe_1_0_0_n15) );
  MUX2_X1 npu_inst_pe_1_0_0_U134 ( .A(npu_inst_pe_1_0_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_0_n2), .Z(
        npu_inst_pe_1_0_0_n14) );
  MUX2_X1 npu_inst_pe_1_0_0_U133 ( .A(npu_inst_pe_1_0_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_0_n2), .Z(
        npu_inst_pe_1_0_0_n13) );
  MUX2_X1 npu_inst_pe_1_0_0_U132 ( .A(npu_inst_pe_1_0_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_0_n2), .Z(
        npu_inst_pe_1_0_0_n12) );
  XOR2_X1 npu_inst_pe_1_0_0_U131 ( .A(npu_inst_pe_1_0_0_int_data_0_), .B(
        int_o_data_npu[56]), .Z(npu_inst_pe_1_0_0_N73) );
  AND2_X1 npu_inst_pe_1_0_0_U130 ( .A1(int_o_data_npu[56]), .A2(
        npu_inst_pe_1_0_0_int_data_0_), .ZN(npu_inst_pe_1_0_0_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_0_U129 ( .A(int_o_data_npu[56]), .B(
        npu_inst_pe_1_0_0_n10), .ZN(npu_inst_pe_1_0_0_N65) );
  OR2_X1 npu_inst_pe_1_0_0_U128 ( .A1(npu_inst_pe_1_0_0_n10), .A2(
        int_o_data_npu[56]), .ZN(npu_inst_pe_1_0_0_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_0_U127 ( .A(int_o_data_npu[58]), .B(
        npu_inst_pe_1_0_0_add_79_carry_2_), .Z(npu_inst_pe_1_0_0_N75) );
  AND2_X1 npu_inst_pe_1_0_0_U126 ( .A1(npu_inst_pe_1_0_0_add_79_carry_2_), 
        .A2(int_o_data_npu[58]), .ZN(npu_inst_pe_1_0_0_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_0_U125 ( .A(int_o_data_npu[59]), .B(
        npu_inst_pe_1_0_0_add_79_carry_3_), .Z(npu_inst_pe_1_0_0_N76) );
  AND2_X1 npu_inst_pe_1_0_0_U124 ( .A1(npu_inst_pe_1_0_0_add_79_carry_3_), 
        .A2(int_o_data_npu[59]), .ZN(npu_inst_pe_1_0_0_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_0_U123 ( .A(int_o_data_npu[60]), .B(
        npu_inst_pe_1_0_0_add_79_carry_4_), .Z(npu_inst_pe_1_0_0_N77) );
  AND2_X1 npu_inst_pe_1_0_0_U122 ( .A1(npu_inst_pe_1_0_0_add_79_carry_4_), 
        .A2(int_o_data_npu[60]), .ZN(npu_inst_pe_1_0_0_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_0_U121 ( .A(int_o_data_npu[61]), .B(
        npu_inst_pe_1_0_0_add_79_carry_5_), .Z(npu_inst_pe_1_0_0_N78) );
  AND2_X1 npu_inst_pe_1_0_0_U120 ( .A1(npu_inst_pe_1_0_0_add_79_carry_5_), 
        .A2(int_o_data_npu[61]), .ZN(npu_inst_pe_1_0_0_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_0_U119 ( .A(int_o_data_npu[62]), .B(
        npu_inst_pe_1_0_0_add_79_carry_6_), .Z(npu_inst_pe_1_0_0_N79) );
  AND2_X1 npu_inst_pe_1_0_0_U118 ( .A1(npu_inst_pe_1_0_0_add_79_carry_6_), 
        .A2(int_o_data_npu[62]), .ZN(npu_inst_pe_1_0_0_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_0_U117 ( .A(int_o_data_npu[63]), .B(
        npu_inst_pe_1_0_0_add_79_carry_7_), .Z(npu_inst_pe_1_0_0_N80) );
  XNOR2_X1 npu_inst_pe_1_0_0_U116 ( .A(npu_inst_pe_1_0_0_sub_77_carry_2_), .B(
        int_o_data_npu[58]), .ZN(npu_inst_pe_1_0_0_N67) );
  OR2_X1 npu_inst_pe_1_0_0_U115 ( .A1(int_o_data_npu[58]), .A2(
        npu_inst_pe_1_0_0_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_0_0_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_0_U114 ( .A(npu_inst_pe_1_0_0_sub_77_carry_3_), .B(
        int_o_data_npu[59]), .ZN(npu_inst_pe_1_0_0_N68) );
  OR2_X1 npu_inst_pe_1_0_0_U113 ( .A1(int_o_data_npu[59]), .A2(
        npu_inst_pe_1_0_0_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_0_0_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_0_U112 ( .A(npu_inst_pe_1_0_0_sub_77_carry_4_), .B(
        int_o_data_npu[60]), .ZN(npu_inst_pe_1_0_0_N69) );
  OR2_X1 npu_inst_pe_1_0_0_U111 ( .A1(int_o_data_npu[60]), .A2(
        npu_inst_pe_1_0_0_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_0_0_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_0_U110 ( .A(npu_inst_pe_1_0_0_sub_77_carry_5_), .B(
        int_o_data_npu[61]), .ZN(npu_inst_pe_1_0_0_N70) );
  OR2_X1 npu_inst_pe_1_0_0_U109 ( .A1(int_o_data_npu[61]), .A2(
        npu_inst_pe_1_0_0_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_0_0_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_0_U108 ( .A(npu_inst_pe_1_0_0_sub_77_carry_6_), .B(
        int_o_data_npu[62]), .ZN(npu_inst_pe_1_0_0_N71) );
  OR2_X1 npu_inst_pe_1_0_0_U107 ( .A1(int_o_data_npu[62]), .A2(
        npu_inst_pe_1_0_0_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_0_0_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_0_U106 ( .A(int_o_data_npu[63]), .B(
        npu_inst_pe_1_0_0_sub_77_carry_7_), .ZN(npu_inst_pe_1_0_0_N72) );
  INV_X1 npu_inst_pe_1_0_0_U105 ( .A(npu_inst_n62), .ZN(npu_inst_pe_1_0_0_n4)
         );
  INV_X1 npu_inst_pe_1_0_0_U104 ( .A(npu_inst_n39), .ZN(npu_inst_pe_1_0_0_n1)
         );
  AOI22_X1 npu_inst_pe_1_0_0_U103 ( .A1(npu_inst_pe_1_0_0_n38), .A2(
        npu_inst_int_data_y_1__0__1_), .B1(npu_inst_pe_1_0_0_n111), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_0_n39) );
  INV_X1 npu_inst_pe_1_0_0_U102 ( .A(npu_inst_pe_1_0_0_n39), .ZN(
        npu_inst_pe_1_0_0_n104) );
  NOR3_X1 npu_inst_pe_1_0_0_U99 ( .A1(npu_inst_pe_1_0_0_n26), .A2(npu_inst_n39), .A3(npu_inst_int_ckg[63]), .ZN(npu_inst_pe_1_0_0_n85) );
  OR2_X1 npu_inst_pe_1_0_0_U98 ( .A1(npu_inst_pe_1_0_0_n85), .A2(npu_inst_n8), 
        .ZN(npu_inst_pe_1_0_0_N84) );
  NAND2_X1 npu_inst_pe_1_0_0_U97 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_0_n60), .ZN(npu_inst_pe_1_0_0_n74) );
  OAI21_X1 npu_inst_pe_1_0_0_U96 ( .B1(npu_inst_pe_1_0_0_n63), .B2(
        npu_inst_pe_1_0_0_n60), .A(npu_inst_pe_1_0_0_n74), .ZN(
        npu_inst_pe_1_0_0_n97) );
  NAND2_X1 npu_inst_pe_1_0_0_U95 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_0_n60), .ZN(npu_inst_pe_1_0_0_n73) );
  OAI21_X1 npu_inst_pe_1_0_0_U94 ( .B1(npu_inst_pe_1_0_0_n61), .B2(
        npu_inst_pe_1_0_0_n60), .A(npu_inst_pe_1_0_0_n73), .ZN(
        npu_inst_pe_1_0_0_n96) );
  NAND2_X1 npu_inst_pe_1_0_0_U93 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_0_n56), .ZN(npu_inst_pe_1_0_0_n72) );
  OAI21_X1 npu_inst_pe_1_0_0_U92 ( .B1(npu_inst_pe_1_0_0_n63), .B2(
        npu_inst_pe_1_0_0_n56), .A(npu_inst_pe_1_0_0_n72), .ZN(
        npu_inst_pe_1_0_0_n95) );
  NAND2_X1 npu_inst_pe_1_0_0_U91 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_0_n56), .ZN(npu_inst_pe_1_0_0_n71) );
  OAI21_X1 npu_inst_pe_1_0_0_U90 ( .B1(npu_inst_pe_1_0_0_n61), .B2(
        npu_inst_pe_1_0_0_n56), .A(npu_inst_pe_1_0_0_n71), .ZN(
        npu_inst_pe_1_0_0_n94) );
  NAND2_X1 npu_inst_pe_1_0_0_U89 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_0_n52), .ZN(npu_inst_pe_1_0_0_n70) );
  OAI21_X1 npu_inst_pe_1_0_0_U88 ( .B1(npu_inst_pe_1_0_0_n63), .B2(
        npu_inst_pe_1_0_0_n52), .A(npu_inst_pe_1_0_0_n70), .ZN(
        npu_inst_pe_1_0_0_n93) );
  NAND2_X1 npu_inst_pe_1_0_0_U87 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_0_n52), .ZN(npu_inst_pe_1_0_0_n69) );
  OAI21_X1 npu_inst_pe_1_0_0_U86 ( .B1(npu_inst_pe_1_0_0_n61), .B2(
        npu_inst_pe_1_0_0_n52), .A(npu_inst_pe_1_0_0_n69), .ZN(
        npu_inst_pe_1_0_0_n92) );
  NAND2_X1 npu_inst_pe_1_0_0_U85 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_0_n48), .ZN(npu_inst_pe_1_0_0_n68) );
  OAI21_X1 npu_inst_pe_1_0_0_U84 ( .B1(npu_inst_pe_1_0_0_n63), .B2(
        npu_inst_pe_1_0_0_n48), .A(npu_inst_pe_1_0_0_n68), .ZN(
        npu_inst_pe_1_0_0_n91) );
  NAND2_X1 npu_inst_pe_1_0_0_U83 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_0_n48), .ZN(npu_inst_pe_1_0_0_n67) );
  OAI21_X1 npu_inst_pe_1_0_0_U82 ( .B1(npu_inst_pe_1_0_0_n61), .B2(
        npu_inst_pe_1_0_0_n48), .A(npu_inst_pe_1_0_0_n67), .ZN(
        npu_inst_pe_1_0_0_n90) );
  NAND2_X1 npu_inst_pe_1_0_0_U81 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_0_n44), .ZN(npu_inst_pe_1_0_0_n66) );
  OAI21_X1 npu_inst_pe_1_0_0_U80 ( .B1(npu_inst_pe_1_0_0_n63), .B2(
        npu_inst_pe_1_0_0_n44), .A(npu_inst_pe_1_0_0_n66), .ZN(
        npu_inst_pe_1_0_0_n89) );
  NAND2_X1 npu_inst_pe_1_0_0_U79 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_0_n44), .ZN(npu_inst_pe_1_0_0_n65) );
  OAI21_X1 npu_inst_pe_1_0_0_U78 ( .B1(npu_inst_pe_1_0_0_n61), .B2(
        npu_inst_pe_1_0_0_n44), .A(npu_inst_pe_1_0_0_n65), .ZN(
        npu_inst_pe_1_0_0_n88) );
  NAND2_X1 npu_inst_pe_1_0_0_U77 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_0_n40), .ZN(npu_inst_pe_1_0_0_n64) );
  OAI21_X1 npu_inst_pe_1_0_0_U76 ( .B1(npu_inst_pe_1_0_0_n63), .B2(
        npu_inst_pe_1_0_0_n40), .A(npu_inst_pe_1_0_0_n64), .ZN(
        npu_inst_pe_1_0_0_n87) );
  NAND2_X1 npu_inst_pe_1_0_0_U75 ( .A1(npu_inst_pe_1_0_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_0_n40), .ZN(npu_inst_pe_1_0_0_n62) );
  OAI21_X1 npu_inst_pe_1_0_0_U74 ( .B1(npu_inst_pe_1_0_0_n61), .B2(
        npu_inst_pe_1_0_0_n40), .A(npu_inst_pe_1_0_0_n62), .ZN(
        npu_inst_pe_1_0_0_n86) );
  AOI22_X1 npu_inst_pe_1_0_0_U73 ( .A1(npu_inst_pe_1_0_0_n38), .A2(
        npu_inst_int_data_y_1__0__0_), .B1(npu_inst_pe_1_0_0_n111), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_0_n37) );
  INV_X1 npu_inst_pe_1_0_0_U72 ( .A(npu_inst_pe_1_0_0_n37), .ZN(
        npu_inst_pe_1_0_0_n110) );
  AOI22_X1 npu_inst_pe_1_0_0_U71 ( .A1(npu_inst_int_data_y_1__0__1_), .A2(
        npu_inst_pe_1_0_0_n58), .B1(npu_inst_pe_1_0_0_n116), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_0_n59) );
  INV_X1 npu_inst_pe_1_0_0_U70 ( .A(npu_inst_pe_1_0_0_n59), .ZN(
        npu_inst_pe_1_0_0_n99) );
  AOI22_X1 npu_inst_pe_1_0_0_U69 ( .A1(npu_inst_int_data_y_1__0__0_), .A2(
        npu_inst_pe_1_0_0_n58), .B1(npu_inst_pe_1_0_0_n116), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_0_n57) );
  INV_X1 npu_inst_pe_1_0_0_U68 ( .A(npu_inst_pe_1_0_0_n57), .ZN(
        npu_inst_pe_1_0_0_n105) );
  AOI22_X1 npu_inst_pe_1_0_0_U67 ( .A1(npu_inst_int_data_y_1__0__1_), .A2(
        npu_inst_pe_1_0_0_n54), .B1(npu_inst_pe_1_0_0_n115), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_0_n55) );
  INV_X1 npu_inst_pe_1_0_0_U66 ( .A(npu_inst_pe_1_0_0_n55), .ZN(
        npu_inst_pe_1_0_0_n100) );
  AOI22_X1 npu_inst_pe_1_0_0_U65 ( .A1(npu_inst_int_data_y_1__0__0_), .A2(
        npu_inst_pe_1_0_0_n54), .B1(npu_inst_pe_1_0_0_n115), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_0_n53) );
  INV_X1 npu_inst_pe_1_0_0_U64 ( .A(npu_inst_pe_1_0_0_n53), .ZN(
        npu_inst_pe_1_0_0_n106) );
  AOI22_X1 npu_inst_pe_1_0_0_U63 ( .A1(npu_inst_int_data_y_1__0__1_), .A2(
        npu_inst_pe_1_0_0_n50), .B1(npu_inst_pe_1_0_0_n114), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_0_n51) );
  INV_X1 npu_inst_pe_1_0_0_U62 ( .A(npu_inst_pe_1_0_0_n51), .ZN(
        npu_inst_pe_1_0_0_n101) );
  AOI22_X1 npu_inst_pe_1_0_0_U61 ( .A1(npu_inst_int_data_y_1__0__0_), .A2(
        npu_inst_pe_1_0_0_n50), .B1(npu_inst_pe_1_0_0_n114), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_0_n49) );
  INV_X1 npu_inst_pe_1_0_0_U60 ( .A(npu_inst_pe_1_0_0_n49), .ZN(
        npu_inst_pe_1_0_0_n107) );
  AOI22_X1 npu_inst_pe_1_0_0_U59 ( .A1(npu_inst_int_data_y_1__0__1_), .A2(
        npu_inst_pe_1_0_0_n46), .B1(npu_inst_pe_1_0_0_n113), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_0_n47) );
  INV_X1 npu_inst_pe_1_0_0_U58 ( .A(npu_inst_pe_1_0_0_n47), .ZN(
        npu_inst_pe_1_0_0_n102) );
  AOI22_X1 npu_inst_pe_1_0_0_U57 ( .A1(npu_inst_int_data_y_1__0__0_), .A2(
        npu_inst_pe_1_0_0_n46), .B1(npu_inst_pe_1_0_0_n113), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_0_n45) );
  INV_X1 npu_inst_pe_1_0_0_U56 ( .A(npu_inst_pe_1_0_0_n45), .ZN(
        npu_inst_pe_1_0_0_n108) );
  AOI22_X1 npu_inst_pe_1_0_0_U55 ( .A1(npu_inst_int_data_y_1__0__1_), .A2(
        npu_inst_pe_1_0_0_n42), .B1(npu_inst_pe_1_0_0_n112), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_0_n43) );
  INV_X1 npu_inst_pe_1_0_0_U54 ( .A(npu_inst_pe_1_0_0_n43), .ZN(
        npu_inst_pe_1_0_0_n103) );
  AOI22_X1 npu_inst_pe_1_0_0_U53 ( .A1(npu_inst_int_data_y_1__0__0_), .A2(
        npu_inst_pe_1_0_0_n42), .B1(npu_inst_pe_1_0_0_n112), .B2(
        npu_inst_pe_1_0_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_0_n41) );
  INV_X1 npu_inst_pe_1_0_0_U52 ( .A(npu_inst_pe_1_0_0_n41), .ZN(
        npu_inst_pe_1_0_0_n109) );
  AOI222_X1 npu_inst_pe_1_0_0_U51 ( .A1(npu_inst_int_data_res_1__0__0_), .A2(
        npu_inst_n8), .B1(npu_inst_pe_1_0_0_N73), .B2(npu_inst_pe_1_0_0_n76), 
        .C1(npu_inst_pe_1_0_0_N65), .C2(npu_inst_pe_1_0_0_n77), .ZN(
        npu_inst_pe_1_0_0_n84) );
  INV_X1 npu_inst_pe_1_0_0_U50 ( .A(npu_inst_pe_1_0_0_n84), .ZN(
        npu_inst_pe_1_0_0_n98) );
  AOI222_X1 npu_inst_pe_1_0_0_U49 ( .A1(npu_inst_n8), .A2(
        npu_inst_int_data_res_1__0__7_), .B1(npu_inst_pe_1_0_0_N80), .B2(
        npu_inst_pe_1_0_0_n76), .C1(npu_inst_pe_1_0_0_N72), .C2(
        npu_inst_pe_1_0_0_n77), .ZN(npu_inst_pe_1_0_0_n75) );
  INV_X1 npu_inst_pe_1_0_0_U48 ( .A(npu_inst_pe_1_0_0_n75), .ZN(
        npu_inst_pe_1_0_0_n30) );
  AOI222_X1 npu_inst_pe_1_0_0_U47 ( .A1(npu_inst_int_data_res_1__0__1_), .A2(
        npu_inst_n8), .B1(npu_inst_pe_1_0_0_N74), .B2(npu_inst_pe_1_0_0_n76), 
        .C1(npu_inst_pe_1_0_0_N66), .C2(npu_inst_pe_1_0_0_n77), .ZN(
        npu_inst_pe_1_0_0_n83) );
  INV_X1 npu_inst_pe_1_0_0_U46 ( .A(npu_inst_pe_1_0_0_n83), .ZN(
        npu_inst_pe_1_0_0_n36) );
  AOI222_X1 npu_inst_pe_1_0_0_U45 ( .A1(npu_inst_int_data_res_1__0__2_), .A2(
        npu_inst_n8), .B1(npu_inst_pe_1_0_0_N75), .B2(npu_inst_pe_1_0_0_n76), 
        .C1(npu_inst_pe_1_0_0_N67), .C2(npu_inst_pe_1_0_0_n77), .ZN(
        npu_inst_pe_1_0_0_n82) );
  INV_X1 npu_inst_pe_1_0_0_U44 ( .A(npu_inst_pe_1_0_0_n82), .ZN(
        npu_inst_pe_1_0_0_n35) );
  AOI222_X1 npu_inst_pe_1_0_0_U43 ( .A1(npu_inst_int_data_res_1__0__3_), .A2(
        npu_inst_n8), .B1(npu_inst_pe_1_0_0_N76), .B2(npu_inst_pe_1_0_0_n76), 
        .C1(npu_inst_pe_1_0_0_N68), .C2(npu_inst_pe_1_0_0_n77), .ZN(
        npu_inst_pe_1_0_0_n81) );
  INV_X1 npu_inst_pe_1_0_0_U42 ( .A(npu_inst_pe_1_0_0_n81), .ZN(
        npu_inst_pe_1_0_0_n34) );
  AOI222_X1 npu_inst_pe_1_0_0_U41 ( .A1(npu_inst_int_data_res_1__0__4_), .A2(
        npu_inst_n8), .B1(npu_inst_pe_1_0_0_N77), .B2(npu_inst_pe_1_0_0_n76), 
        .C1(npu_inst_pe_1_0_0_N69), .C2(npu_inst_pe_1_0_0_n77), .ZN(
        npu_inst_pe_1_0_0_n80) );
  INV_X1 npu_inst_pe_1_0_0_U40 ( .A(npu_inst_pe_1_0_0_n80), .ZN(
        npu_inst_pe_1_0_0_n33) );
  AOI222_X1 npu_inst_pe_1_0_0_U39 ( .A1(npu_inst_int_data_res_1__0__5_), .A2(
        npu_inst_n8), .B1(npu_inst_pe_1_0_0_N78), .B2(npu_inst_pe_1_0_0_n76), 
        .C1(npu_inst_pe_1_0_0_N70), .C2(npu_inst_pe_1_0_0_n77), .ZN(
        npu_inst_pe_1_0_0_n79) );
  INV_X1 npu_inst_pe_1_0_0_U38 ( .A(npu_inst_pe_1_0_0_n79), .ZN(
        npu_inst_pe_1_0_0_n32) );
  AND2_X1 npu_inst_pe_1_0_0_U37 ( .A1(npu_inst_pe_1_0_0_o_data_h_1_), .A2(
        npu_inst_pe_1_0_0_int_q_weight_1_), .ZN(npu_inst_pe_1_0_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_0_U36 ( .A1(npu_inst_pe_1_0_0_o_data_h_0_), .A2(
        npu_inst_pe_1_0_0_int_q_weight_1_), .ZN(npu_inst_pe_1_0_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_0_0_U35 ( .A(npu_inst_pe_1_0_0_int_data_1_), .ZN(
        npu_inst_pe_1_0_0_n11) );
  AOI222_X1 npu_inst_pe_1_0_0_U34 ( .A1(npu_inst_int_data_res_1__0__6_), .A2(
        npu_inst_n8), .B1(npu_inst_pe_1_0_0_N79), .B2(npu_inst_pe_1_0_0_n76), 
        .C1(npu_inst_pe_1_0_0_N71), .C2(npu_inst_pe_1_0_0_n77), .ZN(
        npu_inst_pe_1_0_0_n78) );
  INV_X1 npu_inst_pe_1_0_0_U33 ( .A(npu_inst_pe_1_0_0_n78), .ZN(
        npu_inst_pe_1_0_0_n31) );
  AND2_X1 npu_inst_pe_1_0_0_U32 ( .A1(npu_inst_pe_1_0_0_N93), .A2(npu_inst_n39), .ZN(npu_inst_pe_1_0_0_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_0_U31 ( .A1(npu_inst_n39), .A2(npu_inst_pe_1_0_0_N94), .ZN(npu_inst_pe_1_0_0_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_0_U30 ( .A1(npu_inst_n39), .A2(
        npu_inst_int_data_y_1__0__1_), .B1(npu_inst_pe_1_0_0_n1), .B2(
        npu_inst_int_data_x_0__1__1_), .ZN(npu_inst_pe_1_0_0_n63) );
  AOI22_X1 npu_inst_pe_1_0_0_U29 ( .A1(npu_inst_n39), .A2(
        npu_inst_int_data_y_1__0__0_), .B1(npu_inst_pe_1_0_0_n1), .B2(
        npu_inst_int_data_x_0__1__0_), .ZN(npu_inst_pe_1_0_0_n61) );
  INV_X1 npu_inst_pe_1_0_0_U28 ( .A(npu_inst_pe_1_0_0_int_data_0_), .ZN(
        npu_inst_pe_1_0_0_n10) );
  INV_X1 npu_inst_pe_1_0_0_U27 ( .A(npu_inst_n54), .ZN(npu_inst_pe_1_0_0_n3)
         );
  OR3_X1 npu_inst_pe_1_0_0_U26 ( .A1(npu_inst_n62), .A2(npu_inst_pe_1_0_0_n5), 
        .A3(npu_inst_pe_1_0_0_n3), .ZN(npu_inst_pe_1_0_0_n56) );
  OR3_X1 npu_inst_pe_1_0_0_U25 ( .A1(npu_inst_pe_1_0_0_n3), .A2(
        npu_inst_pe_1_0_0_n5), .A3(npu_inst_pe_1_0_0_n4), .ZN(
        npu_inst_pe_1_0_0_n48) );
  INV_X1 npu_inst_pe_1_0_0_U24 ( .A(npu_inst_pe_1_0_0_n3), .ZN(
        npu_inst_pe_1_0_0_n2) );
  OR3_X1 npu_inst_pe_1_0_0_U23 ( .A1(npu_inst_pe_1_0_0_n2), .A2(
        npu_inst_pe_1_0_0_n5), .A3(npu_inst_pe_1_0_0_n4), .ZN(
        npu_inst_pe_1_0_0_n52) );
  OR3_X1 npu_inst_pe_1_0_0_U22 ( .A1(npu_inst_n62), .A2(npu_inst_pe_1_0_0_n5), 
        .A3(npu_inst_pe_1_0_0_n2), .ZN(npu_inst_pe_1_0_0_n60) );
  NOR2_X1 npu_inst_pe_1_0_0_U21 ( .A1(npu_inst_pe_1_0_0_n60), .A2(
        npu_inst_pe_1_0_0_n1), .ZN(npu_inst_pe_1_0_0_n58) );
  NOR2_X1 npu_inst_pe_1_0_0_U20 ( .A1(npu_inst_pe_1_0_0_n56), .A2(
        npu_inst_pe_1_0_0_n1), .ZN(npu_inst_pe_1_0_0_n54) );
  NOR2_X1 npu_inst_pe_1_0_0_U19 ( .A1(npu_inst_pe_1_0_0_n52), .A2(
        npu_inst_pe_1_0_0_n1), .ZN(npu_inst_pe_1_0_0_n50) );
  NOR2_X1 npu_inst_pe_1_0_0_U18 ( .A1(npu_inst_pe_1_0_0_n48), .A2(
        npu_inst_pe_1_0_0_n1), .ZN(npu_inst_pe_1_0_0_n46) );
  NOR2_X1 npu_inst_pe_1_0_0_U17 ( .A1(npu_inst_pe_1_0_0_n40), .A2(
        npu_inst_pe_1_0_0_n1), .ZN(npu_inst_pe_1_0_0_n38) );
  NOR2_X1 npu_inst_pe_1_0_0_U16 ( .A1(npu_inst_pe_1_0_0_n44), .A2(
        npu_inst_pe_1_0_0_n1), .ZN(npu_inst_pe_1_0_0_n42) );
  BUF_X1 npu_inst_pe_1_0_0_U15 ( .A(npu_inst_n89), .Z(npu_inst_pe_1_0_0_n5) );
  INV_X1 npu_inst_pe_1_0_0_U14 ( .A(npu_inst_n109), .ZN(npu_inst_pe_1_0_0_n9)
         );
  INV_X1 npu_inst_pe_1_0_0_U13 ( .A(npu_inst_pe_1_0_0_n38), .ZN(
        npu_inst_pe_1_0_0_n111) );
  INV_X1 npu_inst_pe_1_0_0_U12 ( .A(npu_inst_pe_1_0_0_n58), .ZN(
        npu_inst_pe_1_0_0_n116) );
  INV_X1 npu_inst_pe_1_0_0_U11 ( .A(npu_inst_pe_1_0_0_n54), .ZN(
        npu_inst_pe_1_0_0_n115) );
  INV_X1 npu_inst_pe_1_0_0_U10 ( .A(npu_inst_pe_1_0_0_n50), .ZN(
        npu_inst_pe_1_0_0_n114) );
  INV_X1 npu_inst_pe_1_0_0_U9 ( .A(npu_inst_pe_1_0_0_n46), .ZN(
        npu_inst_pe_1_0_0_n113) );
  INV_X1 npu_inst_pe_1_0_0_U8 ( .A(npu_inst_pe_1_0_0_n42), .ZN(
        npu_inst_pe_1_0_0_n112) );
  BUF_X1 npu_inst_pe_1_0_0_U7 ( .A(npu_inst_pe_1_0_0_n9), .Z(
        npu_inst_pe_1_0_0_n8) );
  BUF_X1 npu_inst_pe_1_0_0_U6 ( .A(npu_inst_pe_1_0_0_n9), .Z(
        npu_inst_pe_1_0_0_n7) );
  BUF_X1 npu_inst_pe_1_0_0_U5 ( .A(npu_inst_pe_1_0_0_n9), .Z(
        npu_inst_pe_1_0_0_n6) );
  NOR2_X1 npu_inst_pe_1_0_0_U4 ( .A1(npu_inst_pe_1_0_0_int_q_weight_0_), .A2(
        npu_inst_n8), .ZN(npu_inst_pe_1_0_0_n76) );
  NOR2_X1 npu_inst_pe_1_0_0_U3 ( .A1(npu_inst_pe_1_0_0_n27), .A2(npu_inst_n8), 
        .ZN(npu_inst_pe_1_0_0_n77) );
  FA_X1 npu_inst_pe_1_0_0_sub_77_U2_1 ( .A(int_o_data_npu[57]), .B(
        npu_inst_pe_1_0_0_n11), .CI(npu_inst_pe_1_0_0_sub_77_carry_1_), .CO(
        npu_inst_pe_1_0_0_sub_77_carry_2_), .S(npu_inst_pe_1_0_0_N66) );
  FA_X1 npu_inst_pe_1_0_0_add_79_U1_1 ( .A(int_o_data_npu[57]), .B(
        npu_inst_pe_1_0_0_int_data_1_), .CI(npu_inst_pe_1_0_0_add_79_carry_1_), 
        .CO(npu_inst_pe_1_0_0_add_79_carry_2_), .S(npu_inst_pe_1_0_0_N74) );
  NAND3_X1 npu_inst_pe_1_0_0_U101 ( .A1(npu_inst_pe_1_0_0_n3), .A2(
        npu_inst_pe_1_0_0_n4), .A3(npu_inst_pe_1_0_0_n5), .ZN(
        npu_inst_pe_1_0_0_n44) );
  NAND3_X1 npu_inst_pe_1_0_0_U100 ( .A1(npu_inst_pe_1_0_0_n2), .A2(
        npu_inst_pe_1_0_0_n4), .A3(npu_inst_pe_1_0_0_n5), .ZN(
        npu_inst_pe_1_0_0_n40) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_0_n31), .CK(
        npu_inst_pe_1_0_0_net4478), .RN(npu_inst_pe_1_0_0_n6), .Q(
        int_o_data_npu[62]) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_0_n32), .CK(
        npu_inst_pe_1_0_0_net4478), .RN(npu_inst_pe_1_0_0_n6), .Q(
        int_o_data_npu[61]) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_0_n33), .CK(
        npu_inst_pe_1_0_0_net4478), .RN(npu_inst_pe_1_0_0_n6), .Q(
        int_o_data_npu[60]) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_0_n34), .CK(
        npu_inst_pe_1_0_0_net4478), .RN(npu_inst_pe_1_0_0_n6), .Q(
        int_o_data_npu[59]) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_0_n35), .CK(
        npu_inst_pe_1_0_0_net4478), .RN(npu_inst_pe_1_0_0_n6), .Q(
        int_o_data_npu[58]) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_0_n36), .CK(
        npu_inst_pe_1_0_0_net4478), .RN(npu_inst_pe_1_0_0_n6), .Q(
        int_o_data_npu[57]) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_0_n30), .CK(
        npu_inst_pe_1_0_0_net4478), .RN(npu_inst_pe_1_0_0_n6), .Q(
        int_o_data_npu[63]) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_0_n98), .CK(
        npu_inst_pe_1_0_0_net4478), .RN(npu_inst_pe_1_0_0_n6), .Q(
        int_o_data_npu[56]) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_weight_reg_0_ ( .D(npu_inst_n95), .CK(
        npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n6), .Q(
        npu_inst_pe_1_0_0_int_q_weight_0_), .QN(npu_inst_pe_1_0_0_n27) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_weight_reg_1_ ( .D(npu_inst_n101), .CK(
        npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n6), .Q(
        npu_inst_pe_1_0_0_int_q_weight_1_), .QN(npu_inst_pe_1_0_0_n26) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_0_n110), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n6), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_0_n104), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n6), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_0_n109), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n7), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_0_n103), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n7), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_0_n108), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n7), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_0_n102), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n7), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_0_n107), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n7), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_0_n101), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n7), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_0_n106), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n7), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_0_n100), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n7), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_0_n105), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n7), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_0_n99), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n7), .Q(
        npu_inst_pe_1_0_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_0_n86), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n7), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_0_n87), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n7), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_0_n88), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_0_n89), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_0_n90), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_0_n91), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_0_n92), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_0_n93), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_0_n94), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_0_n95), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_0_n96), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_0_n97), 
        .CK(npu_inst_pe_1_0_0_net4484), .RN(npu_inst_pe_1_0_0_n8), .Q(
        npu_inst_pe_1_0_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_0_net4478) );
  CLKGATETST_X1 npu_inst_pe_1_0_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n48), .SE(1'b0), .GCK(npu_inst_pe_1_0_0_net4484) );
  MUX2_X1 npu_inst_pe_1_0_1_U151 ( .A(npu_inst_pe_1_0_1_n29), .B(
        npu_inst_pe_1_0_1_n24), .S(npu_inst_pe_1_0_1_n5), .Z(
        npu_inst_pe_1_0_1_N93) );
  MUX2_X1 npu_inst_pe_1_0_1_U150 ( .A(npu_inst_pe_1_0_1_n28), .B(
        npu_inst_pe_1_0_1_n25), .S(npu_inst_n62), .Z(npu_inst_pe_1_0_1_n29) );
  MUX2_X1 npu_inst_pe_1_0_1_U149 ( .A(npu_inst_pe_1_0_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_v_1__0_), .S(npu_inst_n54), .Z(
        npu_inst_pe_1_0_1_n28) );
  MUX2_X1 npu_inst_pe_1_0_1_U148 ( .A(npu_inst_pe_1_0_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_v_3__0_), .S(npu_inst_n54), .Z(
        npu_inst_pe_1_0_1_n25) );
  MUX2_X1 npu_inst_pe_1_0_1_U147 ( .A(npu_inst_pe_1_0_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_v_5__0_), .S(npu_inst_n54), .Z(
        npu_inst_pe_1_0_1_n24) );
  MUX2_X1 npu_inst_pe_1_0_1_U146 ( .A(npu_inst_pe_1_0_1_n23), .B(
        npu_inst_pe_1_0_1_n20), .S(npu_inst_pe_1_0_1_n5), .Z(
        npu_inst_pe_1_0_1_N94) );
  MUX2_X1 npu_inst_pe_1_0_1_U145 ( .A(npu_inst_pe_1_0_1_n22), .B(
        npu_inst_pe_1_0_1_n21), .S(npu_inst_n62), .Z(npu_inst_pe_1_0_1_n23) );
  MUX2_X1 npu_inst_pe_1_0_1_U144 ( .A(npu_inst_pe_1_0_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_v_1__1_), .S(npu_inst_n54), .Z(
        npu_inst_pe_1_0_1_n22) );
  MUX2_X1 npu_inst_pe_1_0_1_U143 ( .A(npu_inst_pe_1_0_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_v_3__1_), .S(npu_inst_n54), .Z(
        npu_inst_pe_1_0_1_n21) );
  MUX2_X1 npu_inst_pe_1_0_1_U142 ( .A(npu_inst_pe_1_0_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_v_5__1_), .S(npu_inst_n54), .Z(
        npu_inst_pe_1_0_1_n20) );
  MUX2_X1 npu_inst_pe_1_0_1_U141 ( .A(npu_inst_pe_1_0_1_n19), .B(
        npu_inst_pe_1_0_1_n16), .S(npu_inst_pe_1_0_1_n5), .Z(
        npu_inst_int_data_x_0__1__1_) );
  MUX2_X1 npu_inst_pe_1_0_1_U140 ( .A(npu_inst_pe_1_0_1_n18), .B(
        npu_inst_pe_1_0_1_n17), .S(npu_inst_n62), .Z(npu_inst_pe_1_0_1_n19) );
  MUX2_X1 npu_inst_pe_1_0_1_U139 ( .A(npu_inst_pe_1_0_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_h_1__1_), .S(npu_inst_n54), .Z(
        npu_inst_pe_1_0_1_n18) );
  MUX2_X1 npu_inst_pe_1_0_1_U138 ( .A(npu_inst_pe_1_0_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_h_3__1_), .S(npu_inst_n54), .Z(
        npu_inst_pe_1_0_1_n17) );
  MUX2_X1 npu_inst_pe_1_0_1_U137 ( .A(npu_inst_pe_1_0_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_h_5__1_), .S(npu_inst_n54), .Z(
        npu_inst_pe_1_0_1_n16) );
  MUX2_X1 npu_inst_pe_1_0_1_U136 ( .A(npu_inst_pe_1_0_1_n15), .B(
        npu_inst_pe_1_0_1_n12), .S(npu_inst_pe_1_0_1_n5), .Z(
        npu_inst_int_data_x_0__1__0_) );
  MUX2_X1 npu_inst_pe_1_0_1_U135 ( .A(npu_inst_pe_1_0_1_n14), .B(
        npu_inst_pe_1_0_1_n13), .S(npu_inst_n62), .Z(npu_inst_pe_1_0_1_n15) );
  MUX2_X1 npu_inst_pe_1_0_1_U134 ( .A(npu_inst_pe_1_0_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_h_1__0_), .S(npu_inst_n54), .Z(
        npu_inst_pe_1_0_1_n14) );
  MUX2_X1 npu_inst_pe_1_0_1_U133 ( .A(npu_inst_pe_1_0_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_h_3__0_), .S(npu_inst_n54), .Z(
        npu_inst_pe_1_0_1_n13) );
  MUX2_X1 npu_inst_pe_1_0_1_U132 ( .A(npu_inst_pe_1_0_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_1_int_q_reg_h_5__0_), .S(npu_inst_n54), .Z(
        npu_inst_pe_1_0_1_n12) );
  XOR2_X1 npu_inst_pe_1_0_1_U131 ( .A(npu_inst_pe_1_0_1_int_data_0_), .B(
        int_o_data_npu[48]), .Z(npu_inst_pe_1_0_1_N73) );
  AND2_X1 npu_inst_pe_1_0_1_U130 ( .A1(int_o_data_npu[48]), .A2(
        npu_inst_pe_1_0_1_int_data_0_), .ZN(npu_inst_pe_1_0_1_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_1_U129 ( .A(int_o_data_npu[48]), .B(
        npu_inst_pe_1_0_1_n10), .ZN(npu_inst_pe_1_0_1_N65) );
  OR2_X1 npu_inst_pe_1_0_1_U128 ( .A1(npu_inst_pe_1_0_1_n10), .A2(
        int_o_data_npu[48]), .ZN(npu_inst_pe_1_0_1_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_1_U127 ( .A(int_o_data_npu[50]), .B(
        npu_inst_pe_1_0_1_add_79_carry_2_), .Z(npu_inst_pe_1_0_1_N75) );
  AND2_X1 npu_inst_pe_1_0_1_U126 ( .A1(npu_inst_pe_1_0_1_add_79_carry_2_), 
        .A2(int_o_data_npu[50]), .ZN(npu_inst_pe_1_0_1_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_1_U125 ( .A(int_o_data_npu[51]), .B(
        npu_inst_pe_1_0_1_add_79_carry_3_), .Z(npu_inst_pe_1_0_1_N76) );
  AND2_X1 npu_inst_pe_1_0_1_U124 ( .A1(npu_inst_pe_1_0_1_add_79_carry_3_), 
        .A2(int_o_data_npu[51]), .ZN(npu_inst_pe_1_0_1_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_1_U123 ( .A(int_o_data_npu[52]), .B(
        npu_inst_pe_1_0_1_add_79_carry_4_), .Z(npu_inst_pe_1_0_1_N77) );
  AND2_X1 npu_inst_pe_1_0_1_U122 ( .A1(npu_inst_pe_1_0_1_add_79_carry_4_), 
        .A2(int_o_data_npu[52]), .ZN(npu_inst_pe_1_0_1_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_1_U121 ( .A(int_o_data_npu[53]), .B(
        npu_inst_pe_1_0_1_add_79_carry_5_), .Z(npu_inst_pe_1_0_1_N78) );
  AND2_X1 npu_inst_pe_1_0_1_U120 ( .A1(npu_inst_pe_1_0_1_add_79_carry_5_), 
        .A2(int_o_data_npu[53]), .ZN(npu_inst_pe_1_0_1_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_1_U119 ( .A(int_o_data_npu[54]), .B(
        npu_inst_pe_1_0_1_add_79_carry_6_), .Z(npu_inst_pe_1_0_1_N79) );
  AND2_X1 npu_inst_pe_1_0_1_U118 ( .A1(npu_inst_pe_1_0_1_add_79_carry_6_), 
        .A2(int_o_data_npu[54]), .ZN(npu_inst_pe_1_0_1_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_1_U117 ( .A(int_o_data_npu[55]), .B(
        npu_inst_pe_1_0_1_add_79_carry_7_), .Z(npu_inst_pe_1_0_1_N80) );
  XNOR2_X1 npu_inst_pe_1_0_1_U116 ( .A(npu_inst_pe_1_0_1_sub_77_carry_2_), .B(
        int_o_data_npu[50]), .ZN(npu_inst_pe_1_0_1_N67) );
  OR2_X1 npu_inst_pe_1_0_1_U115 ( .A1(int_o_data_npu[50]), .A2(
        npu_inst_pe_1_0_1_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_0_1_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_1_U114 ( .A(npu_inst_pe_1_0_1_sub_77_carry_3_), .B(
        int_o_data_npu[51]), .ZN(npu_inst_pe_1_0_1_N68) );
  OR2_X1 npu_inst_pe_1_0_1_U113 ( .A1(int_o_data_npu[51]), .A2(
        npu_inst_pe_1_0_1_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_0_1_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_1_U112 ( .A(npu_inst_pe_1_0_1_sub_77_carry_4_), .B(
        int_o_data_npu[52]), .ZN(npu_inst_pe_1_0_1_N69) );
  OR2_X1 npu_inst_pe_1_0_1_U111 ( .A1(int_o_data_npu[52]), .A2(
        npu_inst_pe_1_0_1_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_0_1_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_1_U110 ( .A(npu_inst_pe_1_0_1_sub_77_carry_5_), .B(
        int_o_data_npu[53]), .ZN(npu_inst_pe_1_0_1_N70) );
  OR2_X1 npu_inst_pe_1_0_1_U109 ( .A1(int_o_data_npu[53]), .A2(
        npu_inst_pe_1_0_1_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_0_1_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_1_U108 ( .A(npu_inst_pe_1_0_1_sub_77_carry_6_), .B(
        int_o_data_npu[54]), .ZN(npu_inst_pe_1_0_1_N71) );
  OR2_X1 npu_inst_pe_1_0_1_U107 ( .A1(int_o_data_npu[54]), .A2(
        npu_inst_pe_1_0_1_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_0_1_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_1_U106 ( .A(int_o_data_npu[55]), .B(
        npu_inst_pe_1_0_1_sub_77_carry_7_), .ZN(npu_inst_pe_1_0_1_N72) );
  INV_X1 npu_inst_pe_1_0_1_U105 ( .A(npu_inst_n62), .ZN(npu_inst_pe_1_0_1_n4)
         );
  INV_X1 npu_inst_pe_1_0_1_U104 ( .A(npu_inst_n42), .ZN(npu_inst_pe_1_0_1_n2)
         );
  AOI22_X1 npu_inst_pe_1_0_1_U103 ( .A1(npu_inst_int_data_y_1__1__0_), .A2(
        npu_inst_pe_1_0_1_n58), .B1(npu_inst_pe_1_0_1_n116), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_1_n57) );
  INV_X1 npu_inst_pe_1_0_1_U102 ( .A(npu_inst_pe_1_0_1_n57), .ZN(
        npu_inst_pe_1_0_1_n105) );
  AOI22_X1 npu_inst_pe_1_0_1_U99 ( .A1(npu_inst_int_data_y_1__1__0_), .A2(
        npu_inst_pe_1_0_1_n54), .B1(npu_inst_pe_1_0_1_n115), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_1_n53) );
  INV_X1 npu_inst_pe_1_0_1_U98 ( .A(npu_inst_pe_1_0_1_n53), .ZN(
        npu_inst_pe_1_0_1_n106) );
  AOI22_X1 npu_inst_pe_1_0_1_U97 ( .A1(npu_inst_int_data_y_1__1__0_), .A2(
        npu_inst_pe_1_0_1_n50), .B1(npu_inst_pe_1_0_1_n114), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_1_n49) );
  INV_X1 npu_inst_pe_1_0_1_U96 ( .A(npu_inst_pe_1_0_1_n49), .ZN(
        npu_inst_pe_1_0_1_n107) );
  AOI22_X1 npu_inst_pe_1_0_1_U95 ( .A1(npu_inst_int_data_y_1__1__0_), .A2(
        npu_inst_pe_1_0_1_n46), .B1(npu_inst_pe_1_0_1_n113), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_1_n45) );
  INV_X1 npu_inst_pe_1_0_1_U94 ( .A(npu_inst_pe_1_0_1_n45), .ZN(
        npu_inst_pe_1_0_1_n108) );
  AOI22_X1 npu_inst_pe_1_0_1_U93 ( .A1(npu_inst_int_data_y_1__1__0_), .A2(
        npu_inst_pe_1_0_1_n42), .B1(npu_inst_pe_1_0_1_n112), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_1_n41) );
  INV_X1 npu_inst_pe_1_0_1_U92 ( .A(npu_inst_pe_1_0_1_n41), .ZN(
        npu_inst_pe_1_0_1_n109) );
  AOI22_X1 npu_inst_pe_1_0_1_U91 ( .A1(npu_inst_int_data_y_1__1__1_), .A2(
        npu_inst_pe_1_0_1_n58), .B1(npu_inst_pe_1_0_1_n116), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_1_n59) );
  INV_X1 npu_inst_pe_1_0_1_U90 ( .A(npu_inst_pe_1_0_1_n59), .ZN(
        npu_inst_pe_1_0_1_n99) );
  AOI22_X1 npu_inst_pe_1_0_1_U89 ( .A1(npu_inst_int_data_y_1__1__1_), .A2(
        npu_inst_pe_1_0_1_n54), .B1(npu_inst_pe_1_0_1_n115), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_1_n55) );
  INV_X1 npu_inst_pe_1_0_1_U88 ( .A(npu_inst_pe_1_0_1_n55), .ZN(
        npu_inst_pe_1_0_1_n100) );
  AOI22_X1 npu_inst_pe_1_0_1_U87 ( .A1(npu_inst_int_data_y_1__1__1_), .A2(
        npu_inst_pe_1_0_1_n50), .B1(npu_inst_pe_1_0_1_n114), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_1_n51) );
  INV_X1 npu_inst_pe_1_0_1_U86 ( .A(npu_inst_pe_1_0_1_n51), .ZN(
        npu_inst_pe_1_0_1_n101) );
  AOI22_X1 npu_inst_pe_1_0_1_U85 ( .A1(npu_inst_int_data_y_1__1__1_), .A2(
        npu_inst_pe_1_0_1_n46), .B1(npu_inst_pe_1_0_1_n113), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_1_n47) );
  INV_X1 npu_inst_pe_1_0_1_U84 ( .A(npu_inst_pe_1_0_1_n47), .ZN(
        npu_inst_pe_1_0_1_n102) );
  AOI22_X1 npu_inst_pe_1_0_1_U83 ( .A1(npu_inst_int_data_y_1__1__1_), .A2(
        npu_inst_pe_1_0_1_n42), .B1(npu_inst_pe_1_0_1_n112), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_1_n43) );
  INV_X1 npu_inst_pe_1_0_1_U82 ( .A(npu_inst_pe_1_0_1_n43), .ZN(
        npu_inst_pe_1_0_1_n103) );
  AOI22_X1 npu_inst_pe_1_0_1_U81 ( .A1(npu_inst_pe_1_0_1_n38), .A2(
        npu_inst_int_data_y_1__1__1_), .B1(npu_inst_pe_1_0_1_n111), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_1_n39) );
  INV_X1 npu_inst_pe_1_0_1_U80 ( .A(npu_inst_pe_1_0_1_n39), .ZN(
        npu_inst_pe_1_0_1_n104) );
  NAND2_X1 npu_inst_pe_1_0_1_U79 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_1_n60), .ZN(npu_inst_pe_1_0_1_n74) );
  OAI21_X1 npu_inst_pe_1_0_1_U78 ( .B1(npu_inst_pe_1_0_1_n63), .B2(
        npu_inst_pe_1_0_1_n60), .A(npu_inst_pe_1_0_1_n74), .ZN(
        npu_inst_pe_1_0_1_n97) );
  NAND2_X1 npu_inst_pe_1_0_1_U77 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_1_n60), .ZN(npu_inst_pe_1_0_1_n73) );
  OAI21_X1 npu_inst_pe_1_0_1_U76 ( .B1(npu_inst_pe_1_0_1_n61), .B2(
        npu_inst_pe_1_0_1_n60), .A(npu_inst_pe_1_0_1_n73), .ZN(
        npu_inst_pe_1_0_1_n96) );
  NAND2_X1 npu_inst_pe_1_0_1_U75 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_1_n56), .ZN(npu_inst_pe_1_0_1_n72) );
  OAI21_X1 npu_inst_pe_1_0_1_U74 ( .B1(npu_inst_pe_1_0_1_n63), .B2(
        npu_inst_pe_1_0_1_n56), .A(npu_inst_pe_1_0_1_n72), .ZN(
        npu_inst_pe_1_0_1_n95) );
  NAND2_X1 npu_inst_pe_1_0_1_U73 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_1_n56), .ZN(npu_inst_pe_1_0_1_n71) );
  OAI21_X1 npu_inst_pe_1_0_1_U72 ( .B1(npu_inst_pe_1_0_1_n61), .B2(
        npu_inst_pe_1_0_1_n56), .A(npu_inst_pe_1_0_1_n71), .ZN(
        npu_inst_pe_1_0_1_n94) );
  NAND2_X1 npu_inst_pe_1_0_1_U71 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_1_n52), .ZN(npu_inst_pe_1_0_1_n70) );
  OAI21_X1 npu_inst_pe_1_0_1_U70 ( .B1(npu_inst_pe_1_0_1_n63), .B2(
        npu_inst_pe_1_0_1_n52), .A(npu_inst_pe_1_0_1_n70), .ZN(
        npu_inst_pe_1_0_1_n93) );
  NAND2_X1 npu_inst_pe_1_0_1_U69 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_1_n52), .ZN(npu_inst_pe_1_0_1_n69) );
  OAI21_X1 npu_inst_pe_1_0_1_U68 ( .B1(npu_inst_pe_1_0_1_n61), .B2(
        npu_inst_pe_1_0_1_n52), .A(npu_inst_pe_1_0_1_n69), .ZN(
        npu_inst_pe_1_0_1_n92) );
  NAND2_X1 npu_inst_pe_1_0_1_U67 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_1_n48), .ZN(npu_inst_pe_1_0_1_n68) );
  OAI21_X1 npu_inst_pe_1_0_1_U66 ( .B1(npu_inst_pe_1_0_1_n63), .B2(
        npu_inst_pe_1_0_1_n48), .A(npu_inst_pe_1_0_1_n68), .ZN(
        npu_inst_pe_1_0_1_n91) );
  NAND2_X1 npu_inst_pe_1_0_1_U65 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_1_n48), .ZN(npu_inst_pe_1_0_1_n67) );
  OAI21_X1 npu_inst_pe_1_0_1_U64 ( .B1(npu_inst_pe_1_0_1_n61), .B2(
        npu_inst_pe_1_0_1_n48), .A(npu_inst_pe_1_0_1_n67), .ZN(
        npu_inst_pe_1_0_1_n90) );
  NAND2_X1 npu_inst_pe_1_0_1_U63 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_1_n44), .ZN(npu_inst_pe_1_0_1_n66) );
  OAI21_X1 npu_inst_pe_1_0_1_U62 ( .B1(npu_inst_pe_1_0_1_n63), .B2(
        npu_inst_pe_1_0_1_n44), .A(npu_inst_pe_1_0_1_n66), .ZN(
        npu_inst_pe_1_0_1_n89) );
  NAND2_X1 npu_inst_pe_1_0_1_U61 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_1_n44), .ZN(npu_inst_pe_1_0_1_n65) );
  OAI21_X1 npu_inst_pe_1_0_1_U60 ( .B1(npu_inst_pe_1_0_1_n61), .B2(
        npu_inst_pe_1_0_1_n44), .A(npu_inst_pe_1_0_1_n65), .ZN(
        npu_inst_pe_1_0_1_n88) );
  NAND2_X1 npu_inst_pe_1_0_1_U59 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_1_n40), .ZN(npu_inst_pe_1_0_1_n64) );
  OAI21_X1 npu_inst_pe_1_0_1_U58 ( .B1(npu_inst_pe_1_0_1_n63), .B2(
        npu_inst_pe_1_0_1_n40), .A(npu_inst_pe_1_0_1_n64), .ZN(
        npu_inst_pe_1_0_1_n87) );
  NAND2_X1 npu_inst_pe_1_0_1_U57 ( .A1(npu_inst_pe_1_0_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_1_n40), .ZN(npu_inst_pe_1_0_1_n62) );
  OAI21_X1 npu_inst_pe_1_0_1_U56 ( .B1(npu_inst_pe_1_0_1_n61), .B2(
        npu_inst_pe_1_0_1_n40), .A(npu_inst_pe_1_0_1_n62), .ZN(
        npu_inst_pe_1_0_1_n86) );
  AOI22_X1 npu_inst_pe_1_0_1_U55 ( .A1(npu_inst_pe_1_0_1_n38), .A2(
        npu_inst_int_data_y_1__1__0_), .B1(npu_inst_pe_1_0_1_n111), .B2(
        npu_inst_pe_1_0_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_1_n37) );
  INV_X1 npu_inst_pe_1_0_1_U54 ( .A(npu_inst_pe_1_0_1_n37), .ZN(
        npu_inst_pe_1_0_1_n110) );
  AOI222_X1 npu_inst_pe_1_0_1_U53 ( .A1(npu_inst_int_data_res_1__1__0_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N73), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N65), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n84) );
  INV_X1 npu_inst_pe_1_0_1_U52 ( .A(npu_inst_pe_1_0_1_n84), .ZN(
        npu_inst_pe_1_0_1_n98) );
  AOI222_X1 npu_inst_pe_1_0_1_U51 ( .A1(npu_inst_pe_1_0_1_n1), .A2(
        npu_inst_int_data_res_1__1__7_), .B1(npu_inst_pe_1_0_1_N80), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N72), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n75) );
  INV_X1 npu_inst_pe_1_0_1_U50 ( .A(npu_inst_pe_1_0_1_n75), .ZN(
        npu_inst_pe_1_0_1_n30) );
  AOI222_X1 npu_inst_pe_1_0_1_U49 ( .A1(npu_inst_int_data_res_1__1__2_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N75), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N67), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n82) );
  INV_X1 npu_inst_pe_1_0_1_U48 ( .A(npu_inst_pe_1_0_1_n82), .ZN(
        npu_inst_pe_1_0_1_n35) );
  AOI222_X1 npu_inst_pe_1_0_1_U47 ( .A1(npu_inst_int_data_res_1__1__3_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N76), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N68), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n81) );
  INV_X1 npu_inst_pe_1_0_1_U46 ( .A(npu_inst_pe_1_0_1_n81), .ZN(
        npu_inst_pe_1_0_1_n34) );
  AOI222_X1 npu_inst_pe_1_0_1_U45 ( .A1(npu_inst_int_data_res_1__1__4_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N77), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N69), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n80) );
  INV_X1 npu_inst_pe_1_0_1_U44 ( .A(npu_inst_pe_1_0_1_n80), .ZN(
        npu_inst_pe_1_0_1_n33) );
  AOI222_X1 npu_inst_pe_1_0_1_U43 ( .A1(npu_inst_int_data_res_1__1__5_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N78), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N70), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n79) );
  INV_X1 npu_inst_pe_1_0_1_U42 ( .A(npu_inst_pe_1_0_1_n79), .ZN(
        npu_inst_pe_1_0_1_n32) );
  AOI222_X1 npu_inst_pe_1_0_1_U41 ( .A1(npu_inst_int_data_res_1__1__6_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N79), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N71), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n78) );
  INV_X1 npu_inst_pe_1_0_1_U40 ( .A(npu_inst_pe_1_0_1_n78), .ZN(
        npu_inst_pe_1_0_1_n31) );
  NOR3_X1 npu_inst_pe_1_0_1_U39 ( .A1(npu_inst_pe_1_0_1_n26), .A2(npu_inst_n42), .A3(npu_inst_int_ckg[62]), .ZN(npu_inst_pe_1_0_1_n85) );
  OR2_X1 npu_inst_pe_1_0_1_U38 ( .A1(npu_inst_pe_1_0_1_n85), .A2(
        npu_inst_pe_1_0_1_n1), .ZN(npu_inst_pe_1_0_1_N84) );
  AND2_X1 npu_inst_pe_1_0_1_U37 ( .A1(npu_inst_int_data_x_0__1__1_), .A2(
        npu_inst_pe_1_0_1_int_q_weight_1_), .ZN(npu_inst_pe_1_0_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_1_U36 ( .A1(npu_inst_int_data_x_0__1__0_), .A2(
        npu_inst_pe_1_0_1_int_q_weight_1_), .ZN(npu_inst_pe_1_0_1_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_0_1_U35 ( .A(npu_inst_pe_1_0_1_int_data_1_), .ZN(
        npu_inst_pe_1_0_1_n11) );
  AOI222_X1 npu_inst_pe_1_0_1_U34 ( .A1(npu_inst_int_data_res_1__1__1_), .A2(
        npu_inst_pe_1_0_1_n1), .B1(npu_inst_pe_1_0_1_N74), .B2(
        npu_inst_pe_1_0_1_n76), .C1(npu_inst_pe_1_0_1_N66), .C2(
        npu_inst_pe_1_0_1_n77), .ZN(npu_inst_pe_1_0_1_n83) );
  INV_X1 npu_inst_pe_1_0_1_U33 ( .A(npu_inst_pe_1_0_1_n83), .ZN(
        npu_inst_pe_1_0_1_n36) );
  AND2_X1 npu_inst_pe_1_0_1_U32 ( .A1(npu_inst_pe_1_0_1_N93), .A2(npu_inst_n42), .ZN(npu_inst_pe_1_0_1_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_1_U31 ( .A1(npu_inst_n42), .A2(npu_inst_pe_1_0_1_N94), .ZN(npu_inst_pe_1_0_1_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_1_U30 ( .A1(npu_inst_n42), .A2(
        npu_inst_int_data_y_1__1__1_), .B1(npu_inst_pe_1_0_1_n2), .B2(
        npu_inst_int_data_x_0__2__1_), .ZN(npu_inst_pe_1_0_1_n63) );
  AOI22_X1 npu_inst_pe_1_0_1_U29 ( .A1(npu_inst_n42), .A2(
        npu_inst_int_data_y_1__1__0_), .B1(npu_inst_pe_1_0_1_n2), .B2(
        npu_inst_int_data_x_0__2__0_), .ZN(npu_inst_pe_1_0_1_n61) );
  INV_X1 npu_inst_pe_1_0_1_U28 ( .A(npu_inst_pe_1_0_1_int_data_0_), .ZN(
        npu_inst_pe_1_0_1_n10) );
  INV_X1 npu_inst_pe_1_0_1_U27 ( .A(npu_inst_n54), .ZN(npu_inst_pe_1_0_1_n3)
         );
  OR3_X1 npu_inst_pe_1_0_1_U26 ( .A1(npu_inst_n62), .A2(npu_inst_pe_1_0_1_n5), 
        .A3(npu_inst_pe_1_0_1_n3), .ZN(npu_inst_pe_1_0_1_n56) );
  OR3_X1 npu_inst_pe_1_0_1_U25 ( .A1(npu_inst_pe_1_0_1_n3), .A2(
        npu_inst_pe_1_0_1_n5), .A3(npu_inst_pe_1_0_1_n4), .ZN(
        npu_inst_pe_1_0_1_n48) );
  OR3_X1 npu_inst_pe_1_0_1_U24 ( .A1(npu_inst_n54), .A2(npu_inst_pe_1_0_1_n5), 
        .A3(npu_inst_pe_1_0_1_n4), .ZN(npu_inst_pe_1_0_1_n52) );
  OR3_X1 npu_inst_pe_1_0_1_U23 ( .A1(npu_inst_n62), .A2(npu_inst_pe_1_0_1_n5), 
        .A3(npu_inst_n54), .ZN(npu_inst_pe_1_0_1_n60) );
  BUF_X1 npu_inst_pe_1_0_1_U22 ( .A(npu_inst_n31), .Z(npu_inst_pe_1_0_1_n1) );
  NOR2_X1 npu_inst_pe_1_0_1_U21 ( .A1(npu_inst_pe_1_0_1_n60), .A2(
        npu_inst_pe_1_0_1_n2), .ZN(npu_inst_pe_1_0_1_n58) );
  NOR2_X1 npu_inst_pe_1_0_1_U20 ( .A1(npu_inst_pe_1_0_1_n56), .A2(
        npu_inst_pe_1_0_1_n2), .ZN(npu_inst_pe_1_0_1_n54) );
  NOR2_X1 npu_inst_pe_1_0_1_U19 ( .A1(npu_inst_pe_1_0_1_n52), .A2(
        npu_inst_pe_1_0_1_n2), .ZN(npu_inst_pe_1_0_1_n50) );
  NOR2_X1 npu_inst_pe_1_0_1_U18 ( .A1(npu_inst_pe_1_0_1_n48), .A2(
        npu_inst_pe_1_0_1_n2), .ZN(npu_inst_pe_1_0_1_n46) );
  NOR2_X1 npu_inst_pe_1_0_1_U17 ( .A1(npu_inst_pe_1_0_1_n40), .A2(
        npu_inst_pe_1_0_1_n2), .ZN(npu_inst_pe_1_0_1_n38) );
  NOR2_X1 npu_inst_pe_1_0_1_U16 ( .A1(npu_inst_pe_1_0_1_n44), .A2(
        npu_inst_pe_1_0_1_n2), .ZN(npu_inst_pe_1_0_1_n42) );
  BUF_X1 npu_inst_pe_1_0_1_U15 ( .A(npu_inst_n89), .Z(npu_inst_pe_1_0_1_n5) );
  INV_X1 npu_inst_pe_1_0_1_U14 ( .A(npu_inst_n109), .ZN(npu_inst_pe_1_0_1_n9)
         );
  INV_X1 npu_inst_pe_1_0_1_U13 ( .A(npu_inst_pe_1_0_1_n38), .ZN(
        npu_inst_pe_1_0_1_n111) );
  INV_X1 npu_inst_pe_1_0_1_U12 ( .A(npu_inst_pe_1_0_1_n58), .ZN(
        npu_inst_pe_1_0_1_n116) );
  INV_X1 npu_inst_pe_1_0_1_U11 ( .A(npu_inst_pe_1_0_1_n54), .ZN(
        npu_inst_pe_1_0_1_n115) );
  INV_X1 npu_inst_pe_1_0_1_U10 ( .A(npu_inst_pe_1_0_1_n50), .ZN(
        npu_inst_pe_1_0_1_n114) );
  INV_X1 npu_inst_pe_1_0_1_U9 ( .A(npu_inst_pe_1_0_1_n46), .ZN(
        npu_inst_pe_1_0_1_n113) );
  INV_X1 npu_inst_pe_1_0_1_U8 ( .A(npu_inst_pe_1_0_1_n42), .ZN(
        npu_inst_pe_1_0_1_n112) );
  BUF_X1 npu_inst_pe_1_0_1_U7 ( .A(npu_inst_pe_1_0_1_n9), .Z(
        npu_inst_pe_1_0_1_n8) );
  BUF_X1 npu_inst_pe_1_0_1_U6 ( .A(npu_inst_pe_1_0_1_n9), .Z(
        npu_inst_pe_1_0_1_n7) );
  BUF_X1 npu_inst_pe_1_0_1_U5 ( .A(npu_inst_pe_1_0_1_n9), .Z(
        npu_inst_pe_1_0_1_n6) );
  NOR2_X1 npu_inst_pe_1_0_1_U4 ( .A1(npu_inst_pe_1_0_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_1_n1), .ZN(npu_inst_pe_1_0_1_n76) );
  NOR2_X1 npu_inst_pe_1_0_1_U3 ( .A1(npu_inst_pe_1_0_1_n27), .A2(
        npu_inst_pe_1_0_1_n1), .ZN(npu_inst_pe_1_0_1_n77) );
  FA_X1 npu_inst_pe_1_0_1_sub_77_U2_1 ( .A(int_o_data_npu[49]), .B(
        npu_inst_pe_1_0_1_n11), .CI(npu_inst_pe_1_0_1_sub_77_carry_1_), .CO(
        npu_inst_pe_1_0_1_sub_77_carry_2_), .S(npu_inst_pe_1_0_1_N66) );
  FA_X1 npu_inst_pe_1_0_1_add_79_U1_1 ( .A(int_o_data_npu[49]), .B(
        npu_inst_pe_1_0_1_int_data_1_), .CI(npu_inst_pe_1_0_1_add_79_carry_1_), 
        .CO(npu_inst_pe_1_0_1_add_79_carry_2_), .S(npu_inst_pe_1_0_1_N74) );
  NAND3_X1 npu_inst_pe_1_0_1_U101 ( .A1(npu_inst_pe_1_0_1_n3), .A2(
        npu_inst_pe_1_0_1_n4), .A3(npu_inst_pe_1_0_1_n5), .ZN(
        npu_inst_pe_1_0_1_n44) );
  NAND3_X1 npu_inst_pe_1_0_1_U100 ( .A1(npu_inst_n54), .A2(
        npu_inst_pe_1_0_1_n4), .A3(npu_inst_pe_1_0_1_n5), .ZN(
        npu_inst_pe_1_0_1_n40) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_1_n31), .CK(
        npu_inst_pe_1_0_1_net4455), .RN(npu_inst_pe_1_0_1_n6), .Q(
        int_o_data_npu[54]) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_1_n32), .CK(
        npu_inst_pe_1_0_1_net4455), .RN(npu_inst_pe_1_0_1_n6), .Q(
        int_o_data_npu[53]) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_1_n33), .CK(
        npu_inst_pe_1_0_1_net4455), .RN(npu_inst_pe_1_0_1_n6), .Q(
        int_o_data_npu[52]) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_1_n34), .CK(
        npu_inst_pe_1_0_1_net4455), .RN(npu_inst_pe_1_0_1_n6), .Q(
        int_o_data_npu[51]) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_1_n35), .CK(
        npu_inst_pe_1_0_1_net4455), .RN(npu_inst_pe_1_0_1_n6), .Q(
        int_o_data_npu[50]) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_1_n36), .CK(
        npu_inst_pe_1_0_1_net4455), .RN(npu_inst_pe_1_0_1_n6), .Q(
        int_o_data_npu[49]) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_1_n30), .CK(
        npu_inst_pe_1_0_1_net4455), .RN(npu_inst_pe_1_0_1_n6), .Q(
        int_o_data_npu[55]) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_1_n98), .CK(
        npu_inst_pe_1_0_1_net4455), .RN(npu_inst_pe_1_0_1_n6), .Q(
        int_o_data_npu[48]) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_weight_reg_0_ ( .D(npu_inst_n95), .CK(
        npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n6), .Q(
        npu_inst_pe_1_0_1_int_q_weight_0_), .QN(npu_inst_pe_1_0_1_n27) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_weight_reg_1_ ( .D(npu_inst_n101), .CK(
        npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n6), .Q(
        npu_inst_pe_1_0_1_int_q_weight_1_), .QN(npu_inst_pe_1_0_1_n26) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_1_n110), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n6), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_1_n104), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n6), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_1_n109), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_1_n103), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_1_n108), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_1_n102), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_1_n107), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_1_n101), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_1_n106), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_1_n100), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_1_n105), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_1_n99), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_1_n86), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_1_n87), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n7), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_1_n88), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_1_n89), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_1_n90), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_1_n91), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_1_n92), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_1_n93), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_1_n94), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_1_n95), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_1_n96), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_1_n97), 
        .CK(npu_inst_pe_1_0_1_net4461), .RN(npu_inst_pe_1_0_1_n8), .Q(
        npu_inst_pe_1_0_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_1_net4455) );
  CLKGATETST_X1 npu_inst_pe_1_0_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n48), .SE(1'b0), .GCK(npu_inst_pe_1_0_1_net4461) );
  MUX2_X1 npu_inst_pe_1_0_2_U152 ( .A(npu_inst_pe_1_0_2_n30), .B(
        npu_inst_pe_1_0_2_n25), .S(npu_inst_pe_1_0_2_n6), .Z(
        npu_inst_pe_1_0_2_N93) );
  MUX2_X1 npu_inst_pe_1_0_2_U151 ( .A(npu_inst_pe_1_0_2_n29), .B(
        npu_inst_pe_1_0_2_n28), .S(npu_inst_n62), .Z(npu_inst_pe_1_0_2_n30) );
  MUX2_X1 npu_inst_pe_1_0_2_U150 ( .A(npu_inst_pe_1_0_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_2_n3), .Z(
        npu_inst_pe_1_0_2_n29) );
  MUX2_X1 npu_inst_pe_1_0_2_U149 ( .A(npu_inst_pe_1_0_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_2_n3), .Z(
        npu_inst_pe_1_0_2_n28) );
  MUX2_X1 npu_inst_pe_1_0_2_U148 ( .A(npu_inst_pe_1_0_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_2_n3), .Z(
        npu_inst_pe_1_0_2_n25) );
  MUX2_X1 npu_inst_pe_1_0_2_U147 ( .A(npu_inst_pe_1_0_2_n24), .B(
        npu_inst_pe_1_0_2_n21), .S(npu_inst_pe_1_0_2_n6), .Z(
        npu_inst_pe_1_0_2_N94) );
  MUX2_X1 npu_inst_pe_1_0_2_U146 ( .A(npu_inst_pe_1_0_2_n23), .B(
        npu_inst_pe_1_0_2_n22), .S(npu_inst_n62), .Z(npu_inst_pe_1_0_2_n24) );
  MUX2_X1 npu_inst_pe_1_0_2_U145 ( .A(npu_inst_pe_1_0_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_2_n3), .Z(
        npu_inst_pe_1_0_2_n23) );
  MUX2_X1 npu_inst_pe_1_0_2_U144 ( .A(npu_inst_pe_1_0_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_2_n3), .Z(
        npu_inst_pe_1_0_2_n22) );
  MUX2_X1 npu_inst_pe_1_0_2_U143 ( .A(npu_inst_pe_1_0_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_2_n3), .Z(
        npu_inst_pe_1_0_2_n21) );
  MUX2_X1 npu_inst_pe_1_0_2_U142 ( .A(npu_inst_pe_1_0_2_n20), .B(
        npu_inst_pe_1_0_2_n17), .S(npu_inst_pe_1_0_2_n6), .Z(
        npu_inst_int_data_x_0__2__1_) );
  MUX2_X1 npu_inst_pe_1_0_2_U141 ( .A(npu_inst_pe_1_0_2_n19), .B(
        npu_inst_pe_1_0_2_n18), .S(npu_inst_n62), .Z(npu_inst_pe_1_0_2_n20) );
  MUX2_X1 npu_inst_pe_1_0_2_U140 ( .A(npu_inst_pe_1_0_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_2_n3), .Z(
        npu_inst_pe_1_0_2_n19) );
  MUX2_X1 npu_inst_pe_1_0_2_U139 ( .A(npu_inst_pe_1_0_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_2_n3), .Z(
        npu_inst_pe_1_0_2_n18) );
  MUX2_X1 npu_inst_pe_1_0_2_U138 ( .A(npu_inst_pe_1_0_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_2_n3), .Z(
        npu_inst_pe_1_0_2_n17) );
  MUX2_X1 npu_inst_pe_1_0_2_U137 ( .A(npu_inst_pe_1_0_2_n16), .B(
        npu_inst_pe_1_0_2_n13), .S(npu_inst_pe_1_0_2_n6), .Z(
        npu_inst_int_data_x_0__2__0_) );
  MUX2_X1 npu_inst_pe_1_0_2_U136 ( .A(npu_inst_pe_1_0_2_n15), .B(
        npu_inst_pe_1_0_2_n14), .S(npu_inst_n62), .Z(npu_inst_pe_1_0_2_n16) );
  MUX2_X1 npu_inst_pe_1_0_2_U135 ( .A(npu_inst_pe_1_0_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_2_n3), .Z(
        npu_inst_pe_1_0_2_n15) );
  MUX2_X1 npu_inst_pe_1_0_2_U134 ( .A(npu_inst_pe_1_0_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_2_n3), .Z(
        npu_inst_pe_1_0_2_n14) );
  MUX2_X1 npu_inst_pe_1_0_2_U133 ( .A(npu_inst_pe_1_0_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_2_n3), .Z(
        npu_inst_pe_1_0_2_n13) );
  XOR2_X1 npu_inst_pe_1_0_2_U132 ( .A(npu_inst_pe_1_0_2_int_data_0_), .B(
        int_o_data_npu[40]), .Z(npu_inst_pe_1_0_2_N73) );
  AND2_X1 npu_inst_pe_1_0_2_U131 ( .A1(int_o_data_npu[40]), .A2(
        npu_inst_pe_1_0_2_int_data_0_), .ZN(npu_inst_pe_1_0_2_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_2_U130 ( .A(int_o_data_npu[40]), .B(
        npu_inst_pe_1_0_2_n11), .ZN(npu_inst_pe_1_0_2_N65) );
  OR2_X1 npu_inst_pe_1_0_2_U129 ( .A1(npu_inst_pe_1_0_2_n11), .A2(
        int_o_data_npu[40]), .ZN(npu_inst_pe_1_0_2_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_2_U128 ( .A(int_o_data_npu[42]), .B(
        npu_inst_pe_1_0_2_add_79_carry_2_), .Z(npu_inst_pe_1_0_2_N75) );
  AND2_X1 npu_inst_pe_1_0_2_U127 ( .A1(npu_inst_pe_1_0_2_add_79_carry_2_), 
        .A2(int_o_data_npu[42]), .ZN(npu_inst_pe_1_0_2_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_2_U126 ( .A(int_o_data_npu[43]), .B(
        npu_inst_pe_1_0_2_add_79_carry_3_), .Z(npu_inst_pe_1_0_2_N76) );
  AND2_X1 npu_inst_pe_1_0_2_U125 ( .A1(npu_inst_pe_1_0_2_add_79_carry_3_), 
        .A2(int_o_data_npu[43]), .ZN(npu_inst_pe_1_0_2_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_2_U124 ( .A(int_o_data_npu[44]), .B(
        npu_inst_pe_1_0_2_add_79_carry_4_), .Z(npu_inst_pe_1_0_2_N77) );
  AND2_X1 npu_inst_pe_1_0_2_U123 ( .A1(npu_inst_pe_1_0_2_add_79_carry_4_), 
        .A2(int_o_data_npu[44]), .ZN(npu_inst_pe_1_0_2_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_2_U122 ( .A(int_o_data_npu[45]), .B(
        npu_inst_pe_1_0_2_add_79_carry_5_), .Z(npu_inst_pe_1_0_2_N78) );
  AND2_X1 npu_inst_pe_1_0_2_U121 ( .A1(npu_inst_pe_1_0_2_add_79_carry_5_), 
        .A2(int_o_data_npu[45]), .ZN(npu_inst_pe_1_0_2_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_2_U120 ( .A(int_o_data_npu[46]), .B(
        npu_inst_pe_1_0_2_add_79_carry_6_), .Z(npu_inst_pe_1_0_2_N79) );
  AND2_X1 npu_inst_pe_1_0_2_U119 ( .A1(npu_inst_pe_1_0_2_add_79_carry_6_), 
        .A2(int_o_data_npu[46]), .ZN(npu_inst_pe_1_0_2_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_2_U118 ( .A(int_o_data_npu[47]), .B(
        npu_inst_pe_1_0_2_add_79_carry_7_), .Z(npu_inst_pe_1_0_2_N80) );
  XNOR2_X1 npu_inst_pe_1_0_2_U117 ( .A(npu_inst_pe_1_0_2_sub_77_carry_2_), .B(
        int_o_data_npu[42]), .ZN(npu_inst_pe_1_0_2_N67) );
  OR2_X1 npu_inst_pe_1_0_2_U116 ( .A1(int_o_data_npu[42]), .A2(
        npu_inst_pe_1_0_2_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_0_2_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_2_U115 ( .A(npu_inst_pe_1_0_2_sub_77_carry_3_), .B(
        int_o_data_npu[43]), .ZN(npu_inst_pe_1_0_2_N68) );
  OR2_X1 npu_inst_pe_1_0_2_U114 ( .A1(int_o_data_npu[43]), .A2(
        npu_inst_pe_1_0_2_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_0_2_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_2_U113 ( .A(npu_inst_pe_1_0_2_sub_77_carry_4_), .B(
        int_o_data_npu[44]), .ZN(npu_inst_pe_1_0_2_N69) );
  OR2_X1 npu_inst_pe_1_0_2_U112 ( .A1(int_o_data_npu[44]), .A2(
        npu_inst_pe_1_0_2_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_0_2_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_2_U111 ( .A(npu_inst_pe_1_0_2_sub_77_carry_5_), .B(
        int_o_data_npu[45]), .ZN(npu_inst_pe_1_0_2_N70) );
  OR2_X1 npu_inst_pe_1_0_2_U110 ( .A1(int_o_data_npu[45]), .A2(
        npu_inst_pe_1_0_2_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_0_2_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_2_U109 ( .A(npu_inst_pe_1_0_2_sub_77_carry_6_), .B(
        int_o_data_npu[46]), .ZN(npu_inst_pe_1_0_2_N71) );
  OR2_X1 npu_inst_pe_1_0_2_U108 ( .A1(int_o_data_npu[46]), .A2(
        npu_inst_pe_1_0_2_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_0_2_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_2_U107 ( .A(int_o_data_npu[47]), .B(
        npu_inst_pe_1_0_2_sub_77_carry_7_), .ZN(npu_inst_pe_1_0_2_N72) );
  INV_X1 npu_inst_pe_1_0_2_U106 ( .A(npu_inst_n62), .ZN(npu_inst_pe_1_0_2_n5)
         );
  INV_X1 npu_inst_pe_1_0_2_U105 ( .A(npu_inst_n42), .ZN(npu_inst_pe_1_0_2_n2)
         );
  AOI22_X1 npu_inst_pe_1_0_2_U104 ( .A1(npu_inst_int_data_y_1__2__0_), .A2(
        npu_inst_pe_1_0_2_n58), .B1(npu_inst_pe_1_0_2_n117), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_2_n57) );
  INV_X1 npu_inst_pe_1_0_2_U103 ( .A(npu_inst_pe_1_0_2_n57), .ZN(
        npu_inst_pe_1_0_2_n106) );
  AOI22_X1 npu_inst_pe_1_0_2_U102 ( .A1(npu_inst_int_data_y_1__2__0_), .A2(
        npu_inst_pe_1_0_2_n54), .B1(npu_inst_pe_1_0_2_n116), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_2_n53) );
  INV_X1 npu_inst_pe_1_0_2_U99 ( .A(npu_inst_pe_1_0_2_n53), .ZN(
        npu_inst_pe_1_0_2_n107) );
  AOI22_X1 npu_inst_pe_1_0_2_U98 ( .A1(npu_inst_int_data_y_1__2__0_), .A2(
        npu_inst_pe_1_0_2_n50), .B1(npu_inst_pe_1_0_2_n115), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_2_n49) );
  INV_X1 npu_inst_pe_1_0_2_U97 ( .A(npu_inst_pe_1_0_2_n49), .ZN(
        npu_inst_pe_1_0_2_n108) );
  AOI22_X1 npu_inst_pe_1_0_2_U96 ( .A1(npu_inst_int_data_y_1__2__0_), .A2(
        npu_inst_pe_1_0_2_n46), .B1(npu_inst_pe_1_0_2_n114), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_2_n45) );
  INV_X1 npu_inst_pe_1_0_2_U95 ( .A(npu_inst_pe_1_0_2_n45), .ZN(
        npu_inst_pe_1_0_2_n109) );
  AOI22_X1 npu_inst_pe_1_0_2_U94 ( .A1(npu_inst_int_data_y_1__2__0_), .A2(
        npu_inst_pe_1_0_2_n42), .B1(npu_inst_pe_1_0_2_n113), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_2_n41) );
  INV_X1 npu_inst_pe_1_0_2_U93 ( .A(npu_inst_pe_1_0_2_n41), .ZN(
        npu_inst_pe_1_0_2_n110) );
  AOI22_X1 npu_inst_pe_1_0_2_U92 ( .A1(npu_inst_int_data_y_1__2__1_), .A2(
        npu_inst_pe_1_0_2_n58), .B1(npu_inst_pe_1_0_2_n117), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_2_n59) );
  INV_X1 npu_inst_pe_1_0_2_U91 ( .A(npu_inst_pe_1_0_2_n59), .ZN(
        npu_inst_pe_1_0_2_n100) );
  AOI22_X1 npu_inst_pe_1_0_2_U90 ( .A1(npu_inst_int_data_y_1__2__1_), .A2(
        npu_inst_pe_1_0_2_n54), .B1(npu_inst_pe_1_0_2_n116), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_2_n55) );
  INV_X1 npu_inst_pe_1_0_2_U89 ( .A(npu_inst_pe_1_0_2_n55), .ZN(
        npu_inst_pe_1_0_2_n101) );
  AOI22_X1 npu_inst_pe_1_0_2_U88 ( .A1(npu_inst_int_data_y_1__2__1_), .A2(
        npu_inst_pe_1_0_2_n50), .B1(npu_inst_pe_1_0_2_n115), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_2_n51) );
  INV_X1 npu_inst_pe_1_0_2_U87 ( .A(npu_inst_pe_1_0_2_n51), .ZN(
        npu_inst_pe_1_0_2_n102) );
  AOI22_X1 npu_inst_pe_1_0_2_U86 ( .A1(npu_inst_int_data_y_1__2__1_), .A2(
        npu_inst_pe_1_0_2_n46), .B1(npu_inst_pe_1_0_2_n114), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_2_n47) );
  INV_X1 npu_inst_pe_1_0_2_U85 ( .A(npu_inst_pe_1_0_2_n47), .ZN(
        npu_inst_pe_1_0_2_n103) );
  AOI22_X1 npu_inst_pe_1_0_2_U84 ( .A1(npu_inst_int_data_y_1__2__1_), .A2(
        npu_inst_pe_1_0_2_n42), .B1(npu_inst_pe_1_0_2_n113), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_2_n43) );
  INV_X1 npu_inst_pe_1_0_2_U83 ( .A(npu_inst_pe_1_0_2_n43), .ZN(
        npu_inst_pe_1_0_2_n104) );
  AOI22_X1 npu_inst_pe_1_0_2_U82 ( .A1(npu_inst_pe_1_0_2_n38), .A2(
        npu_inst_int_data_y_1__2__1_), .B1(npu_inst_pe_1_0_2_n112), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_2_n39) );
  INV_X1 npu_inst_pe_1_0_2_U81 ( .A(npu_inst_pe_1_0_2_n39), .ZN(
        npu_inst_pe_1_0_2_n105) );
  NAND2_X1 npu_inst_pe_1_0_2_U80 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_2_n60), .ZN(npu_inst_pe_1_0_2_n74) );
  OAI21_X1 npu_inst_pe_1_0_2_U79 ( .B1(npu_inst_pe_1_0_2_n63), .B2(
        npu_inst_pe_1_0_2_n60), .A(npu_inst_pe_1_0_2_n74), .ZN(
        npu_inst_pe_1_0_2_n97) );
  NAND2_X1 npu_inst_pe_1_0_2_U78 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_2_n60), .ZN(npu_inst_pe_1_0_2_n73) );
  OAI21_X1 npu_inst_pe_1_0_2_U77 ( .B1(npu_inst_pe_1_0_2_n61), .B2(
        npu_inst_pe_1_0_2_n60), .A(npu_inst_pe_1_0_2_n73), .ZN(
        npu_inst_pe_1_0_2_n96) );
  NAND2_X1 npu_inst_pe_1_0_2_U76 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_2_n56), .ZN(npu_inst_pe_1_0_2_n72) );
  OAI21_X1 npu_inst_pe_1_0_2_U75 ( .B1(npu_inst_pe_1_0_2_n63), .B2(
        npu_inst_pe_1_0_2_n56), .A(npu_inst_pe_1_0_2_n72), .ZN(
        npu_inst_pe_1_0_2_n95) );
  NAND2_X1 npu_inst_pe_1_0_2_U74 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_2_n56), .ZN(npu_inst_pe_1_0_2_n71) );
  OAI21_X1 npu_inst_pe_1_0_2_U73 ( .B1(npu_inst_pe_1_0_2_n61), .B2(
        npu_inst_pe_1_0_2_n56), .A(npu_inst_pe_1_0_2_n71), .ZN(
        npu_inst_pe_1_0_2_n94) );
  NAND2_X1 npu_inst_pe_1_0_2_U72 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_2_n52), .ZN(npu_inst_pe_1_0_2_n70) );
  OAI21_X1 npu_inst_pe_1_0_2_U71 ( .B1(npu_inst_pe_1_0_2_n63), .B2(
        npu_inst_pe_1_0_2_n52), .A(npu_inst_pe_1_0_2_n70), .ZN(
        npu_inst_pe_1_0_2_n93) );
  NAND2_X1 npu_inst_pe_1_0_2_U70 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_2_n52), .ZN(npu_inst_pe_1_0_2_n69) );
  OAI21_X1 npu_inst_pe_1_0_2_U69 ( .B1(npu_inst_pe_1_0_2_n61), .B2(
        npu_inst_pe_1_0_2_n52), .A(npu_inst_pe_1_0_2_n69), .ZN(
        npu_inst_pe_1_0_2_n92) );
  NAND2_X1 npu_inst_pe_1_0_2_U68 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_2_n48), .ZN(npu_inst_pe_1_0_2_n68) );
  OAI21_X1 npu_inst_pe_1_0_2_U67 ( .B1(npu_inst_pe_1_0_2_n63), .B2(
        npu_inst_pe_1_0_2_n48), .A(npu_inst_pe_1_0_2_n68), .ZN(
        npu_inst_pe_1_0_2_n91) );
  NAND2_X1 npu_inst_pe_1_0_2_U66 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_2_n48), .ZN(npu_inst_pe_1_0_2_n67) );
  OAI21_X1 npu_inst_pe_1_0_2_U65 ( .B1(npu_inst_pe_1_0_2_n61), .B2(
        npu_inst_pe_1_0_2_n48), .A(npu_inst_pe_1_0_2_n67), .ZN(
        npu_inst_pe_1_0_2_n90) );
  NAND2_X1 npu_inst_pe_1_0_2_U64 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_2_n44), .ZN(npu_inst_pe_1_0_2_n66) );
  OAI21_X1 npu_inst_pe_1_0_2_U63 ( .B1(npu_inst_pe_1_0_2_n63), .B2(
        npu_inst_pe_1_0_2_n44), .A(npu_inst_pe_1_0_2_n66), .ZN(
        npu_inst_pe_1_0_2_n89) );
  NAND2_X1 npu_inst_pe_1_0_2_U62 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_2_n44), .ZN(npu_inst_pe_1_0_2_n65) );
  OAI21_X1 npu_inst_pe_1_0_2_U61 ( .B1(npu_inst_pe_1_0_2_n61), .B2(
        npu_inst_pe_1_0_2_n44), .A(npu_inst_pe_1_0_2_n65), .ZN(
        npu_inst_pe_1_0_2_n88) );
  NAND2_X1 npu_inst_pe_1_0_2_U60 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_2_n40), .ZN(npu_inst_pe_1_0_2_n64) );
  OAI21_X1 npu_inst_pe_1_0_2_U59 ( .B1(npu_inst_pe_1_0_2_n63), .B2(
        npu_inst_pe_1_0_2_n40), .A(npu_inst_pe_1_0_2_n64), .ZN(
        npu_inst_pe_1_0_2_n87) );
  NAND2_X1 npu_inst_pe_1_0_2_U58 ( .A1(npu_inst_pe_1_0_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_2_n40), .ZN(npu_inst_pe_1_0_2_n62) );
  OAI21_X1 npu_inst_pe_1_0_2_U57 ( .B1(npu_inst_pe_1_0_2_n61), .B2(
        npu_inst_pe_1_0_2_n40), .A(npu_inst_pe_1_0_2_n62), .ZN(
        npu_inst_pe_1_0_2_n86) );
  AOI22_X1 npu_inst_pe_1_0_2_U56 ( .A1(npu_inst_pe_1_0_2_n38), .A2(
        npu_inst_int_data_y_1__2__0_), .B1(npu_inst_pe_1_0_2_n112), .B2(
        npu_inst_pe_1_0_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_2_n37) );
  INV_X1 npu_inst_pe_1_0_2_U55 ( .A(npu_inst_pe_1_0_2_n37), .ZN(
        npu_inst_pe_1_0_2_n111) );
  AOI222_X1 npu_inst_pe_1_0_2_U54 ( .A1(npu_inst_int_data_res_1__2__0_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N73), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N65), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n84) );
  INV_X1 npu_inst_pe_1_0_2_U53 ( .A(npu_inst_pe_1_0_2_n84), .ZN(
        npu_inst_pe_1_0_2_n99) );
  AOI222_X1 npu_inst_pe_1_0_2_U52 ( .A1(npu_inst_pe_1_0_2_n1), .A2(
        npu_inst_int_data_res_1__2__7_), .B1(npu_inst_pe_1_0_2_N80), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N72), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n75) );
  INV_X1 npu_inst_pe_1_0_2_U51 ( .A(npu_inst_pe_1_0_2_n75), .ZN(
        npu_inst_pe_1_0_2_n31) );
  AOI222_X1 npu_inst_pe_1_0_2_U50 ( .A1(npu_inst_int_data_res_1__2__2_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N75), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N67), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n82) );
  INV_X1 npu_inst_pe_1_0_2_U49 ( .A(npu_inst_pe_1_0_2_n82), .ZN(
        npu_inst_pe_1_0_2_n36) );
  AOI222_X1 npu_inst_pe_1_0_2_U48 ( .A1(npu_inst_int_data_res_1__2__3_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N76), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N68), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n81) );
  INV_X1 npu_inst_pe_1_0_2_U47 ( .A(npu_inst_pe_1_0_2_n81), .ZN(
        npu_inst_pe_1_0_2_n35) );
  AOI222_X1 npu_inst_pe_1_0_2_U46 ( .A1(npu_inst_int_data_res_1__2__4_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N77), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N69), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n80) );
  INV_X1 npu_inst_pe_1_0_2_U45 ( .A(npu_inst_pe_1_0_2_n80), .ZN(
        npu_inst_pe_1_0_2_n34) );
  AOI222_X1 npu_inst_pe_1_0_2_U44 ( .A1(npu_inst_int_data_res_1__2__5_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N78), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N70), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n79) );
  INV_X1 npu_inst_pe_1_0_2_U43 ( .A(npu_inst_pe_1_0_2_n79), .ZN(
        npu_inst_pe_1_0_2_n33) );
  AOI222_X1 npu_inst_pe_1_0_2_U42 ( .A1(npu_inst_int_data_res_1__2__6_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N79), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N71), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n78) );
  INV_X1 npu_inst_pe_1_0_2_U41 ( .A(npu_inst_pe_1_0_2_n78), .ZN(
        npu_inst_pe_1_0_2_n32) );
  NOR3_X1 npu_inst_pe_1_0_2_U40 ( .A1(npu_inst_pe_1_0_2_n26), .A2(npu_inst_n42), .A3(npu_inst_int_ckg[61]), .ZN(npu_inst_pe_1_0_2_n85) );
  OR2_X1 npu_inst_pe_1_0_2_U39 ( .A1(npu_inst_pe_1_0_2_n85), .A2(
        npu_inst_pe_1_0_2_n1), .ZN(npu_inst_pe_1_0_2_N84) );
  AND2_X1 npu_inst_pe_1_0_2_U38 ( .A1(npu_inst_int_data_x_0__2__1_), .A2(
        npu_inst_pe_1_0_2_int_q_weight_1_), .ZN(npu_inst_pe_1_0_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_2_U37 ( .A1(npu_inst_int_data_x_0__2__0_), .A2(
        npu_inst_pe_1_0_2_int_q_weight_1_), .ZN(npu_inst_pe_1_0_2_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_0_2_U36 ( .A(npu_inst_pe_1_0_2_int_data_1_), .ZN(
        npu_inst_pe_1_0_2_n12) );
  AOI222_X1 npu_inst_pe_1_0_2_U35 ( .A1(npu_inst_int_data_res_1__2__1_), .A2(
        npu_inst_pe_1_0_2_n1), .B1(npu_inst_pe_1_0_2_N74), .B2(
        npu_inst_pe_1_0_2_n76), .C1(npu_inst_pe_1_0_2_N66), .C2(
        npu_inst_pe_1_0_2_n77), .ZN(npu_inst_pe_1_0_2_n83) );
  INV_X1 npu_inst_pe_1_0_2_U34 ( .A(npu_inst_pe_1_0_2_n83), .ZN(
        npu_inst_pe_1_0_2_n98) );
  AND2_X1 npu_inst_pe_1_0_2_U33 ( .A1(npu_inst_pe_1_0_2_N93), .A2(npu_inst_n42), .ZN(npu_inst_pe_1_0_2_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_2_U32 ( .A1(npu_inst_n42), .A2(npu_inst_pe_1_0_2_N94), .ZN(npu_inst_pe_1_0_2_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_2_U31 ( .A1(npu_inst_n42), .A2(
        npu_inst_int_data_y_1__2__1_), .B1(npu_inst_pe_1_0_2_n2), .B2(
        npu_inst_int_data_x_0__3__1_), .ZN(npu_inst_pe_1_0_2_n63) );
  AOI22_X1 npu_inst_pe_1_0_2_U30 ( .A1(npu_inst_n42), .A2(
        npu_inst_int_data_y_1__2__0_), .B1(npu_inst_pe_1_0_2_n2), .B2(
        npu_inst_int_data_x_0__3__0_), .ZN(npu_inst_pe_1_0_2_n61) );
  INV_X1 npu_inst_pe_1_0_2_U29 ( .A(npu_inst_pe_1_0_2_int_data_0_), .ZN(
        npu_inst_pe_1_0_2_n11) );
  INV_X1 npu_inst_pe_1_0_2_U28 ( .A(npu_inst_n54), .ZN(npu_inst_pe_1_0_2_n4)
         );
  OR3_X1 npu_inst_pe_1_0_2_U27 ( .A1(npu_inst_n62), .A2(npu_inst_pe_1_0_2_n6), 
        .A3(npu_inst_pe_1_0_2_n4), .ZN(npu_inst_pe_1_0_2_n56) );
  OR3_X1 npu_inst_pe_1_0_2_U26 ( .A1(npu_inst_pe_1_0_2_n4), .A2(
        npu_inst_pe_1_0_2_n6), .A3(npu_inst_pe_1_0_2_n5), .ZN(
        npu_inst_pe_1_0_2_n48) );
  INV_X1 npu_inst_pe_1_0_2_U25 ( .A(npu_inst_pe_1_0_2_n4), .ZN(
        npu_inst_pe_1_0_2_n3) );
  OR3_X1 npu_inst_pe_1_0_2_U24 ( .A1(npu_inst_pe_1_0_2_n3), .A2(
        npu_inst_pe_1_0_2_n6), .A3(npu_inst_pe_1_0_2_n5), .ZN(
        npu_inst_pe_1_0_2_n52) );
  OR3_X1 npu_inst_pe_1_0_2_U23 ( .A1(npu_inst_n62), .A2(npu_inst_pe_1_0_2_n6), 
        .A3(npu_inst_pe_1_0_2_n3), .ZN(npu_inst_pe_1_0_2_n60) );
  BUF_X1 npu_inst_pe_1_0_2_U22 ( .A(npu_inst_n31), .Z(npu_inst_pe_1_0_2_n1) );
  NOR2_X1 npu_inst_pe_1_0_2_U21 ( .A1(npu_inst_pe_1_0_2_n60), .A2(
        npu_inst_pe_1_0_2_n2), .ZN(npu_inst_pe_1_0_2_n58) );
  NOR2_X1 npu_inst_pe_1_0_2_U20 ( .A1(npu_inst_pe_1_0_2_n56), .A2(
        npu_inst_pe_1_0_2_n2), .ZN(npu_inst_pe_1_0_2_n54) );
  NOR2_X1 npu_inst_pe_1_0_2_U19 ( .A1(npu_inst_pe_1_0_2_n52), .A2(
        npu_inst_pe_1_0_2_n2), .ZN(npu_inst_pe_1_0_2_n50) );
  NOR2_X1 npu_inst_pe_1_0_2_U18 ( .A1(npu_inst_pe_1_0_2_n48), .A2(
        npu_inst_pe_1_0_2_n2), .ZN(npu_inst_pe_1_0_2_n46) );
  NOR2_X1 npu_inst_pe_1_0_2_U17 ( .A1(npu_inst_pe_1_0_2_n40), .A2(
        npu_inst_pe_1_0_2_n2), .ZN(npu_inst_pe_1_0_2_n38) );
  NOR2_X1 npu_inst_pe_1_0_2_U16 ( .A1(npu_inst_pe_1_0_2_n44), .A2(
        npu_inst_pe_1_0_2_n2), .ZN(npu_inst_pe_1_0_2_n42) );
  BUF_X1 npu_inst_pe_1_0_2_U15 ( .A(npu_inst_n89), .Z(npu_inst_pe_1_0_2_n6) );
  INV_X1 npu_inst_pe_1_0_2_U14 ( .A(npu_inst_n109), .ZN(npu_inst_pe_1_0_2_n10)
         );
  INV_X1 npu_inst_pe_1_0_2_U13 ( .A(npu_inst_pe_1_0_2_n38), .ZN(
        npu_inst_pe_1_0_2_n112) );
  INV_X1 npu_inst_pe_1_0_2_U12 ( .A(npu_inst_pe_1_0_2_n58), .ZN(
        npu_inst_pe_1_0_2_n117) );
  INV_X1 npu_inst_pe_1_0_2_U11 ( .A(npu_inst_pe_1_0_2_n54), .ZN(
        npu_inst_pe_1_0_2_n116) );
  INV_X1 npu_inst_pe_1_0_2_U10 ( .A(npu_inst_pe_1_0_2_n50), .ZN(
        npu_inst_pe_1_0_2_n115) );
  INV_X1 npu_inst_pe_1_0_2_U9 ( .A(npu_inst_pe_1_0_2_n46), .ZN(
        npu_inst_pe_1_0_2_n114) );
  INV_X1 npu_inst_pe_1_0_2_U8 ( .A(npu_inst_pe_1_0_2_n42), .ZN(
        npu_inst_pe_1_0_2_n113) );
  BUF_X1 npu_inst_pe_1_0_2_U7 ( .A(npu_inst_pe_1_0_2_n10), .Z(
        npu_inst_pe_1_0_2_n9) );
  BUF_X1 npu_inst_pe_1_0_2_U6 ( .A(npu_inst_pe_1_0_2_n10), .Z(
        npu_inst_pe_1_0_2_n8) );
  BUF_X1 npu_inst_pe_1_0_2_U5 ( .A(npu_inst_pe_1_0_2_n10), .Z(
        npu_inst_pe_1_0_2_n7) );
  NOR2_X1 npu_inst_pe_1_0_2_U4 ( .A1(npu_inst_pe_1_0_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_2_n1), .ZN(npu_inst_pe_1_0_2_n76) );
  NOR2_X1 npu_inst_pe_1_0_2_U3 ( .A1(npu_inst_pe_1_0_2_n27), .A2(
        npu_inst_pe_1_0_2_n1), .ZN(npu_inst_pe_1_0_2_n77) );
  FA_X1 npu_inst_pe_1_0_2_sub_77_U2_1 ( .A(int_o_data_npu[41]), .B(
        npu_inst_pe_1_0_2_n12), .CI(npu_inst_pe_1_0_2_sub_77_carry_1_), .CO(
        npu_inst_pe_1_0_2_sub_77_carry_2_), .S(npu_inst_pe_1_0_2_N66) );
  FA_X1 npu_inst_pe_1_0_2_add_79_U1_1 ( .A(int_o_data_npu[41]), .B(
        npu_inst_pe_1_0_2_int_data_1_), .CI(npu_inst_pe_1_0_2_add_79_carry_1_), 
        .CO(npu_inst_pe_1_0_2_add_79_carry_2_), .S(npu_inst_pe_1_0_2_N74) );
  NAND3_X1 npu_inst_pe_1_0_2_U101 ( .A1(npu_inst_pe_1_0_2_n4), .A2(
        npu_inst_pe_1_0_2_n5), .A3(npu_inst_pe_1_0_2_n6), .ZN(
        npu_inst_pe_1_0_2_n44) );
  NAND3_X1 npu_inst_pe_1_0_2_U100 ( .A1(npu_inst_pe_1_0_2_n3), .A2(
        npu_inst_pe_1_0_2_n5), .A3(npu_inst_pe_1_0_2_n6), .ZN(
        npu_inst_pe_1_0_2_n40) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_2_n32), .CK(
        npu_inst_pe_1_0_2_net4432), .RN(npu_inst_pe_1_0_2_n7), .Q(
        int_o_data_npu[46]) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_2_n33), .CK(
        npu_inst_pe_1_0_2_net4432), .RN(npu_inst_pe_1_0_2_n7), .Q(
        int_o_data_npu[45]) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_2_n34), .CK(
        npu_inst_pe_1_0_2_net4432), .RN(npu_inst_pe_1_0_2_n7), .Q(
        int_o_data_npu[44]) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_2_n35), .CK(
        npu_inst_pe_1_0_2_net4432), .RN(npu_inst_pe_1_0_2_n7), .Q(
        int_o_data_npu[43]) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_2_n36), .CK(
        npu_inst_pe_1_0_2_net4432), .RN(npu_inst_pe_1_0_2_n7), .Q(
        int_o_data_npu[42]) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_2_n98), .CK(
        npu_inst_pe_1_0_2_net4432), .RN(npu_inst_pe_1_0_2_n7), .Q(
        int_o_data_npu[41]) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_2_n31), .CK(
        npu_inst_pe_1_0_2_net4432), .RN(npu_inst_pe_1_0_2_n7), .Q(
        int_o_data_npu[47]) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_2_n99), .CK(
        npu_inst_pe_1_0_2_net4432), .RN(npu_inst_pe_1_0_2_n7), .Q(
        int_o_data_npu[40]) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_weight_reg_0_ ( .D(npu_inst_n95), .CK(
        npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n7), .Q(
        npu_inst_pe_1_0_2_int_q_weight_0_), .QN(npu_inst_pe_1_0_2_n27) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_weight_reg_1_ ( .D(npu_inst_n101), .CK(
        npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n7), .Q(
        npu_inst_pe_1_0_2_int_q_weight_1_), .QN(npu_inst_pe_1_0_2_n26) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_2_n111), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n7), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_2_n105), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n7), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_2_n110), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_2_n104), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_2_n109), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_2_n103), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_2_n108), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_2_n102), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_2_n107), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_2_n101), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_2_n106), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_2_n100), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_2_n86), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_2_n87), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n8), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_2_n88), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_2_n89), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_2_n90), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_2_n91), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_2_n92), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_2_n93), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_2_n94), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_2_n95), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_2_n96), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_2_n97), 
        .CK(npu_inst_pe_1_0_2_net4438), .RN(npu_inst_pe_1_0_2_n9), .Q(
        npu_inst_pe_1_0_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_2_net4432) );
  CLKGATETST_X1 npu_inst_pe_1_0_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n48), .SE(1'b0), .GCK(npu_inst_pe_1_0_2_net4438) );
  MUX2_X1 npu_inst_pe_1_0_3_U153 ( .A(npu_inst_pe_1_0_3_n31), .B(
        npu_inst_pe_1_0_3_n28), .S(npu_inst_pe_1_0_3_n7), .Z(
        npu_inst_pe_1_0_3_N93) );
  MUX2_X1 npu_inst_pe_1_0_3_U152 ( .A(npu_inst_pe_1_0_3_n30), .B(
        npu_inst_pe_1_0_3_n29), .S(npu_inst_pe_1_0_3_n5), .Z(
        npu_inst_pe_1_0_3_n31) );
  MUX2_X1 npu_inst_pe_1_0_3_U151 ( .A(npu_inst_pe_1_0_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_3_n3), .Z(
        npu_inst_pe_1_0_3_n30) );
  MUX2_X1 npu_inst_pe_1_0_3_U150 ( .A(npu_inst_pe_1_0_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_3_n3), .Z(
        npu_inst_pe_1_0_3_n29) );
  MUX2_X1 npu_inst_pe_1_0_3_U149 ( .A(npu_inst_pe_1_0_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_3_n3), .Z(
        npu_inst_pe_1_0_3_n28) );
  MUX2_X1 npu_inst_pe_1_0_3_U148 ( .A(npu_inst_pe_1_0_3_n25), .B(
        npu_inst_pe_1_0_3_n22), .S(npu_inst_pe_1_0_3_n7), .Z(
        npu_inst_pe_1_0_3_N94) );
  MUX2_X1 npu_inst_pe_1_0_3_U147 ( .A(npu_inst_pe_1_0_3_n24), .B(
        npu_inst_pe_1_0_3_n23), .S(npu_inst_pe_1_0_3_n5), .Z(
        npu_inst_pe_1_0_3_n25) );
  MUX2_X1 npu_inst_pe_1_0_3_U146 ( .A(npu_inst_pe_1_0_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_3_n3), .Z(
        npu_inst_pe_1_0_3_n24) );
  MUX2_X1 npu_inst_pe_1_0_3_U145 ( .A(npu_inst_pe_1_0_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_3_n3), .Z(
        npu_inst_pe_1_0_3_n23) );
  MUX2_X1 npu_inst_pe_1_0_3_U144 ( .A(npu_inst_pe_1_0_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_3_n3), .Z(
        npu_inst_pe_1_0_3_n22) );
  MUX2_X1 npu_inst_pe_1_0_3_U143 ( .A(npu_inst_pe_1_0_3_n21), .B(
        npu_inst_pe_1_0_3_n18), .S(npu_inst_pe_1_0_3_n7), .Z(
        npu_inst_int_data_x_0__3__1_) );
  MUX2_X1 npu_inst_pe_1_0_3_U142 ( .A(npu_inst_pe_1_0_3_n20), .B(
        npu_inst_pe_1_0_3_n19), .S(npu_inst_pe_1_0_3_n5), .Z(
        npu_inst_pe_1_0_3_n21) );
  MUX2_X1 npu_inst_pe_1_0_3_U141 ( .A(npu_inst_pe_1_0_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_3_n3), .Z(
        npu_inst_pe_1_0_3_n20) );
  MUX2_X1 npu_inst_pe_1_0_3_U140 ( .A(npu_inst_pe_1_0_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_3_n3), .Z(
        npu_inst_pe_1_0_3_n19) );
  MUX2_X1 npu_inst_pe_1_0_3_U139 ( .A(npu_inst_pe_1_0_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_3_n3), .Z(
        npu_inst_pe_1_0_3_n18) );
  MUX2_X1 npu_inst_pe_1_0_3_U138 ( .A(npu_inst_pe_1_0_3_n17), .B(
        npu_inst_pe_1_0_3_n14), .S(npu_inst_pe_1_0_3_n7), .Z(
        npu_inst_int_data_x_0__3__0_) );
  MUX2_X1 npu_inst_pe_1_0_3_U137 ( .A(npu_inst_pe_1_0_3_n16), .B(
        npu_inst_pe_1_0_3_n15), .S(npu_inst_pe_1_0_3_n5), .Z(
        npu_inst_pe_1_0_3_n17) );
  MUX2_X1 npu_inst_pe_1_0_3_U136 ( .A(npu_inst_pe_1_0_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_3_n3), .Z(
        npu_inst_pe_1_0_3_n16) );
  MUX2_X1 npu_inst_pe_1_0_3_U135 ( .A(npu_inst_pe_1_0_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_3_n3), .Z(
        npu_inst_pe_1_0_3_n15) );
  MUX2_X1 npu_inst_pe_1_0_3_U134 ( .A(npu_inst_pe_1_0_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_3_n3), .Z(
        npu_inst_pe_1_0_3_n14) );
  XOR2_X1 npu_inst_pe_1_0_3_U133 ( .A(npu_inst_pe_1_0_3_int_data_0_), .B(
        int_o_data_npu[32]), .Z(npu_inst_pe_1_0_3_N73) );
  AND2_X1 npu_inst_pe_1_0_3_U132 ( .A1(int_o_data_npu[32]), .A2(
        npu_inst_pe_1_0_3_int_data_0_), .ZN(npu_inst_pe_1_0_3_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_3_U131 ( .A(int_o_data_npu[32]), .B(
        npu_inst_pe_1_0_3_n12), .ZN(npu_inst_pe_1_0_3_N65) );
  OR2_X1 npu_inst_pe_1_0_3_U130 ( .A1(npu_inst_pe_1_0_3_n12), .A2(
        int_o_data_npu[32]), .ZN(npu_inst_pe_1_0_3_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_3_U129 ( .A(int_o_data_npu[34]), .B(
        npu_inst_pe_1_0_3_add_79_carry_2_), .Z(npu_inst_pe_1_0_3_N75) );
  AND2_X1 npu_inst_pe_1_0_3_U128 ( .A1(npu_inst_pe_1_0_3_add_79_carry_2_), 
        .A2(int_o_data_npu[34]), .ZN(npu_inst_pe_1_0_3_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_3_U127 ( .A(int_o_data_npu[35]), .B(
        npu_inst_pe_1_0_3_add_79_carry_3_), .Z(npu_inst_pe_1_0_3_N76) );
  AND2_X1 npu_inst_pe_1_0_3_U126 ( .A1(npu_inst_pe_1_0_3_add_79_carry_3_), 
        .A2(int_o_data_npu[35]), .ZN(npu_inst_pe_1_0_3_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_3_U125 ( .A(int_o_data_npu[36]), .B(
        npu_inst_pe_1_0_3_add_79_carry_4_), .Z(npu_inst_pe_1_0_3_N77) );
  AND2_X1 npu_inst_pe_1_0_3_U124 ( .A1(npu_inst_pe_1_0_3_add_79_carry_4_), 
        .A2(int_o_data_npu[36]), .ZN(npu_inst_pe_1_0_3_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_3_U123 ( .A(int_o_data_npu[37]), .B(
        npu_inst_pe_1_0_3_add_79_carry_5_), .Z(npu_inst_pe_1_0_3_N78) );
  AND2_X1 npu_inst_pe_1_0_3_U122 ( .A1(npu_inst_pe_1_0_3_add_79_carry_5_), 
        .A2(int_o_data_npu[37]), .ZN(npu_inst_pe_1_0_3_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_3_U121 ( .A(int_o_data_npu[38]), .B(
        npu_inst_pe_1_0_3_add_79_carry_6_), .Z(npu_inst_pe_1_0_3_N79) );
  AND2_X1 npu_inst_pe_1_0_3_U120 ( .A1(npu_inst_pe_1_0_3_add_79_carry_6_), 
        .A2(int_o_data_npu[38]), .ZN(npu_inst_pe_1_0_3_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_3_U119 ( .A(int_o_data_npu[39]), .B(
        npu_inst_pe_1_0_3_add_79_carry_7_), .Z(npu_inst_pe_1_0_3_N80) );
  XNOR2_X1 npu_inst_pe_1_0_3_U118 ( .A(npu_inst_pe_1_0_3_sub_77_carry_2_), .B(
        int_o_data_npu[34]), .ZN(npu_inst_pe_1_0_3_N67) );
  OR2_X1 npu_inst_pe_1_0_3_U117 ( .A1(int_o_data_npu[34]), .A2(
        npu_inst_pe_1_0_3_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_0_3_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_3_U116 ( .A(npu_inst_pe_1_0_3_sub_77_carry_3_), .B(
        int_o_data_npu[35]), .ZN(npu_inst_pe_1_0_3_N68) );
  OR2_X1 npu_inst_pe_1_0_3_U115 ( .A1(int_o_data_npu[35]), .A2(
        npu_inst_pe_1_0_3_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_0_3_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_3_U114 ( .A(npu_inst_pe_1_0_3_sub_77_carry_4_), .B(
        int_o_data_npu[36]), .ZN(npu_inst_pe_1_0_3_N69) );
  OR2_X1 npu_inst_pe_1_0_3_U113 ( .A1(int_o_data_npu[36]), .A2(
        npu_inst_pe_1_0_3_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_0_3_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_3_U112 ( .A(npu_inst_pe_1_0_3_sub_77_carry_5_), .B(
        int_o_data_npu[37]), .ZN(npu_inst_pe_1_0_3_N70) );
  OR2_X1 npu_inst_pe_1_0_3_U111 ( .A1(int_o_data_npu[37]), .A2(
        npu_inst_pe_1_0_3_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_0_3_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_3_U110 ( .A(npu_inst_pe_1_0_3_sub_77_carry_6_), .B(
        int_o_data_npu[38]), .ZN(npu_inst_pe_1_0_3_N71) );
  OR2_X1 npu_inst_pe_1_0_3_U109 ( .A1(int_o_data_npu[38]), .A2(
        npu_inst_pe_1_0_3_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_0_3_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_3_U108 ( .A(int_o_data_npu[39]), .B(
        npu_inst_pe_1_0_3_sub_77_carry_7_), .ZN(npu_inst_pe_1_0_3_N72) );
  INV_X1 npu_inst_pe_1_0_3_U107 ( .A(npu_inst_n62), .ZN(npu_inst_pe_1_0_3_n6)
         );
  INV_X1 npu_inst_pe_1_0_3_U106 ( .A(npu_inst_pe_1_0_3_n6), .ZN(
        npu_inst_pe_1_0_3_n5) );
  INV_X1 npu_inst_pe_1_0_3_U105 ( .A(npu_inst_n42), .ZN(npu_inst_pe_1_0_3_n2)
         );
  AOI22_X1 npu_inst_pe_1_0_3_U104 ( .A1(npu_inst_int_data_y_1__3__0_), .A2(
        npu_inst_pe_1_0_3_n58), .B1(npu_inst_pe_1_0_3_n118), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_3_n57) );
  INV_X1 npu_inst_pe_1_0_3_U103 ( .A(npu_inst_pe_1_0_3_n57), .ZN(
        npu_inst_pe_1_0_3_n107) );
  AOI22_X1 npu_inst_pe_1_0_3_U102 ( .A1(npu_inst_int_data_y_1__3__0_), .A2(
        npu_inst_pe_1_0_3_n54), .B1(npu_inst_pe_1_0_3_n117), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_3_n53) );
  INV_X1 npu_inst_pe_1_0_3_U99 ( .A(npu_inst_pe_1_0_3_n53), .ZN(
        npu_inst_pe_1_0_3_n108) );
  AOI22_X1 npu_inst_pe_1_0_3_U98 ( .A1(npu_inst_int_data_y_1__3__0_), .A2(
        npu_inst_pe_1_0_3_n50), .B1(npu_inst_pe_1_0_3_n116), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_3_n49) );
  INV_X1 npu_inst_pe_1_0_3_U97 ( .A(npu_inst_pe_1_0_3_n49), .ZN(
        npu_inst_pe_1_0_3_n109) );
  AOI22_X1 npu_inst_pe_1_0_3_U96 ( .A1(npu_inst_int_data_y_1__3__0_), .A2(
        npu_inst_pe_1_0_3_n46), .B1(npu_inst_pe_1_0_3_n115), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_3_n45) );
  INV_X1 npu_inst_pe_1_0_3_U95 ( .A(npu_inst_pe_1_0_3_n45), .ZN(
        npu_inst_pe_1_0_3_n110) );
  AOI22_X1 npu_inst_pe_1_0_3_U94 ( .A1(npu_inst_int_data_y_1__3__0_), .A2(
        npu_inst_pe_1_0_3_n42), .B1(npu_inst_pe_1_0_3_n114), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_3_n41) );
  INV_X1 npu_inst_pe_1_0_3_U93 ( .A(npu_inst_pe_1_0_3_n41), .ZN(
        npu_inst_pe_1_0_3_n111) );
  AOI22_X1 npu_inst_pe_1_0_3_U92 ( .A1(npu_inst_int_data_y_1__3__1_), .A2(
        npu_inst_pe_1_0_3_n58), .B1(npu_inst_pe_1_0_3_n118), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_3_n59) );
  INV_X1 npu_inst_pe_1_0_3_U91 ( .A(npu_inst_pe_1_0_3_n59), .ZN(
        npu_inst_pe_1_0_3_n101) );
  AOI22_X1 npu_inst_pe_1_0_3_U90 ( .A1(npu_inst_int_data_y_1__3__1_), .A2(
        npu_inst_pe_1_0_3_n54), .B1(npu_inst_pe_1_0_3_n117), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_3_n55) );
  INV_X1 npu_inst_pe_1_0_3_U89 ( .A(npu_inst_pe_1_0_3_n55), .ZN(
        npu_inst_pe_1_0_3_n102) );
  AOI22_X1 npu_inst_pe_1_0_3_U88 ( .A1(npu_inst_int_data_y_1__3__1_), .A2(
        npu_inst_pe_1_0_3_n50), .B1(npu_inst_pe_1_0_3_n116), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_3_n51) );
  INV_X1 npu_inst_pe_1_0_3_U87 ( .A(npu_inst_pe_1_0_3_n51), .ZN(
        npu_inst_pe_1_0_3_n103) );
  AOI22_X1 npu_inst_pe_1_0_3_U86 ( .A1(npu_inst_int_data_y_1__3__1_), .A2(
        npu_inst_pe_1_0_3_n46), .B1(npu_inst_pe_1_0_3_n115), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_3_n47) );
  INV_X1 npu_inst_pe_1_0_3_U85 ( .A(npu_inst_pe_1_0_3_n47), .ZN(
        npu_inst_pe_1_0_3_n104) );
  AOI22_X1 npu_inst_pe_1_0_3_U84 ( .A1(npu_inst_int_data_y_1__3__1_), .A2(
        npu_inst_pe_1_0_3_n42), .B1(npu_inst_pe_1_0_3_n114), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_3_n43) );
  INV_X1 npu_inst_pe_1_0_3_U83 ( .A(npu_inst_pe_1_0_3_n43), .ZN(
        npu_inst_pe_1_0_3_n105) );
  AOI22_X1 npu_inst_pe_1_0_3_U82 ( .A1(npu_inst_pe_1_0_3_n38), .A2(
        npu_inst_int_data_y_1__3__1_), .B1(npu_inst_pe_1_0_3_n113), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_3_n39) );
  INV_X1 npu_inst_pe_1_0_3_U81 ( .A(npu_inst_pe_1_0_3_n39), .ZN(
        npu_inst_pe_1_0_3_n106) );
  NAND2_X1 npu_inst_pe_1_0_3_U80 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_3_n60), .ZN(npu_inst_pe_1_0_3_n74) );
  OAI21_X1 npu_inst_pe_1_0_3_U79 ( .B1(npu_inst_pe_1_0_3_n63), .B2(
        npu_inst_pe_1_0_3_n60), .A(npu_inst_pe_1_0_3_n74), .ZN(
        npu_inst_pe_1_0_3_n97) );
  NAND2_X1 npu_inst_pe_1_0_3_U78 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_3_n60), .ZN(npu_inst_pe_1_0_3_n73) );
  OAI21_X1 npu_inst_pe_1_0_3_U77 ( .B1(npu_inst_pe_1_0_3_n61), .B2(
        npu_inst_pe_1_0_3_n60), .A(npu_inst_pe_1_0_3_n73), .ZN(
        npu_inst_pe_1_0_3_n96) );
  NAND2_X1 npu_inst_pe_1_0_3_U76 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_3_n56), .ZN(npu_inst_pe_1_0_3_n72) );
  OAI21_X1 npu_inst_pe_1_0_3_U75 ( .B1(npu_inst_pe_1_0_3_n63), .B2(
        npu_inst_pe_1_0_3_n56), .A(npu_inst_pe_1_0_3_n72), .ZN(
        npu_inst_pe_1_0_3_n95) );
  NAND2_X1 npu_inst_pe_1_0_3_U74 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_3_n56), .ZN(npu_inst_pe_1_0_3_n71) );
  OAI21_X1 npu_inst_pe_1_0_3_U73 ( .B1(npu_inst_pe_1_0_3_n61), .B2(
        npu_inst_pe_1_0_3_n56), .A(npu_inst_pe_1_0_3_n71), .ZN(
        npu_inst_pe_1_0_3_n94) );
  NAND2_X1 npu_inst_pe_1_0_3_U72 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_3_n52), .ZN(npu_inst_pe_1_0_3_n70) );
  OAI21_X1 npu_inst_pe_1_0_3_U71 ( .B1(npu_inst_pe_1_0_3_n63), .B2(
        npu_inst_pe_1_0_3_n52), .A(npu_inst_pe_1_0_3_n70), .ZN(
        npu_inst_pe_1_0_3_n93) );
  NAND2_X1 npu_inst_pe_1_0_3_U70 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_3_n52), .ZN(npu_inst_pe_1_0_3_n69) );
  OAI21_X1 npu_inst_pe_1_0_3_U69 ( .B1(npu_inst_pe_1_0_3_n61), .B2(
        npu_inst_pe_1_0_3_n52), .A(npu_inst_pe_1_0_3_n69), .ZN(
        npu_inst_pe_1_0_3_n92) );
  NAND2_X1 npu_inst_pe_1_0_3_U68 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_3_n48), .ZN(npu_inst_pe_1_0_3_n68) );
  OAI21_X1 npu_inst_pe_1_0_3_U67 ( .B1(npu_inst_pe_1_0_3_n63), .B2(
        npu_inst_pe_1_0_3_n48), .A(npu_inst_pe_1_0_3_n68), .ZN(
        npu_inst_pe_1_0_3_n91) );
  NAND2_X1 npu_inst_pe_1_0_3_U66 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_3_n48), .ZN(npu_inst_pe_1_0_3_n67) );
  OAI21_X1 npu_inst_pe_1_0_3_U65 ( .B1(npu_inst_pe_1_0_3_n61), .B2(
        npu_inst_pe_1_0_3_n48), .A(npu_inst_pe_1_0_3_n67), .ZN(
        npu_inst_pe_1_0_3_n90) );
  NAND2_X1 npu_inst_pe_1_0_3_U64 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_3_n44), .ZN(npu_inst_pe_1_0_3_n66) );
  OAI21_X1 npu_inst_pe_1_0_3_U63 ( .B1(npu_inst_pe_1_0_3_n63), .B2(
        npu_inst_pe_1_0_3_n44), .A(npu_inst_pe_1_0_3_n66), .ZN(
        npu_inst_pe_1_0_3_n89) );
  NAND2_X1 npu_inst_pe_1_0_3_U62 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_3_n44), .ZN(npu_inst_pe_1_0_3_n65) );
  OAI21_X1 npu_inst_pe_1_0_3_U61 ( .B1(npu_inst_pe_1_0_3_n61), .B2(
        npu_inst_pe_1_0_3_n44), .A(npu_inst_pe_1_0_3_n65), .ZN(
        npu_inst_pe_1_0_3_n88) );
  NAND2_X1 npu_inst_pe_1_0_3_U60 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_3_n40), .ZN(npu_inst_pe_1_0_3_n64) );
  OAI21_X1 npu_inst_pe_1_0_3_U59 ( .B1(npu_inst_pe_1_0_3_n63), .B2(
        npu_inst_pe_1_0_3_n40), .A(npu_inst_pe_1_0_3_n64), .ZN(
        npu_inst_pe_1_0_3_n87) );
  NAND2_X1 npu_inst_pe_1_0_3_U58 ( .A1(npu_inst_pe_1_0_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_3_n40), .ZN(npu_inst_pe_1_0_3_n62) );
  OAI21_X1 npu_inst_pe_1_0_3_U57 ( .B1(npu_inst_pe_1_0_3_n61), .B2(
        npu_inst_pe_1_0_3_n40), .A(npu_inst_pe_1_0_3_n62), .ZN(
        npu_inst_pe_1_0_3_n86) );
  AOI22_X1 npu_inst_pe_1_0_3_U56 ( .A1(npu_inst_pe_1_0_3_n38), .A2(
        npu_inst_int_data_y_1__3__0_), .B1(npu_inst_pe_1_0_3_n113), .B2(
        npu_inst_pe_1_0_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_3_n37) );
  INV_X1 npu_inst_pe_1_0_3_U55 ( .A(npu_inst_pe_1_0_3_n37), .ZN(
        npu_inst_pe_1_0_3_n112) );
  AOI222_X1 npu_inst_pe_1_0_3_U54 ( .A1(npu_inst_int_data_res_1__3__0_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N73), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N65), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n84) );
  INV_X1 npu_inst_pe_1_0_3_U53 ( .A(npu_inst_pe_1_0_3_n84), .ZN(
        npu_inst_pe_1_0_3_n100) );
  AOI222_X1 npu_inst_pe_1_0_3_U52 ( .A1(npu_inst_pe_1_0_3_n1), .A2(
        npu_inst_int_data_res_1__3__7_), .B1(npu_inst_pe_1_0_3_N80), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N72), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n75) );
  INV_X1 npu_inst_pe_1_0_3_U51 ( .A(npu_inst_pe_1_0_3_n75), .ZN(
        npu_inst_pe_1_0_3_n32) );
  AOI222_X1 npu_inst_pe_1_0_3_U50 ( .A1(npu_inst_int_data_res_1__3__2_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N75), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N67), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n82) );
  INV_X1 npu_inst_pe_1_0_3_U49 ( .A(npu_inst_pe_1_0_3_n82), .ZN(
        npu_inst_pe_1_0_3_n98) );
  AOI222_X1 npu_inst_pe_1_0_3_U48 ( .A1(npu_inst_int_data_res_1__3__3_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N76), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N68), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n81) );
  INV_X1 npu_inst_pe_1_0_3_U47 ( .A(npu_inst_pe_1_0_3_n81), .ZN(
        npu_inst_pe_1_0_3_n36) );
  AOI222_X1 npu_inst_pe_1_0_3_U46 ( .A1(npu_inst_int_data_res_1__3__4_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N77), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N69), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n80) );
  INV_X1 npu_inst_pe_1_0_3_U45 ( .A(npu_inst_pe_1_0_3_n80), .ZN(
        npu_inst_pe_1_0_3_n35) );
  AOI222_X1 npu_inst_pe_1_0_3_U44 ( .A1(npu_inst_int_data_res_1__3__5_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N78), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N70), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n79) );
  INV_X1 npu_inst_pe_1_0_3_U43 ( .A(npu_inst_pe_1_0_3_n79), .ZN(
        npu_inst_pe_1_0_3_n34) );
  AOI222_X1 npu_inst_pe_1_0_3_U42 ( .A1(npu_inst_int_data_res_1__3__6_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N79), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N71), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n78) );
  INV_X1 npu_inst_pe_1_0_3_U41 ( .A(npu_inst_pe_1_0_3_n78), .ZN(
        npu_inst_pe_1_0_3_n33) );
  NOR3_X1 npu_inst_pe_1_0_3_U40 ( .A1(npu_inst_pe_1_0_3_n26), .A2(npu_inst_n42), .A3(npu_inst_int_ckg[60]), .ZN(npu_inst_pe_1_0_3_n85) );
  OR2_X1 npu_inst_pe_1_0_3_U39 ( .A1(npu_inst_pe_1_0_3_n85), .A2(
        npu_inst_pe_1_0_3_n1), .ZN(npu_inst_pe_1_0_3_N84) );
  AND2_X1 npu_inst_pe_1_0_3_U38 ( .A1(npu_inst_int_data_x_0__3__1_), .A2(
        npu_inst_pe_1_0_3_int_q_weight_1_), .ZN(npu_inst_pe_1_0_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_3_U37 ( .A1(npu_inst_int_data_x_0__3__0_), .A2(
        npu_inst_pe_1_0_3_int_q_weight_1_), .ZN(npu_inst_pe_1_0_3_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_0_3_U36 ( .A(npu_inst_pe_1_0_3_int_data_1_), .ZN(
        npu_inst_pe_1_0_3_n13) );
  AOI222_X1 npu_inst_pe_1_0_3_U35 ( .A1(npu_inst_int_data_res_1__3__1_), .A2(
        npu_inst_pe_1_0_3_n1), .B1(npu_inst_pe_1_0_3_N74), .B2(
        npu_inst_pe_1_0_3_n76), .C1(npu_inst_pe_1_0_3_N66), .C2(
        npu_inst_pe_1_0_3_n77), .ZN(npu_inst_pe_1_0_3_n83) );
  INV_X1 npu_inst_pe_1_0_3_U34 ( .A(npu_inst_pe_1_0_3_n83), .ZN(
        npu_inst_pe_1_0_3_n99) );
  AND2_X1 npu_inst_pe_1_0_3_U33 ( .A1(npu_inst_pe_1_0_3_N93), .A2(npu_inst_n42), .ZN(npu_inst_pe_1_0_3_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_3_U32 ( .A1(npu_inst_n42), .A2(npu_inst_pe_1_0_3_N94), .ZN(npu_inst_pe_1_0_3_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_3_U31 ( .A1(npu_inst_n42), .A2(
        npu_inst_int_data_y_1__3__1_), .B1(npu_inst_pe_1_0_3_n2), .B2(
        npu_inst_int_data_x_0__4__1_), .ZN(npu_inst_pe_1_0_3_n63) );
  AOI22_X1 npu_inst_pe_1_0_3_U30 ( .A1(npu_inst_n42), .A2(
        npu_inst_int_data_y_1__3__0_), .B1(npu_inst_pe_1_0_3_n2), .B2(
        npu_inst_int_data_x_0__4__0_), .ZN(npu_inst_pe_1_0_3_n61) );
  INV_X1 npu_inst_pe_1_0_3_U29 ( .A(npu_inst_pe_1_0_3_int_data_0_), .ZN(
        npu_inst_pe_1_0_3_n12) );
  INV_X1 npu_inst_pe_1_0_3_U28 ( .A(npu_inst_n54), .ZN(npu_inst_pe_1_0_3_n4)
         );
  OR3_X1 npu_inst_pe_1_0_3_U27 ( .A1(npu_inst_pe_1_0_3_n5), .A2(
        npu_inst_pe_1_0_3_n7), .A3(npu_inst_pe_1_0_3_n4), .ZN(
        npu_inst_pe_1_0_3_n56) );
  OR3_X1 npu_inst_pe_1_0_3_U26 ( .A1(npu_inst_pe_1_0_3_n4), .A2(
        npu_inst_pe_1_0_3_n7), .A3(npu_inst_pe_1_0_3_n6), .ZN(
        npu_inst_pe_1_0_3_n48) );
  INV_X1 npu_inst_pe_1_0_3_U25 ( .A(npu_inst_pe_1_0_3_n4), .ZN(
        npu_inst_pe_1_0_3_n3) );
  OR3_X1 npu_inst_pe_1_0_3_U24 ( .A1(npu_inst_pe_1_0_3_n3), .A2(
        npu_inst_pe_1_0_3_n7), .A3(npu_inst_pe_1_0_3_n6), .ZN(
        npu_inst_pe_1_0_3_n52) );
  OR3_X1 npu_inst_pe_1_0_3_U23 ( .A1(npu_inst_pe_1_0_3_n5), .A2(
        npu_inst_pe_1_0_3_n7), .A3(npu_inst_pe_1_0_3_n3), .ZN(
        npu_inst_pe_1_0_3_n60) );
  BUF_X1 npu_inst_pe_1_0_3_U22 ( .A(npu_inst_n31), .Z(npu_inst_pe_1_0_3_n1) );
  NOR2_X1 npu_inst_pe_1_0_3_U21 ( .A1(npu_inst_pe_1_0_3_n60), .A2(
        npu_inst_pe_1_0_3_n2), .ZN(npu_inst_pe_1_0_3_n58) );
  NOR2_X1 npu_inst_pe_1_0_3_U20 ( .A1(npu_inst_pe_1_0_3_n56), .A2(
        npu_inst_pe_1_0_3_n2), .ZN(npu_inst_pe_1_0_3_n54) );
  NOR2_X1 npu_inst_pe_1_0_3_U19 ( .A1(npu_inst_pe_1_0_3_n52), .A2(
        npu_inst_pe_1_0_3_n2), .ZN(npu_inst_pe_1_0_3_n50) );
  NOR2_X1 npu_inst_pe_1_0_3_U18 ( .A1(npu_inst_pe_1_0_3_n48), .A2(
        npu_inst_pe_1_0_3_n2), .ZN(npu_inst_pe_1_0_3_n46) );
  NOR2_X1 npu_inst_pe_1_0_3_U17 ( .A1(npu_inst_pe_1_0_3_n40), .A2(
        npu_inst_pe_1_0_3_n2), .ZN(npu_inst_pe_1_0_3_n38) );
  NOR2_X1 npu_inst_pe_1_0_3_U16 ( .A1(npu_inst_pe_1_0_3_n44), .A2(
        npu_inst_pe_1_0_3_n2), .ZN(npu_inst_pe_1_0_3_n42) );
  BUF_X1 npu_inst_pe_1_0_3_U15 ( .A(npu_inst_n89), .Z(npu_inst_pe_1_0_3_n7) );
  INV_X1 npu_inst_pe_1_0_3_U14 ( .A(npu_inst_n109), .ZN(npu_inst_pe_1_0_3_n11)
         );
  INV_X1 npu_inst_pe_1_0_3_U13 ( .A(npu_inst_pe_1_0_3_n38), .ZN(
        npu_inst_pe_1_0_3_n113) );
  INV_X1 npu_inst_pe_1_0_3_U12 ( .A(npu_inst_pe_1_0_3_n58), .ZN(
        npu_inst_pe_1_0_3_n118) );
  INV_X1 npu_inst_pe_1_0_3_U11 ( .A(npu_inst_pe_1_0_3_n54), .ZN(
        npu_inst_pe_1_0_3_n117) );
  INV_X1 npu_inst_pe_1_0_3_U10 ( .A(npu_inst_pe_1_0_3_n50), .ZN(
        npu_inst_pe_1_0_3_n116) );
  INV_X1 npu_inst_pe_1_0_3_U9 ( .A(npu_inst_pe_1_0_3_n46), .ZN(
        npu_inst_pe_1_0_3_n115) );
  INV_X1 npu_inst_pe_1_0_3_U8 ( .A(npu_inst_pe_1_0_3_n42), .ZN(
        npu_inst_pe_1_0_3_n114) );
  BUF_X1 npu_inst_pe_1_0_3_U7 ( .A(npu_inst_pe_1_0_3_n11), .Z(
        npu_inst_pe_1_0_3_n10) );
  BUF_X1 npu_inst_pe_1_0_3_U6 ( .A(npu_inst_pe_1_0_3_n11), .Z(
        npu_inst_pe_1_0_3_n9) );
  BUF_X1 npu_inst_pe_1_0_3_U5 ( .A(npu_inst_pe_1_0_3_n11), .Z(
        npu_inst_pe_1_0_3_n8) );
  NOR2_X1 npu_inst_pe_1_0_3_U4 ( .A1(npu_inst_pe_1_0_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_3_n1), .ZN(npu_inst_pe_1_0_3_n76) );
  NOR2_X1 npu_inst_pe_1_0_3_U3 ( .A1(npu_inst_pe_1_0_3_n27), .A2(
        npu_inst_pe_1_0_3_n1), .ZN(npu_inst_pe_1_0_3_n77) );
  FA_X1 npu_inst_pe_1_0_3_sub_77_U2_1 ( .A(int_o_data_npu[33]), .B(
        npu_inst_pe_1_0_3_n13), .CI(npu_inst_pe_1_0_3_sub_77_carry_1_), .CO(
        npu_inst_pe_1_0_3_sub_77_carry_2_), .S(npu_inst_pe_1_0_3_N66) );
  FA_X1 npu_inst_pe_1_0_3_add_79_U1_1 ( .A(int_o_data_npu[33]), .B(
        npu_inst_pe_1_0_3_int_data_1_), .CI(npu_inst_pe_1_0_3_add_79_carry_1_), 
        .CO(npu_inst_pe_1_0_3_add_79_carry_2_), .S(npu_inst_pe_1_0_3_N74) );
  NAND3_X1 npu_inst_pe_1_0_3_U101 ( .A1(npu_inst_pe_1_0_3_n4), .A2(
        npu_inst_pe_1_0_3_n6), .A3(npu_inst_pe_1_0_3_n7), .ZN(
        npu_inst_pe_1_0_3_n44) );
  NAND3_X1 npu_inst_pe_1_0_3_U100 ( .A1(npu_inst_pe_1_0_3_n3), .A2(
        npu_inst_pe_1_0_3_n6), .A3(npu_inst_pe_1_0_3_n7), .ZN(
        npu_inst_pe_1_0_3_n40) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_3_n33), .CK(
        npu_inst_pe_1_0_3_net4409), .RN(npu_inst_pe_1_0_3_n8), .Q(
        int_o_data_npu[38]) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_3_n34), .CK(
        npu_inst_pe_1_0_3_net4409), .RN(npu_inst_pe_1_0_3_n8), .Q(
        int_o_data_npu[37]) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_3_n35), .CK(
        npu_inst_pe_1_0_3_net4409), .RN(npu_inst_pe_1_0_3_n8), .Q(
        int_o_data_npu[36]) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_3_n36), .CK(
        npu_inst_pe_1_0_3_net4409), .RN(npu_inst_pe_1_0_3_n8), .Q(
        int_o_data_npu[35]) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_3_n98), .CK(
        npu_inst_pe_1_0_3_net4409), .RN(npu_inst_pe_1_0_3_n8), .Q(
        int_o_data_npu[34]) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_3_n99), .CK(
        npu_inst_pe_1_0_3_net4409), .RN(npu_inst_pe_1_0_3_n8), .Q(
        int_o_data_npu[33]) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_3_n32), .CK(
        npu_inst_pe_1_0_3_net4409), .RN(npu_inst_pe_1_0_3_n8), .Q(
        int_o_data_npu[39]) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_3_n100), 
        .CK(npu_inst_pe_1_0_3_net4409), .RN(npu_inst_pe_1_0_3_n8), .Q(
        int_o_data_npu[32]) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_weight_reg_0_ ( .D(npu_inst_n95), .CK(
        npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n8), .Q(
        npu_inst_pe_1_0_3_int_q_weight_0_), .QN(npu_inst_pe_1_0_3_n27) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_weight_reg_1_ ( .D(npu_inst_n101), .CK(
        npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n8), .Q(
        npu_inst_pe_1_0_3_int_q_weight_1_), .QN(npu_inst_pe_1_0_3_n26) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_3_n112), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n8), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_3_n106), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n8), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_3_n111), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_3_n105), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_3_n110), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_3_n104), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_3_n109), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_3_n103), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_3_n108), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_3_n102), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_3_n107), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_3_n101), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_3_n86), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_3_n87), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n9), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_3_n88), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_3_n89), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_3_n90), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_3_n91), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_3_n92), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_3_n93), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_3_n94), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_3_n95), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_3_n96), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_3_n97), 
        .CK(npu_inst_pe_1_0_3_net4415), .RN(npu_inst_pe_1_0_3_n10), .Q(
        npu_inst_pe_1_0_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_3_net4409) );
  CLKGATETST_X1 npu_inst_pe_1_0_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n48), .SE(1'b0), .GCK(npu_inst_pe_1_0_3_net4415) );
  MUX2_X1 npu_inst_pe_1_0_4_U152 ( .A(npu_inst_pe_1_0_4_n30), .B(
        npu_inst_pe_1_0_4_n25), .S(npu_inst_pe_1_0_4_n6), .Z(
        npu_inst_pe_1_0_4_N93) );
  MUX2_X1 npu_inst_pe_1_0_4_U151 ( .A(npu_inst_pe_1_0_4_n29), .B(
        npu_inst_pe_1_0_4_n28), .S(npu_inst_n61), .Z(npu_inst_pe_1_0_4_n30) );
  MUX2_X1 npu_inst_pe_1_0_4_U150 ( .A(npu_inst_pe_1_0_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_4_n3), .Z(
        npu_inst_pe_1_0_4_n29) );
  MUX2_X1 npu_inst_pe_1_0_4_U149 ( .A(npu_inst_pe_1_0_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_4_n3), .Z(
        npu_inst_pe_1_0_4_n28) );
  MUX2_X1 npu_inst_pe_1_0_4_U148 ( .A(npu_inst_pe_1_0_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_4_n3), .Z(
        npu_inst_pe_1_0_4_n25) );
  MUX2_X1 npu_inst_pe_1_0_4_U147 ( .A(npu_inst_pe_1_0_4_n24), .B(
        npu_inst_pe_1_0_4_n21), .S(npu_inst_pe_1_0_4_n6), .Z(
        npu_inst_pe_1_0_4_N94) );
  MUX2_X1 npu_inst_pe_1_0_4_U146 ( .A(npu_inst_pe_1_0_4_n23), .B(
        npu_inst_pe_1_0_4_n22), .S(npu_inst_n61), .Z(npu_inst_pe_1_0_4_n24) );
  MUX2_X1 npu_inst_pe_1_0_4_U145 ( .A(npu_inst_pe_1_0_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_4_n3), .Z(
        npu_inst_pe_1_0_4_n23) );
  MUX2_X1 npu_inst_pe_1_0_4_U144 ( .A(npu_inst_pe_1_0_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_4_n3), .Z(
        npu_inst_pe_1_0_4_n22) );
  MUX2_X1 npu_inst_pe_1_0_4_U143 ( .A(npu_inst_pe_1_0_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_4_n3), .Z(
        npu_inst_pe_1_0_4_n21) );
  MUX2_X1 npu_inst_pe_1_0_4_U142 ( .A(npu_inst_pe_1_0_4_n20), .B(
        npu_inst_pe_1_0_4_n17), .S(npu_inst_pe_1_0_4_n6), .Z(
        npu_inst_int_data_x_0__4__1_) );
  MUX2_X1 npu_inst_pe_1_0_4_U141 ( .A(npu_inst_pe_1_0_4_n19), .B(
        npu_inst_pe_1_0_4_n18), .S(npu_inst_n61), .Z(npu_inst_pe_1_0_4_n20) );
  MUX2_X1 npu_inst_pe_1_0_4_U140 ( .A(npu_inst_pe_1_0_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_4_n3), .Z(
        npu_inst_pe_1_0_4_n19) );
  MUX2_X1 npu_inst_pe_1_0_4_U139 ( .A(npu_inst_pe_1_0_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_4_n3), .Z(
        npu_inst_pe_1_0_4_n18) );
  MUX2_X1 npu_inst_pe_1_0_4_U138 ( .A(npu_inst_pe_1_0_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_4_n3), .Z(
        npu_inst_pe_1_0_4_n17) );
  MUX2_X1 npu_inst_pe_1_0_4_U137 ( .A(npu_inst_pe_1_0_4_n16), .B(
        npu_inst_pe_1_0_4_n13), .S(npu_inst_pe_1_0_4_n6), .Z(
        npu_inst_int_data_x_0__4__0_) );
  MUX2_X1 npu_inst_pe_1_0_4_U136 ( .A(npu_inst_pe_1_0_4_n15), .B(
        npu_inst_pe_1_0_4_n14), .S(npu_inst_n61), .Z(npu_inst_pe_1_0_4_n16) );
  MUX2_X1 npu_inst_pe_1_0_4_U135 ( .A(npu_inst_pe_1_0_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_4_n3), .Z(
        npu_inst_pe_1_0_4_n15) );
  MUX2_X1 npu_inst_pe_1_0_4_U134 ( .A(npu_inst_pe_1_0_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_4_n3), .Z(
        npu_inst_pe_1_0_4_n14) );
  MUX2_X1 npu_inst_pe_1_0_4_U133 ( .A(npu_inst_pe_1_0_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_4_n3), .Z(
        npu_inst_pe_1_0_4_n13) );
  XOR2_X1 npu_inst_pe_1_0_4_U132 ( .A(npu_inst_pe_1_0_4_int_data_0_), .B(
        int_o_data_npu[24]), .Z(npu_inst_pe_1_0_4_N73) );
  AND2_X1 npu_inst_pe_1_0_4_U131 ( .A1(int_o_data_npu[24]), .A2(
        npu_inst_pe_1_0_4_int_data_0_), .ZN(npu_inst_pe_1_0_4_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_4_U130 ( .A(int_o_data_npu[24]), .B(
        npu_inst_pe_1_0_4_n11), .ZN(npu_inst_pe_1_0_4_N65) );
  OR2_X1 npu_inst_pe_1_0_4_U129 ( .A1(npu_inst_pe_1_0_4_n11), .A2(
        int_o_data_npu[24]), .ZN(npu_inst_pe_1_0_4_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_4_U128 ( .A(int_o_data_npu[26]), .B(
        npu_inst_pe_1_0_4_add_79_carry_2_), .Z(npu_inst_pe_1_0_4_N75) );
  AND2_X1 npu_inst_pe_1_0_4_U127 ( .A1(npu_inst_pe_1_0_4_add_79_carry_2_), 
        .A2(int_o_data_npu[26]), .ZN(npu_inst_pe_1_0_4_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_4_U126 ( .A(int_o_data_npu[27]), .B(
        npu_inst_pe_1_0_4_add_79_carry_3_), .Z(npu_inst_pe_1_0_4_N76) );
  AND2_X1 npu_inst_pe_1_0_4_U125 ( .A1(npu_inst_pe_1_0_4_add_79_carry_3_), 
        .A2(int_o_data_npu[27]), .ZN(npu_inst_pe_1_0_4_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_4_U124 ( .A(int_o_data_npu[28]), .B(
        npu_inst_pe_1_0_4_add_79_carry_4_), .Z(npu_inst_pe_1_0_4_N77) );
  AND2_X1 npu_inst_pe_1_0_4_U123 ( .A1(npu_inst_pe_1_0_4_add_79_carry_4_), 
        .A2(int_o_data_npu[28]), .ZN(npu_inst_pe_1_0_4_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_4_U122 ( .A(int_o_data_npu[29]), .B(
        npu_inst_pe_1_0_4_add_79_carry_5_), .Z(npu_inst_pe_1_0_4_N78) );
  AND2_X1 npu_inst_pe_1_0_4_U121 ( .A1(npu_inst_pe_1_0_4_add_79_carry_5_), 
        .A2(int_o_data_npu[29]), .ZN(npu_inst_pe_1_0_4_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_4_U120 ( .A(int_o_data_npu[30]), .B(
        npu_inst_pe_1_0_4_add_79_carry_6_), .Z(npu_inst_pe_1_0_4_N79) );
  AND2_X1 npu_inst_pe_1_0_4_U119 ( .A1(npu_inst_pe_1_0_4_add_79_carry_6_), 
        .A2(int_o_data_npu[30]), .ZN(npu_inst_pe_1_0_4_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_4_U118 ( .A(int_o_data_npu[31]), .B(
        npu_inst_pe_1_0_4_add_79_carry_7_), .Z(npu_inst_pe_1_0_4_N80) );
  XNOR2_X1 npu_inst_pe_1_0_4_U117 ( .A(npu_inst_pe_1_0_4_sub_77_carry_2_), .B(
        int_o_data_npu[26]), .ZN(npu_inst_pe_1_0_4_N67) );
  OR2_X1 npu_inst_pe_1_0_4_U116 ( .A1(int_o_data_npu[26]), .A2(
        npu_inst_pe_1_0_4_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_0_4_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_4_U115 ( .A(npu_inst_pe_1_0_4_sub_77_carry_3_), .B(
        int_o_data_npu[27]), .ZN(npu_inst_pe_1_0_4_N68) );
  OR2_X1 npu_inst_pe_1_0_4_U114 ( .A1(int_o_data_npu[27]), .A2(
        npu_inst_pe_1_0_4_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_0_4_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_4_U113 ( .A(npu_inst_pe_1_0_4_sub_77_carry_4_), .B(
        int_o_data_npu[28]), .ZN(npu_inst_pe_1_0_4_N69) );
  OR2_X1 npu_inst_pe_1_0_4_U112 ( .A1(int_o_data_npu[28]), .A2(
        npu_inst_pe_1_0_4_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_0_4_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_4_U111 ( .A(npu_inst_pe_1_0_4_sub_77_carry_5_), .B(
        int_o_data_npu[29]), .ZN(npu_inst_pe_1_0_4_N70) );
  OR2_X1 npu_inst_pe_1_0_4_U110 ( .A1(int_o_data_npu[29]), .A2(
        npu_inst_pe_1_0_4_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_0_4_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_4_U109 ( .A(npu_inst_pe_1_0_4_sub_77_carry_6_), .B(
        int_o_data_npu[30]), .ZN(npu_inst_pe_1_0_4_N71) );
  OR2_X1 npu_inst_pe_1_0_4_U108 ( .A1(int_o_data_npu[30]), .A2(
        npu_inst_pe_1_0_4_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_0_4_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_4_U107 ( .A(int_o_data_npu[31]), .B(
        npu_inst_pe_1_0_4_sub_77_carry_7_), .ZN(npu_inst_pe_1_0_4_N72) );
  INV_X1 npu_inst_pe_1_0_4_U106 ( .A(npu_inst_n61), .ZN(npu_inst_pe_1_0_4_n5)
         );
  INV_X1 npu_inst_pe_1_0_4_U105 ( .A(npu_inst_n42), .ZN(npu_inst_pe_1_0_4_n2)
         );
  AOI22_X1 npu_inst_pe_1_0_4_U104 ( .A1(npu_inst_int_data_y_1__4__0_), .A2(
        npu_inst_pe_1_0_4_n58), .B1(npu_inst_pe_1_0_4_n117), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_4_n57) );
  INV_X1 npu_inst_pe_1_0_4_U103 ( .A(npu_inst_pe_1_0_4_n57), .ZN(
        npu_inst_pe_1_0_4_n106) );
  AOI22_X1 npu_inst_pe_1_0_4_U102 ( .A1(npu_inst_int_data_y_1__4__0_), .A2(
        npu_inst_pe_1_0_4_n54), .B1(npu_inst_pe_1_0_4_n116), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_4_n53) );
  INV_X1 npu_inst_pe_1_0_4_U99 ( .A(npu_inst_pe_1_0_4_n53), .ZN(
        npu_inst_pe_1_0_4_n107) );
  AOI22_X1 npu_inst_pe_1_0_4_U98 ( .A1(npu_inst_int_data_y_1__4__0_), .A2(
        npu_inst_pe_1_0_4_n50), .B1(npu_inst_pe_1_0_4_n115), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_4_n49) );
  INV_X1 npu_inst_pe_1_0_4_U97 ( .A(npu_inst_pe_1_0_4_n49), .ZN(
        npu_inst_pe_1_0_4_n108) );
  AOI22_X1 npu_inst_pe_1_0_4_U96 ( .A1(npu_inst_int_data_y_1__4__0_), .A2(
        npu_inst_pe_1_0_4_n46), .B1(npu_inst_pe_1_0_4_n114), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_4_n45) );
  INV_X1 npu_inst_pe_1_0_4_U95 ( .A(npu_inst_pe_1_0_4_n45), .ZN(
        npu_inst_pe_1_0_4_n109) );
  AOI22_X1 npu_inst_pe_1_0_4_U94 ( .A1(npu_inst_int_data_y_1__4__0_), .A2(
        npu_inst_pe_1_0_4_n42), .B1(npu_inst_pe_1_0_4_n113), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_4_n41) );
  INV_X1 npu_inst_pe_1_0_4_U93 ( .A(npu_inst_pe_1_0_4_n41), .ZN(
        npu_inst_pe_1_0_4_n110) );
  AOI22_X1 npu_inst_pe_1_0_4_U92 ( .A1(npu_inst_int_data_y_1__4__1_), .A2(
        npu_inst_pe_1_0_4_n58), .B1(npu_inst_pe_1_0_4_n117), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_4_n59) );
  INV_X1 npu_inst_pe_1_0_4_U91 ( .A(npu_inst_pe_1_0_4_n59), .ZN(
        npu_inst_pe_1_0_4_n100) );
  AOI22_X1 npu_inst_pe_1_0_4_U90 ( .A1(npu_inst_int_data_y_1__4__1_), .A2(
        npu_inst_pe_1_0_4_n54), .B1(npu_inst_pe_1_0_4_n116), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_4_n55) );
  INV_X1 npu_inst_pe_1_0_4_U89 ( .A(npu_inst_pe_1_0_4_n55), .ZN(
        npu_inst_pe_1_0_4_n101) );
  AOI22_X1 npu_inst_pe_1_0_4_U88 ( .A1(npu_inst_int_data_y_1__4__1_), .A2(
        npu_inst_pe_1_0_4_n50), .B1(npu_inst_pe_1_0_4_n115), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_4_n51) );
  INV_X1 npu_inst_pe_1_0_4_U87 ( .A(npu_inst_pe_1_0_4_n51), .ZN(
        npu_inst_pe_1_0_4_n102) );
  AOI22_X1 npu_inst_pe_1_0_4_U86 ( .A1(npu_inst_int_data_y_1__4__1_), .A2(
        npu_inst_pe_1_0_4_n46), .B1(npu_inst_pe_1_0_4_n114), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_4_n47) );
  INV_X1 npu_inst_pe_1_0_4_U85 ( .A(npu_inst_pe_1_0_4_n47), .ZN(
        npu_inst_pe_1_0_4_n103) );
  AOI22_X1 npu_inst_pe_1_0_4_U84 ( .A1(npu_inst_int_data_y_1__4__1_), .A2(
        npu_inst_pe_1_0_4_n42), .B1(npu_inst_pe_1_0_4_n113), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_4_n43) );
  INV_X1 npu_inst_pe_1_0_4_U83 ( .A(npu_inst_pe_1_0_4_n43), .ZN(
        npu_inst_pe_1_0_4_n104) );
  AOI22_X1 npu_inst_pe_1_0_4_U82 ( .A1(npu_inst_pe_1_0_4_n38), .A2(
        npu_inst_int_data_y_1__4__1_), .B1(npu_inst_pe_1_0_4_n112), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_4_n39) );
  INV_X1 npu_inst_pe_1_0_4_U81 ( .A(npu_inst_pe_1_0_4_n39), .ZN(
        npu_inst_pe_1_0_4_n105) );
  NOR3_X1 npu_inst_pe_1_0_4_U80 ( .A1(npu_inst_pe_1_0_4_n26), .A2(npu_inst_n42), .A3(npu_inst_int_ckg[59]), .ZN(npu_inst_pe_1_0_4_n85) );
  OR2_X1 npu_inst_pe_1_0_4_U79 ( .A1(npu_inst_pe_1_0_4_n85), .A2(
        npu_inst_pe_1_0_4_n1), .ZN(npu_inst_pe_1_0_4_N84) );
  NAND2_X1 npu_inst_pe_1_0_4_U78 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_4_n60), .ZN(npu_inst_pe_1_0_4_n74) );
  OAI21_X1 npu_inst_pe_1_0_4_U77 ( .B1(npu_inst_pe_1_0_4_n63), .B2(
        npu_inst_pe_1_0_4_n60), .A(npu_inst_pe_1_0_4_n74), .ZN(
        npu_inst_pe_1_0_4_n97) );
  NAND2_X1 npu_inst_pe_1_0_4_U76 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_4_n60), .ZN(npu_inst_pe_1_0_4_n73) );
  OAI21_X1 npu_inst_pe_1_0_4_U75 ( .B1(npu_inst_pe_1_0_4_n61), .B2(
        npu_inst_pe_1_0_4_n60), .A(npu_inst_pe_1_0_4_n73), .ZN(
        npu_inst_pe_1_0_4_n96) );
  NAND2_X1 npu_inst_pe_1_0_4_U74 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_4_n56), .ZN(npu_inst_pe_1_0_4_n72) );
  OAI21_X1 npu_inst_pe_1_0_4_U73 ( .B1(npu_inst_pe_1_0_4_n63), .B2(
        npu_inst_pe_1_0_4_n56), .A(npu_inst_pe_1_0_4_n72), .ZN(
        npu_inst_pe_1_0_4_n95) );
  NAND2_X1 npu_inst_pe_1_0_4_U72 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_4_n56), .ZN(npu_inst_pe_1_0_4_n71) );
  OAI21_X1 npu_inst_pe_1_0_4_U71 ( .B1(npu_inst_pe_1_0_4_n61), .B2(
        npu_inst_pe_1_0_4_n56), .A(npu_inst_pe_1_0_4_n71), .ZN(
        npu_inst_pe_1_0_4_n94) );
  NAND2_X1 npu_inst_pe_1_0_4_U70 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_4_n52), .ZN(npu_inst_pe_1_0_4_n70) );
  OAI21_X1 npu_inst_pe_1_0_4_U69 ( .B1(npu_inst_pe_1_0_4_n63), .B2(
        npu_inst_pe_1_0_4_n52), .A(npu_inst_pe_1_0_4_n70), .ZN(
        npu_inst_pe_1_0_4_n93) );
  NAND2_X1 npu_inst_pe_1_0_4_U68 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_4_n52), .ZN(npu_inst_pe_1_0_4_n69) );
  OAI21_X1 npu_inst_pe_1_0_4_U67 ( .B1(npu_inst_pe_1_0_4_n61), .B2(
        npu_inst_pe_1_0_4_n52), .A(npu_inst_pe_1_0_4_n69), .ZN(
        npu_inst_pe_1_0_4_n92) );
  NAND2_X1 npu_inst_pe_1_0_4_U66 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_4_n48), .ZN(npu_inst_pe_1_0_4_n68) );
  OAI21_X1 npu_inst_pe_1_0_4_U65 ( .B1(npu_inst_pe_1_0_4_n63), .B2(
        npu_inst_pe_1_0_4_n48), .A(npu_inst_pe_1_0_4_n68), .ZN(
        npu_inst_pe_1_0_4_n91) );
  NAND2_X1 npu_inst_pe_1_0_4_U64 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_4_n48), .ZN(npu_inst_pe_1_0_4_n67) );
  OAI21_X1 npu_inst_pe_1_0_4_U63 ( .B1(npu_inst_pe_1_0_4_n61), .B2(
        npu_inst_pe_1_0_4_n48), .A(npu_inst_pe_1_0_4_n67), .ZN(
        npu_inst_pe_1_0_4_n90) );
  NAND2_X1 npu_inst_pe_1_0_4_U62 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_4_n44), .ZN(npu_inst_pe_1_0_4_n66) );
  OAI21_X1 npu_inst_pe_1_0_4_U61 ( .B1(npu_inst_pe_1_0_4_n63), .B2(
        npu_inst_pe_1_0_4_n44), .A(npu_inst_pe_1_0_4_n66), .ZN(
        npu_inst_pe_1_0_4_n89) );
  NAND2_X1 npu_inst_pe_1_0_4_U60 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_4_n44), .ZN(npu_inst_pe_1_0_4_n65) );
  OAI21_X1 npu_inst_pe_1_0_4_U59 ( .B1(npu_inst_pe_1_0_4_n61), .B2(
        npu_inst_pe_1_0_4_n44), .A(npu_inst_pe_1_0_4_n65), .ZN(
        npu_inst_pe_1_0_4_n88) );
  NAND2_X1 npu_inst_pe_1_0_4_U58 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_4_n40), .ZN(npu_inst_pe_1_0_4_n64) );
  OAI21_X1 npu_inst_pe_1_0_4_U57 ( .B1(npu_inst_pe_1_0_4_n63), .B2(
        npu_inst_pe_1_0_4_n40), .A(npu_inst_pe_1_0_4_n64), .ZN(
        npu_inst_pe_1_0_4_n87) );
  NAND2_X1 npu_inst_pe_1_0_4_U56 ( .A1(npu_inst_pe_1_0_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_4_n40), .ZN(npu_inst_pe_1_0_4_n62) );
  OAI21_X1 npu_inst_pe_1_0_4_U55 ( .B1(npu_inst_pe_1_0_4_n61), .B2(
        npu_inst_pe_1_0_4_n40), .A(npu_inst_pe_1_0_4_n62), .ZN(
        npu_inst_pe_1_0_4_n86) );
  AOI22_X1 npu_inst_pe_1_0_4_U54 ( .A1(npu_inst_pe_1_0_4_n38), .A2(
        npu_inst_int_data_y_1__4__0_), .B1(npu_inst_pe_1_0_4_n112), .B2(
        npu_inst_pe_1_0_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_4_n37) );
  INV_X1 npu_inst_pe_1_0_4_U53 ( .A(npu_inst_pe_1_0_4_n37), .ZN(
        npu_inst_pe_1_0_4_n111) );
  AOI222_X1 npu_inst_pe_1_0_4_U52 ( .A1(npu_inst_int_data_res_1__4__0_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N73), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N65), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n84) );
  INV_X1 npu_inst_pe_1_0_4_U51 ( .A(npu_inst_pe_1_0_4_n84), .ZN(
        npu_inst_pe_1_0_4_n99) );
  AOI222_X1 npu_inst_pe_1_0_4_U50 ( .A1(npu_inst_pe_1_0_4_n1), .A2(
        npu_inst_int_data_res_1__4__7_), .B1(npu_inst_pe_1_0_4_N80), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N72), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n75) );
  INV_X1 npu_inst_pe_1_0_4_U49 ( .A(npu_inst_pe_1_0_4_n75), .ZN(
        npu_inst_pe_1_0_4_n31) );
  AOI222_X1 npu_inst_pe_1_0_4_U48 ( .A1(npu_inst_int_data_res_1__4__2_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N75), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N67), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n82) );
  INV_X1 npu_inst_pe_1_0_4_U47 ( .A(npu_inst_pe_1_0_4_n82), .ZN(
        npu_inst_pe_1_0_4_n36) );
  AOI222_X1 npu_inst_pe_1_0_4_U46 ( .A1(npu_inst_int_data_res_1__4__3_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N76), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N68), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n81) );
  INV_X1 npu_inst_pe_1_0_4_U45 ( .A(npu_inst_pe_1_0_4_n81), .ZN(
        npu_inst_pe_1_0_4_n35) );
  AOI222_X1 npu_inst_pe_1_0_4_U44 ( .A1(npu_inst_int_data_res_1__4__4_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N77), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N69), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n80) );
  INV_X1 npu_inst_pe_1_0_4_U43 ( .A(npu_inst_pe_1_0_4_n80), .ZN(
        npu_inst_pe_1_0_4_n34) );
  AOI222_X1 npu_inst_pe_1_0_4_U42 ( .A1(npu_inst_int_data_res_1__4__5_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N78), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N70), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n79) );
  INV_X1 npu_inst_pe_1_0_4_U41 ( .A(npu_inst_pe_1_0_4_n79), .ZN(
        npu_inst_pe_1_0_4_n33) );
  AOI222_X1 npu_inst_pe_1_0_4_U40 ( .A1(npu_inst_int_data_res_1__4__6_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N79), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N71), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n78) );
  INV_X1 npu_inst_pe_1_0_4_U39 ( .A(npu_inst_pe_1_0_4_n78), .ZN(
        npu_inst_pe_1_0_4_n32) );
  AND2_X1 npu_inst_pe_1_0_4_U38 ( .A1(npu_inst_int_data_x_0__4__1_), .A2(
        npu_inst_pe_1_0_4_int_q_weight_1_), .ZN(npu_inst_pe_1_0_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_4_U37 ( .A1(npu_inst_int_data_x_0__4__0_), .A2(
        npu_inst_pe_1_0_4_int_q_weight_1_), .ZN(npu_inst_pe_1_0_4_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_0_4_U36 ( .A(npu_inst_pe_1_0_4_int_data_1_), .ZN(
        npu_inst_pe_1_0_4_n12) );
  AOI222_X1 npu_inst_pe_1_0_4_U35 ( .A1(npu_inst_int_data_res_1__4__1_), .A2(
        npu_inst_pe_1_0_4_n1), .B1(npu_inst_pe_1_0_4_N74), .B2(
        npu_inst_pe_1_0_4_n76), .C1(npu_inst_pe_1_0_4_N66), .C2(
        npu_inst_pe_1_0_4_n77), .ZN(npu_inst_pe_1_0_4_n83) );
  INV_X1 npu_inst_pe_1_0_4_U34 ( .A(npu_inst_pe_1_0_4_n83), .ZN(
        npu_inst_pe_1_0_4_n98) );
  AND2_X1 npu_inst_pe_1_0_4_U33 ( .A1(npu_inst_pe_1_0_4_N93), .A2(npu_inst_n42), .ZN(npu_inst_pe_1_0_4_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_4_U32 ( .A1(npu_inst_n42), .A2(npu_inst_pe_1_0_4_N94), .ZN(npu_inst_pe_1_0_4_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_4_U31 ( .A1(npu_inst_n42), .A2(
        npu_inst_int_data_y_1__4__1_), .B1(npu_inst_pe_1_0_4_n2), .B2(
        npu_inst_int_data_x_0__5__1_), .ZN(npu_inst_pe_1_0_4_n63) );
  AOI22_X1 npu_inst_pe_1_0_4_U30 ( .A1(npu_inst_n42), .A2(
        npu_inst_int_data_y_1__4__0_), .B1(npu_inst_pe_1_0_4_n2), .B2(
        npu_inst_int_data_x_0__5__0_), .ZN(npu_inst_pe_1_0_4_n61) );
  INV_X1 npu_inst_pe_1_0_4_U29 ( .A(npu_inst_pe_1_0_4_int_data_0_), .ZN(
        npu_inst_pe_1_0_4_n11) );
  INV_X1 npu_inst_pe_1_0_4_U28 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_0_4_n4)
         );
  OR3_X1 npu_inst_pe_1_0_4_U27 ( .A1(npu_inst_n61), .A2(npu_inst_pe_1_0_4_n6), 
        .A3(npu_inst_pe_1_0_4_n4), .ZN(npu_inst_pe_1_0_4_n56) );
  OR3_X1 npu_inst_pe_1_0_4_U26 ( .A1(npu_inst_pe_1_0_4_n4), .A2(
        npu_inst_pe_1_0_4_n6), .A3(npu_inst_pe_1_0_4_n5), .ZN(
        npu_inst_pe_1_0_4_n48) );
  INV_X1 npu_inst_pe_1_0_4_U25 ( .A(npu_inst_pe_1_0_4_n4), .ZN(
        npu_inst_pe_1_0_4_n3) );
  OR3_X1 npu_inst_pe_1_0_4_U24 ( .A1(npu_inst_pe_1_0_4_n3), .A2(
        npu_inst_pe_1_0_4_n6), .A3(npu_inst_pe_1_0_4_n5), .ZN(
        npu_inst_pe_1_0_4_n52) );
  OR3_X1 npu_inst_pe_1_0_4_U23 ( .A1(npu_inst_n61), .A2(npu_inst_pe_1_0_4_n6), 
        .A3(npu_inst_pe_1_0_4_n3), .ZN(npu_inst_pe_1_0_4_n60) );
  BUF_X1 npu_inst_pe_1_0_4_U22 ( .A(npu_inst_n30), .Z(npu_inst_pe_1_0_4_n1) );
  NOR2_X1 npu_inst_pe_1_0_4_U21 ( .A1(npu_inst_pe_1_0_4_n60), .A2(
        npu_inst_pe_1_0_4_n2), .ZN(npu_inst_pe_1_0_4_n58) );
  NOR2_X1 npu_inst_pe_1_0_4_U20 ( .A1(npu_inst_pe_1_0_4_n56), .A2(
        npu_inst_pe_1_0_4_n2), .ZN(npu_inst_pe_1_0_4_n54) );
  NOR2_X1 npu_inst_pe_1_0_4_U19 ( .A1(npu_inst_pe_1_0_4_n52), .A2(
        npu_inst_pe_1_0_4_n2), .ZN(npu_inst_pe_1_0_4_n50) );
  NOR2_X1 npu_inst_pe_1_0_4_U18 ( .A1(npu_inst_pe_1_0_4_n48), .A2(
        npu_inst_pe_1_0_4_n2), .ZN(npu_inst_pe_1_0_4_n46) );
  NOR2_X1 npu_inst_pe_1_0_4_U17 ( .A1(npu_inst_pe_1_0_4_n40), .A2(
        npu_inst_pe_1_0_4_n2), .ZN(npu_inst_pe_1_0_4_n38) );
  NOR2_X1 npu_inst_pe_1_0_4_U16 ( .A1(npu_inst_pe_1_0_4_n44), .A2(
        npu_inst_pe_1_0_4_n2), .ZN(npu_inst_pe_1_0_4_n42) );
  BUF_X1 npu_inst_pe_1_0_4_U15 ( .A(npu_inst_n88), .Z(npu_inst_pe_1_0_4_n6) );
  INV_X1 npu_inst_pe_1_0_4_U14 ( .A(npu_inst_n108), .ZN(npu_inst_pe_1_0_4_n10)
         );
  INV_X1 npu_inst_pe_1_0_4_U13 ( .A(npu_inst_pe_1_0_4_n38), .ZN(
        npu_inst_pe_1_0_4_n112) );
  INV_X1 npu_inst_pe_1_0_4_U12 ( .A(npu_inst_pe_1_0_4_n58), .ZN(
        npu_inst_pe_1_0_4_n117) );
  INV_X1 npu_inst_pe_1_0_4_U11 ( .A(npu_inst_pe_1_0_4_n54), .ZN(
        npu_inst_pe_1_0_4_n116) );
  INV_X1 npu_inst_pe_1_0_4_U10 ( .A(npu_inst_pe_1_0_4_n50), .ZN(
        npu_inst_pe_1_0_4_n115) );
  INV_X1 npu_inst_pe_1_0_4_U9 ( .A(npu_inst_pe_1_0_4_n46), .ZN(
        npu_inst_pe_1_0_4_n114) );
  INV_X1 npu_inst_pe_1_0_4_U8 ( .A(npu_inst_pe_1_0_4_n42), .ZN(
        npu_inst_pe_1_0_4_n113) );
  BUF_X1 npu_inst_pe_1_0_4_U7 ( .A(npu_inst_pe_1_0_4_n10), .Z(
        npu_inst_pe_1_0_4_n9) );
  BUF_X1 npu_inst_pe_1_0_4_U6 ( .A(npu_inst_pe_1_0_4_n10), .Z(
        npu_inst_pe_1_0_4_n8) );
  BUF_X1 npu_inst_pe_1_0_4_U5 ( .A(npu_inst_pe_1_0_4_n10), .Z(
        npu_inst_pe_1_0_4_n7) );
  NOR2_X1 npu_inst_pe_1_0_4_U4 ( .A1(npu_inst_pe_1_0_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_4_n1), .ZN(npu_inst_pe_1_0_4_n76) );
  NOR2_X1 npu_inst_pe_1_0_4_U3 ( .A1(npu_inst_pe_1_0_4_n27), .A2(
        npu_inst_pe_1_0_4_n1), .ZN(npu_inst_pe_1_0_4_n77) );
  FA_X1 npu_inst_pe_1_0_4_sub_77_U2_1 ( .A(int_o_data_npu[25]), .B(
        npu_inst_pe_1_0_4_n12), .CI(npu_inst_pe_1_0_4_sub_77_carry_1_), .CO(
        npu_inst_pe_1_0_4_sub_77_carry_2_), .S(npu_inst_pe_1_0_4_N66) );
  FA_X1 npu_inst_pe_1_0_4_add_79_U1_1 ( .A(int_o_data_npu[25]), .B(
        npu_inst_pe_1_0_4_int_data_1_), .CI(npu_inst_pe_1_0_4_add_79_carry_1_), 
        .CO(npu_inst_pe_1_0_4_add_79_carry_2_), .S(npu_inst_pe_1_0_4_N74) );
  NAND3_X1 npu_inst_pe_1_0_4_U101 ( .A1(npu_inst_pe_1_0_4_n4), .A2(
        npu_inst_pe_1_0_4_n5), .A3(npu_inst_pe_1_0_4_n6), .ZN(
        npu_inst_pe_1_0_4_n44) );
  NAND3_X1 npu_inst_pe_1_0_4_U100 ( .A1(npu_inst_pe_1_0_4_n3), .A2(
        npu_inst_pe_1_0_4_n5), .A3(npu_inst_pe_1_0_4_n6), .ZN(
        npu_inst_pe_1_0_4_n40) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_4_n32), .CK(
        npu_inst_pe_1_0_4_net4386), .RN(npu_inst_pe_1_0_4_n7), .Q(
        int_o_data_npu[30]) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_4_n33), .CK(
        npu_inst_pe_1_0_4_net4386), .RN(npu_inst_pe_1_0_4_n7), .Q(
        int_o_data_npu[29]) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_4_n34), .CK(
        npu_inst_pe_1_0_4_net4386), .RN(npu_inst_pe_1_0_4_n7), .Q(
        int_o_data_npu[28]) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_4_n35), .CK(
        npu_inst_pe_1_0_4_net4386), .RN(npu_inst_pe_1_0_4_n7), .Q(
        int_o_data_npu[27]) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_4_n36), .CK(
        npu_inst_pe_1_0_4_net4386), .RN(npu_inst_pe_1_0_4_n7), .Q(
        int_o_data_npu[26]) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_4_n98), .CK(
        npu_inst_pe_1_0_4_net4386), .RN(npu_inst_pe_1_0_4_n7), .Q(
        int_o_data_npu[25]) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_4_n31), .CK(
        npu_inst_pe_1_0_4_net4386), .RN(npu_inst_pe_1_0_4_n7), .Q(
        int_o_data_npu[31]) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_4_n99), .CK(
        npu_inst_pe_1_0_4_net4386), .RN(npu_inst_pe_1_0_4_n7), .Q(
        int_o_data_npu[24]) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_weight_reg_0_ ( .D(npu_inst_n94), .CK(
        npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n7), .Q(
        npu_inst_pe_1_0_4_int_q_weight_0_), .QN(npu_inst_pe_1_0_4_n27) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_weight_reg_1_ ( .D(npu_inst_n100), .CK(
        npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n7), .Q(
        npu_inst_pe_1_0_4_int_q_weight_1_), .QN(npu_inst_pe_1_0_4_n26) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_4_n111), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n7), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_4_n105), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n7), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_4_n110), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_4_n104), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_4_n109), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_4_n103), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_4_n108), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_4_n102), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_4_n107), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_4_n101), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_4_n106), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_4_n100), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_4_n86), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_4_n87), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n8), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_4_n88), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_4_n89), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_4_n90), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_4_n91), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_4_n92), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_4_n93), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_4_n94), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_4_n95), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_4_n96), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_4_n97), 
        .CK(npu_inst_pe_1_0_4_net4392), .RN(npu_inst_pe_1_0_4_n9), .Q(
        npu_inst_pe_1_0_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_4_net4386) );
  CLKGATETST_X1 npu_inst_pe_1_0_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n48), .SE(1'b0), .GCK(npu_inst_pe_1_0_4_net4392) );
  MUX2_X1 npu_inst_pe_1_0_5_U153 ( .A(npu_inst_pe_1_0_5_n31), .B(
        npu_inst_pe_1_0_5_n28), .S(npu_inst_pe_1_0_5_n7), .Z(
        npu_inst_pe_1_0_5_N93) );
  MUX2_X1 npu_inst_pe_1_0_5_U152 ( .A(npu_inst_pe_1_0_5_n30), .B(
        npu_inst_pe_1_0_5_n29), .S(npu_inst_pe_1_0_5_n5), .Z(
        npu_inst_pe_1_0_5_n31) );
  MUX2_X1 npu_inst_pe_1_0_5_U151 ( .A(npu_inst_pe_1_0_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_5_n3), .Z(
        npu_inst_pe_1_0_5_n30) );
  MUX2_X1 npu_inst_pe_1_0_5_U150 ( .A(npu_inst_pe_1_0_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_5_n3), .Z(
        npu_inst_pe_1_0_5_n29) );
  MUX2_X1 npu_inst_pe_1_0_5_U149 ( .A(npu_inst_pe_1_0_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_5_n3), .Z(
        npu_inst_pe_1_0_5_n28) );
  MUX2_X1 npu_inst_pe_1_0_5_U148 ( .A(npu_inst_pe_1_0_5_n25), .B(
        npu_inst_pe_1_0_5_n22), .S(npu_inst_pe_1_0_5_n7), .Z(
        npu_inst_pe_1_0_5_N94) );
  MUX2_X1 npu_inst_pe_1_0_5_U147 ( .A(npu_inst_pe_1_0_5_n24), .B(
        npu_inst_pe_1_0_5_n23), .S(npu_inst_pe_1_0_5_n5), .Z(
        npu_inst_pe_1_0_5_n25) );
  MUX2_X1 npu_inst_pe_1_0_5_U146 ( .A(npu_inst_pe_1_0_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_5_n3), .Z(
        npu_inst_pe_1_0_5_n24) );
  MUX2_X1 npu_inst_pe_1_0_5_U145 ( .A(npu_inst_pe_1_0_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_5_n3), .Z(
        npu_inst_pe_1_0_5_n23) );
  MUX2_X1 npu_inst_pe_1_0_5_U144 ( .A(npu_inst_pe_1_0_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_5_n3), .Z(
        npu_inst_pe_1_0_5_n22) );
  MUX2_X1 npu_inst_pe_1_0_5_U143 ( .A(npu_inst_pe_1_0_5_n21), .B(
        npu_inst_pe_1_0_5_n18), .S(npu_inst_pe_1_0_5_n7), .Z(
        npu_inst_int_data_x_0__5__1_) );
  MUX2_X1 npu_inst_pe_1_0_5_U142 ( .A(npu_inst_pe_1_0_5_n20), .B(
        npu_inst_pe_1_0_5_n19), .S(npu_inst_pe_1_0_5_n5), .Z(
        npu_inst_pe_1_0_5_n21) );
  MUX2_X1 npu_inst_pe_1_0_5_U141 ( .A(npu_inst_pe_1_0_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_5_n3), .Z(
        npu_inst_pe_1_0_5_n20) );
  MUX2_X1 npu_inst_pe_1_0_5_U140 ( .A(npu_inst_pe_1_0_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_5_n3), .Z(
        npu_inst_pe_1_0_5_n19) );
  MUX2_X1 npu_inst_pe_1_0_5_U139 ( .A(npu_inst_pe_1_0_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_5_n3), .Z(
        npu_inst_pe_1_0_5_n18) );
  MUX2_X1 npu_inst_pe_1_0_5_U138 ( .A(npu_inst_pe_1_0_5_n17), .B(
        npu_inst_pe_1_0_5_n14), .S(npu_inst_pe_1_0_5_n7), .Z(
        npu_inst_int_data_x_0__5__0_) );
  MUX2_X1 npu_inst_pe_1_0_5_U137 ( .A(npu_inst_pe_1_0_5_n16), .B(
        npu_inst_pe_1_0_5_n15), .S(npu_inst_pe_1_0_5_n5), .Z(
        npu_inst_pe_1_0_5_n17) );
  MUX2_X1 npu_inst_pe_1_0_5_U136 ( .A(npu_inst_pe_1_0_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_5_n3), .Z(
        npu_inst_pe_1_0_5_n16) );
  MUX2_X1 npu_inst_pe_1_0_5_U135 ( .A(npu_inst_pe_1_0_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_5_n3), .Z(
        npu_inst_pe_1_0_5_n15) );
  MUX2_X1 npu_inst_pe_1_0_5_U134 ( .A(npu_inst_pe_1_0_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_5_n3), .Z(
        npu_inst_pe_1_0_5_n14) );
  XOR2_X1 npu_inst_pe_1_0_5_U133 ( .A(npu_inst_pe_1_0_5_int_data_0_), .B(
        int_o_data_npu[16]), .Z(npu_inst_pe_1_0_5_N73) );
  AND2_X1 npu_inst_pe_1_0_5_U132 ( .A1(int_o_data_npu[16]), .A2(
        npu_inst_pe_1_0_5_int_data_0_), .ZN(npu_inst_pe_1_0_5_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_5_U131 ( .A(int_o_data_npu[16]), .B(
        npu_inst_pe_1_0_5_n12), .ZN(npu_inst_pe_1_0_5_N65) );
  OR2_X1 npu_inst_pe_1_0_5_U130 ( .A1(npu_inst_pe_1_0_5_n12), .A2(
        int_o_data_npu[16]), .ZN(npu_inst_pe_1_0_5_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_5_U129 ( .A(int_o_data_npu[18]), .B(
        npu_inst_pe_1_0_5_add_79_carry_2_), .Z(npu_inst_pe_1_0_5_N75) );
  AND2_X1 npu_inst_pe_1_0_5_U128 ( .A1(npu_inst_pe_1_0_5_add_79_carry_2_), 
        .A2(int_o_data_npu[18]), .ZN(npu_inst_pe_1_0_5_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_5_U127 ( .A(int_o_data_npu[19]), .B(
        npu_inst_pe_1_0_5_add_79_carry_3_), .Z(npu_inst_pe_1_0_5_N76) );
  AND2_X1 npu_inst_pe_1_0_5_U126 ( .A1(npu_inst_pe_1_0_5_add_79_carry_3_), 
        .A2(int_o_data_npu[19]), .ZN(npu_inst_pe_1_0_5_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_5_U125 ( .A(int_o_data_npu[20]), .B(
        npu_inst_pe_1_0_5_add_79_carry_4_), .Z(npu_inst_pe_1_0_5_N77) );
  AND2_X1 npu_inst_pe_1_0_5_U124 ( .A1(npu_inst_pe_1_0_5_add_79_carry_4_), 
        .A2(int_o_data_npu[20]), .ZN(npu_inst_pe_1_0_5_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_5_U123 ( .A(int_o_data_npu[21]), .B(
        npu_inst_pe_1_0_5_add_79_carry_5_), .Z(npu_inst_pe_1_0_5_N78) );
  AND2_X1 npu_inst_pe_1_0_5_U122 ( .A1(npu_inst_pe_1_0_5_add_79_carry_5_), 
        .A2(int_o_data_npu[21]), .ZN(npu_inst_pe_1_0_5_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_5_U121 ( .A(int_o_data_npu[22]), .B(
        npu_inst_pe_1_0_5_add_79_carry_6_), .Z(npu_inst_pe_1_0_5_N79) );
  AND2_X1 npu_inst_pe_1_0_5_U120 ( .A1(npu_inst_pe_1_0_5_add_79_carry_6_), 
        .A2(int_o_data_npu[22]), .ZN(npu_inst_pe_1_0_5_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_5_U119 ( .A(int_o_data_npu[23]), .B(
        npu_inst_pe_1_0_5_add_79_carry_7_), .Z(npu_inst_pe_1_0_5_N80) );
  XNOR2_X1 npu_inst_pe_1_0_5_U118 ( .A(npu_inst_pe_1_0_5_sub_77_carry_2_), .B(
        int_o_data_npu[18]), .ZN(npu_inst_pe_1_0_5_N67) );
  OR2_X1 npu_inst_pe_1_0_5_U117 ( .A1(int_o_data_npu[18]), .A2(
        npu_inst_pe_1_0_5_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_0_5_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_5_U116 ( .A(npu_inst_pe_1_0_5_sub_77_carry_3_), .B(
        int_o_data_npu[19]), .ZN(npu_inst_pe_1_0_5_N68) );
  OR2_X1 npu_inst_pe_1_0_5_U115 ( .A1(int_o_data_npu[19]), .A2(
        npu_inst_pe_1_0_5_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_0_5_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_5_U114 ( .A(npu_inst_pe_1_0_5_sub_77_carry_4_), .B(
        int_o_data_npu[20]), .ZN(npu_inst_pe_1_0_5_N69) );
  OR2_X1 npu_inst_pe_1_0_5_U113 ( .A1(int_o_data_npu[20]), .A2(
        npu_inst_pe_1_0_5_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_0_5_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_5_U112 ( .A(npu_inst_pe_1_0_5_sub_77_carry_5_), .B(
        int_o_data_npu[21]), .ZN(npu_inst_pe_1_0_5_N70) );
  OR2_X1 npu_inst_pe_1_0_5_U111 ( .A1(int_o_data_npu[21]), .A2(
        npu_inst_pe_1_0_5_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_0_5_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_5_U110 ( .A(npu_inst_pe_1_0_5_sub_77_carry_6_), .B(
        int_o_data_npu[22]), .ZN(npu_inst_pe_1_0_5_N71) );
  OR2_X1 npu_inst_pe_1_0_5_U109 ( .A1(int_o_data_npu[22]), .A2(
        npu_inst_pe_1_0_5_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_0_5_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_5_U108 ( .A(int_o_data_npu[23]), .B(
        npu_inst_pe_1_0_5_sub_77_carry_7_), .ZN(npu_inst_pe_1_0_5_N72) );
  INV_X1 npu_inst_pe_1_0_5_U107 ( .A(npu_inst_n61), .ZN(npu_inst_pe_1_0_5_n6)
         );
  INV_X1 npu_inst_pe_1_0_5_U106 ( .A(npu_inst_pe_1_0_5_n6), .ZN(
        npu_inst_pe_1_0_5_n5) );
  INV_X1 npu_inst_pe_1_0_5_U105 ( .A(npu_inst_n42), .ZN(npu_inst_pe_1_0_5_n2)
         );
  AOI22_X1 npu_inst_pe_1_0_5_U104 ( .A1(npu_inst_int_data_y_1__5__0_), .A2(
        npu_inst_pe_1_0_5_n58), .B1(npu_inst_pe_1_0_5_n118), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_5_n57) );
  INV_X1 npu_inst_pe_1_0_5_U103 ( .A(npu_inst_pe_1_0_5_n57), .ZN(
        npu_inst_pe_1_0_5_n107) );
  AOI22_X1 npu_inst_pe_1_0_5_U102 ( .A1(npu_inst_int_data_y_1__5__0_), .A2(
        npu_inst_pe_1_0_5_n54), .B1(npu_inst_pe_1_0_5_n117), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_5_n53) );
  INV_X1 npu_inst_pe_1_0_5_U99 ( .A(npu_inst_pe_1_0_5_n53), .ZN(
        npu_inst_pe_1_0_5_n108) );
  AOI22_X1 npu_inst_pe_1_0_5_U98 ( .A1(npu_inst_int_data_y_1__5__0_), .A2(
        npu_inst_pe_1_0_5_n50), .B1(npu_inst_pe_1_0_5_n116), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_5_n49) );
  INV_X1 npu_inst_pe_1_0_5_U97 ( .A(npu_inst_pe_1_0_5_n49), .ZN(
        npu_inst_pe_1_0_5_n109) );
  AOI22_X1 npu_inst_pe_1_0_5_U96 ( .A1(npu_inst_int_data_y_1__5__0_), .A2(
        npu_inst_pe_1_0_5_n46), .B1(npu_inst_pe_1_0_5_n115), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_5_n45) );
  INV_X1 npu_inst_pe_1_0_5_U95 ( .A(npu_inst_pe_1_0_5_n45), .ZN(
        npu_inst_pe_1_0_5_n110) );
  AOI22_X1 npu_inst_pe_1_0_5_U94 ( .A1(npu_inst_int_data_y_1__5__0_), .A2(
        npu_inst_pe_1_0_5_n42), .B1(npu_inst_pe_1_0_5_n114), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_5_n41) );
  INV_X1 npu_inst_pe_1_0_5_U93 ( .A(npu_inst_pe_1_0_5_n41), .ZN(
        npu_inst_pe_1_0_5_n111) );
  AOI22_X1 npu_inst_pe_1_0_5_U92 ( .A1(npu_inst_int_data_y_1__5__1_), .A2(
        npu_inst_pe_1_0_5_n58), .B1(npu_inst_pe_1_0_5_n118), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_5_n59) );
  INV_X1 npu_inst_pe_1_0_5_U91 ( .A(npu_inst_pe_1_0_5_n59), .ZN(
        npu_inst_pe_1_0_5_n101) );
  AOI22_X1 npu_inst_pe_1_0_5_U90 ( .A1(npu_inst_int_data_y_1__5__1_), .A2(
        npu_inst_pe_1_0_5_n54), .B1(npu_inst_pe_1_0_5_n117), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_5_n55) );
  INV_X1 npu_inst_pe_1_0_5_U89 ( .A(npu_inst_pe_1_0_5_n55), .ZN(
        npu_inst_pe_1_0_5_n102) );
  AOI22_X1 npu_inst_pe_1_0_5_U88 ( .A1(npu_inst_int_data_y_1__5__1_), .A2(
        npu_inst_pe_1_0_5_n50), .B1(npu_inst_pe_1_0_5_n116), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_5_n51) );
  INV_X1 npu_inst_pe_1_0_5_U87 ( .A(npu_inst_pe_1_0_5_n51), .ZN(
        npu_inst_pe_1_0_5_n103) );
  AOI22_X1 npu_inst_pe_1_0_5_U86 ( .A1(npu_inst_int_data_y_1__5__1_), .A2(
        npu_inst_pe_1_0_5_n46), .B1(npu_inst_pe_1_0_5_n115), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_5_n47) );
  INV_X1 npu_inst_pe_1_0_5_U85 ( .A(npu_inst_pe_1_0_5_n47), .ZN(
        npu_inst_pe_1_0_5_n104) );
  AOI22_X1 npu_inst_pe_1_0_5_U84 ( .A1(npu_inst_int_data_y_1__5__1_), .A2(
        npu_inst_pe_1_0_5_n42), .B1(npu_inst_pe_1_0_5_n114), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_5_n43) );
  INV_X1 npu_inst_pe_1_0_5_U83 ( .A(npu_inst_pe_1_0_5_n43), .ZN(
        npu_inst_pe_1_0_5_n105) );
  AOI22_X1 npu_inst_pe_1_0_5_U82 ( .A1(npu_inst_pe_1_0_5_n38), .A2(
        npu_inst_int_data_y_1__5__1_), .B1(npu_inst_pe_1_0_5_n113), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_5_n39) );
  INV_X1 npu_inst_pe_1_0_5_U81 ( .A(npu_inst_pe_1_0_5_n39), .ZN(
        npu_inst_pe_1_0_5_n106) );
  NAND2_X1 npu_inst_pe_1_0_5_U80 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_5_n60), .ZN(npu_inst_pe_1_0_5_n74) );
  OAI21_X1 npu_inst_pe_1_0_5_U79 ( .B1(npu_inst_pe_1_0_5_n63), .B2(
        npu_inst_pe_1_0_5_n60), .A(npu_inst_pe_1_0_5_n74), .ZN(
        npu_inst_pe_1_0_5_n97) );
  NAND2_X1 npu_inst_pe_1_0_5_U78 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_5_n60), .ZN(npu_inst_pe_1_0_5_n73) );
  OAI21_X1 npu_inst_pe_1_0_5_U77 ( .B1(npu_inst_pe_1_0_5_n61), .B2(
        npu_inst_pe_1_0_5_n60), .A(npu_inst_pe_1_0_5_n73), .ZN(
        npu_inst_pe_1_0_5_n96) );
  NAND2_X1 npu_inst_pe_1_0_5_U76 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_5_n56), .ZN(npu_inst_pe_1_0_5_n72) );
  OAI21_X1 npu_inst_pe_1_0_5_U75 ( .B1(npu_inst_pe_1_0_5_n63), .B2(
        npu_inst_pe_1_0_5_n56), .A(npu_inst_pe_1_0_5_n72), .ZN(
        npu_inst_pe_1_0_5_n95) );
  NAND2_X1 npu_inst_pe_1_0_5_U74 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_5_n56), .ZN(npu_inst_pe_1_0_5_n71) );
  OAI21_X1 npu_inst_pe_1_0_5_U73 ( .B1(npu_inst_pe_1_0_5_n61), .B2(
        npu_inst_pe_1_0_5_n56), .A(npu_inst_pe_1_0_5_n71), .ZN(
        npu_inst_pe_1_0_5_n94) );
  NAND2_X1 npu_inst_pe_1_0_5_U72 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_5_n52), .ZN(npu_inst_pe_1_0_5_n70) );
  OAI21_X1 npu_inst_pe_1_0_5_U71 ( .B1(npu_inst_pe_1_0_5_n63), .B2(
        npu_inst_pe_1_0_5_n52), .A(npu_inst_pe_1_0_5_n70), .ZN(
        npu_inst_pe_1_0_5_n93) );
  NAND2_X1 npu_inst_pe_1_0_5_U70 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_5_n52), .ZN(npu_inst_pe_1_0_5_n69) );
  OAI21_X1 npu_inst_pe_1_0_5_U69 ( .B1(npu_inst_pe_1_0_5_n61), .B2(
        npu_inst_pe_1_0_5_n52), .A(npu_inst_pe_1_0_5_n69), .ZN(
        npu_inst_pe_1_0_5_n92) );
  NAND2_X1 npu_inst_pe_1_0_5_U68 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_5_n48), .ZN(npu_inst_pe_1_0_5_n68) );
  OAI21_X1 npu_inst_pe_1_0_5_U67 ( .B1(npu_inst_pe_1_0_5_n63), .B2(
        npu_inst_pe_1_0_5_n48), .A(npu_inst_pe_1_0_5_n68), .ZN(
        npu_inst_pe_1_0_5_n91) );
  NAND2_X1 npu_inst_pe_1_0_5_U66 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_5_n48), .ZN(npu_inst_pe_1_0_5_n67) );
  OAI21_X1 npu_inst_pe_1_0_5_U65 ( .B1(npu_inst_pe_1_0_5_n61), .B2(
        npu_inst_pe_1_0_5_n48), .A(npu_inst_pe_1_0_5_n67), .ZN(
        npu_inst_pe_1_0_5_n90) );
  NAND2_X1 npu_inst_pe_1_0_5_U64 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_5_n44), .ZN(npu_inst_pe_1_0_5_n66) );
  OAI21_X1 npu_inst_pe_1_0_5_U63 ( .B1(npu_inst_pe_1_0_5_n63), .B2(
        npu_inst_pe_1_0_5_n44), .A(npu_inst_pe_1_0_5_n66), .ZN(
        npu_inst_pe_1_0_5_n89) );
  NAND2_X1 npu_inst_pe_1_0_5_U62 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_5_n44), .ZN(npu_inst_pe_1_0_5_n65) );
  OAI21_X1 npu_inst_pe_1_0_5_U61 ( .B1(npu_inst_pe_1_0_5_n61), .B2(
        npu_inst_pe_1_0_5_n44), .A(npu_inst_pe_1_0_5_n65), .ZN(
        npu_inst_pe_1_0_5_n88) );
  NAND2_X1 npu_inst_pe_1_0_5_U60 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_5_n40), .ZN(npu_inst_pe_1_0_5_n64) );
  OAI21_X1 npu_inst_pe_1_0_5_U59 ( .B1(npu_inst_pe_1_0_5_n63), .B2(
        npu_inst_pe_1_0_5_n40), .A(npu_inst_pe_1_0_5_n64), .ZN(
        npu_inst_pe_1_0_5_n87) );
  NAND2_X1 npu_inst_pe_1_0_5_U58 ( .A1(npu_inst_pe_1_0_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_5_n40), .ZN(npu_inst_pe_1_0_5_n62) );
  OAI21_X1 npu_inst_pe_1_0_5_U57 ( .B1(npu_inst_pe_1_0_5_n61), .B2(
        npu_inst_pe_1_0_5_n40), .A(npu_inst_pe_1_0_5_n62), .ZN(
        npu_inst_pe_1_0_5_n86) );
  AOI22_X1 npu_inst_pe_1_0_5_U56 ( .A1(npu_inst_pe_1_0_5_n38), .A2(
        npu_inst_int_data_y_1__5__0_), .B1(npu_inst_pe_1_0_5_n113), .B2(
        npu_inst_pe_1_0_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_5_n37) );
  INV_X1 npu_inst_pe_1_0_5_U55 ( .A(npu_inst_pe_1_0_5_n37), .ZN(
        npu_inst_pe_1_0_5_n112) );
  AOI222_X1 npu_inst_pe_1_0_5_U54 ( .A1(npu_inst_int_data_res_1__5__0_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N73), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N65), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n84) );
  INV_X1 npu_inst_pe_1_0_5_U53 ( .A(npu_inst_pe_1_0_5_n84), .ZN(
        npu_inst_pe_1_0_5_n100) );
  AOI222_X1 npu_inst_pe_1_0_5_U52 ( .A1(npu_inst_pe_1_0_5_n1), .A2(
        npu_inst_int_data_res_1__5__7_), .B1(npu_inst_pe_1_0_5_N80), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N72), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n75) );
  INV_X1 npu_inst_pe_1_0_5_U51 ( .A(npu_inst_pe_1_0_5_n75), .ZN(
        npu_inst_pe_1_0_5_n32) );
  AOI222_X1 npu_inst_pe_1_0_5_U50 ( .A1(npu_inst_int_data_res_1__5__2_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N75), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N67), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n82) );
  INV_X1 npu_inst_pe_1_0_5_U49 ( .A(npu_inst_pe_1_0_5_n82), .ZN(
        npu_inst_pe_1_0_5_n98) );
  AOI222_X1 npu_inst_pe_1_0_5_U48 ( .A1(npu_inst_int_data_res_1__5__3_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N76), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N68), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n81) );
  INV_X1 npu_inst_pe_1_0_5_U47 ( .A(npu_inst_pe_1_0_5_n81), .ZN(
        npu_inst_pe_1_0_5_n36) );
  AOI222_X1 npu_inst_pe_1_0_5_U46 ( .A1(npu_inst_int_data_res_1__5__4_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N77), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N69), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n80) );
  INV_X1 npu_inst_pe_1_0_5_U45 ( .A(npu_inst_pe_1_0_5_n80), .ZN(
        npu_inst_pe_1_0_5_n35) );
  AOI222_X1 npu_inst_pe_1_0_5_U44 ( .A1(npu_inst_int_data_res_1__5__5_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N78), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N70), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n79) );
  INV_X1 npu_inst_pe_1_0_5_U43 ( .A(npu_inst_pe_1_0_5_n79), .ZN(
        npu_inst_pe_1_0_5_n34) );
  AOI222_X1 npu_inst_pe_1_0_5_U42 ( .A1(npu_inst_int_data_res_1__5__6_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N79), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N71), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n78) );
  INV_X1 npu_inst_pe_1_0_5_U41 ( .A(npu_inst_pe_1_0_5_n78), .ZN(
        npu_inst_pe_1_0_5_n33) );
  NOR3_X1 npu_inst_pe_1_0_5_U40 ( .A1(npu_inst_pe_1_0_5_n26), .A2(npu_inst_n42), .A3(npu_inst_int_ckg[58]), .ZN(npu_inst_pe_1_0_5_n85) );
  OR2_X1 npu_inst_pe_1_0_5_U39 ( .A1(npu_inst_pe_1_0_5_n85), .A2(
        npu_inst_pe_1_0_5_n1), .ZN(npu_inst_pe_1_0_5_N84) );
  AND2_X1 npu_inst_pe_1_0_5_U38 ( .A1(npu_inst_int_data_x_0__5__1_), .A2(
        npu_inst_pe_1_0_5_int_q_weight_1_), .ZN(npu_inst_pe_1_0_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_5_U37 ( .A1(npu_inst_int_data_x_0__5__0_), .A2(
        npu_inst_pe_1_0_5_int_q_weight_1_), .ZN(npu_inst_pe_1_0_5_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_0_5_U36 ( .A(npu_inst_pe_1_0_5_int_data_1_), .ZN(
        npu_inst_pe_1_0_5_n13) );
  AOI222_X1 npu_inst_pe_1_0_5_U35 ( .A1(npu_inst_int_data_res_1__5__1_), .A2(
        npu_inst_pe_1_0_5_n1), .B1(npu_inst_pe_1_0_5_N74), .B2(
        npu_inst_pe_1_0_5_n76), .C1(npu_inst_pe_1_0_5_N66), .C2(
        npu_inst_pe_1_0_5_n77), .ZN(npu_inst_pe_1_0_5_n83) );
  INV_X1 npu_inst_pe_1_0_5_U34 ( .A(npu_inst_pe_1_0_5_n83), .ZN(
        npu_inst_pe_1_0_5_n99) );
  AND2_X1 npu_inst_pe_1_0_5_U33 ( .A1(npu_inst_pe_1_0_5_N93), .A2(npu_inst_n42), .ZN(npu_inst_pe_1_0_5_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_5_U32 ( .A1(npu_inst_n42), .A2(npu_inst_pe_1_0_5_N94), .ZN(npu_inst_pe_1_0_5_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_5_U31 ( .A1(npu_inst_n42), .A2(
        npu_inst_int_data_y_1__5__1_), .B1(npu_inst_pe_1_0_5_n2), .B2(
        npu_inst_int_data_x_0__6__1_), .ZN(npu_inst_pe_1_0_5_n63) );
  AOI22_X1 npu_inst_pe_1_0_5_U30 ( .A1(npu_inst_n42), .A2(
        npu_inst_int_data_y_1__5__0_), .B1(npu_inst_pe_1_0_5_n2), .B2(
        npu_inst_int_data_x_0__6__0_), .ZN(npu_inst_pe_1_0_5_n61) );
  INV_X1 npu_inst_pe_1_0_5_U29 ( .A(npu_inst_pe_1_0_5_int_data_0_), .ZN(
        npu_inst_pe_1_0_5_n12) );
  INV_X1 npu_inst_pe_1_0_5_U28 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_0_5_n4)
         );
  OR3_X1 npu_inst_pe_1_0_5_U27 ( .A1(npu_inst_pe_1_0_5_n5), .A2(
        npu_inst_pe_1_0_5_n7), .A3(npu_inst_pe_1_0_5_n4), .ZN(
        npu_inst_pe_1_0_5_n56) );
  OR3_X1 npu_inst_pe_1_0_5_U26 ( .A1(npu_inst_pe_1_0_5_n4), .A2(
        npu_inst_pe_1_0_5_n7), .A3(npu_inst_pe_1_0_5_n6), .ZN(
        npu_inst_pe_1_0_5_n48) );
  INV_X1 npu_inst_pe_1_0_5_U25 ( .A(npu_inst_pe_1_0_5_n4), .ZN(
        npu_inst_pe_1_0_5_n3) );
  OR3_X1 npu_inst_pe_1_0_5_U24 ( .A1(npu_inst_pe_1_0_5_n3), .A2(
        npu_inst_pe_1_0_5_n7), .A3(npu_inst_pe_1_0_5_n6), .ZN(
        npu_inst_pe_1_0_5_n52) );
  OR3_X1 npu_inst_pe_1_0_5_U23 ( .A1(npu_inst_pe_1_0_5_n5), .A2(
        npu_inst_pe_1_0_5_n7), .A3(npu_inst_pe_1_0_5_n3), .ZN(
        npu_inst_pe_1_0_5_n60) );
  BUF_X1 npu_inst_pe_1_0_5_U22 ( .A(npu_inst_n30), .Z(npu_inst_pe_1_0_5_n1) );
  NOR2_X1 npu_inst_pe_1_0_5_U21 ( .A1(npu_inst_pe_1_0_5_n60), .A2(
        npu_inst_pe_1_0_5_n2), .ZN(npu_inst_pe_1_0_5_n58) );
  NOR2_X1 npu_inst_pe_1_0_5_U20 ( .A1(npu_inst_pe_1_0_5_n56), .A2(
        npu_inst_pe_1_0_5_n2), .ZN(npu_inst_pe_1_0_5_n54) );
  NOR2_X1 npu_inst_pe_1_0_5_U19 ( .A1(npu_inst_pe_1_0_5_n52), .A2(
        npu_inst_pe_1_0_5_n2), .ZN(npu_inst_pe_1_0_5_n50) );
  NOR2_X1 npu_inst_pe_1_0_5_U18 ( .A1(npu_inst_pe_1_0_5_n48), .A2(
        npu_inst_pe_1_0_5_n2), .ZN(npu_inst_pe_1_0_5_n46) );
  NOR2_X1 npu_inst_pe_1_0_5_U17 ( .A1(npu_inst_pe_1_0_5_n40), .A2(
        npu_inst_pe_1_0_5_n2), .ZN(npu_inst_pe_1_0_5_n38) );
  NOR2_X1 npu_inst_pe_1_0_5_U16 ( .A1(npu_inst_pe_1_0_5_n44), .A2(
        npu_inst_pe_1_0_5_n2), .ZN(npu_inst_pe_1_0_5_n42) );
  BUF_X1 npu_inst_pe_1_0_5_U15 ( .A(npu_inst_n88), .Z(npu_inst_pe_1_0_5_n7) );
  INV_X1 npu_inst_pe_1_0_5_U14 ( .A(npu_inst_n108), .ZN(npu_inst_pe_1_0_5_n11)
         );
  INV_X1 npu_inst_pe_1_0_5_U13 ( .A(npu_inst_pe_1_0_5_n38), .ZN(
        npu_inst_pe_1_0_5_n113) );
  INV_X1 npu_inst_pe_1_0_5_U12 ( .A(npu_inst_pe_1_0_5_n58), .ZN(
        npu_inst_pe_1_0_5_n118) );
  INV_X1 npu_inst_pe_1_0_5_U11 ( .A(npu_inst_pe_1_0_5_n54), .ZN(
        npu_inst_pe_1_0_5_n117) );
  INV_X1 npu_inst_pe_1_0_5_U10 ( .A(npu_inst_pe_1_0_5_n50), .ZN(
        npu_inst_pe_1_0_5_n116) );
  INV_X1 npu_inst_pe_1_0_5_U9 ( .A(npu_inst_pe_1_0_5_n46), .ZN(
        npu_inst_pe_1_0_5_n115) );
  INV_X1 npu_inst_pe_1_0_5_U8 ( .A(npu_inst_pe_1_0_5_n42), .ZN(
        npu_inst_pe_1_0_5_n114) );
  BUF_X1 npu_inst_pe_1_0_5_U7 ( .A(npu_inst_pe_1_0_5_n11), .Z(
        npu_inst_pe_1_0_5_n10) );
  BUF_X1 npu_inst_pe_1_0_5_U6 ( .A(npu_inst_pe_1_0_5_n11), .Z(
        npu_inst_pe_1_0_5_n9) );
  BUF_X1 npu_inst_pe_1_0_5_U5 ( .A(npu_inst_pe_1_0_5_n11), .Z(
        npu_inst_pe_1_0_5_n8) );
  NOR2_X1 npu_inst_pe_1_0_5_U4 ( .A1(npu_inst_pe_1_0_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_5_n1), .ZN(npu_inst_pe_1_0_5_n76) );
  NOR2_X1 npu_inst_pe_1_0_5_U3 ( .A1(npu_inst_pe_1_0_5_n27), .A2(
        npu_inst_pe_1_0_5_n1), .ZN(npu_inst_pe_1_0_5_n77) );
  FA_X1 npu_inst_pe_1_0_5_sub_77_U2_1 ( .A(int_o_data_npu[17]), .B(
        npu_inst_pe_1_0_5_n13), .CI(npu_inst_pe_1_0_5_sub_77_carry_1_), .CO(
        npu_inst_pe_1_0_5_sub_77_carry_2_), .S(npu_inst_pe_1_0_5_N66) );
  FA_X1 npu_inst_pe_1_0_5_add_79_U1_1 ( .A(int_o_data_npu[17]), .B(
        npu_inst_pe_1_0_5_int_data_1_), .CI(npu_inst_pe_1_0_5_add_79_carry_1_), 
        .CO(npu_inst_pe_1_0_5_add_79_carry_2_), .S(npu_inst_pe_1_0_5_N74) );
  NAND3_X1 npu_inst_pe_1_0_5_U101 ( .A1(npu_inst_pe_1_0_5_n4), .A2(
        npu_inst_pe_1_0_5_n6), .A3(npu_inst_pe_1_0_5_n7), .ZN(
        npu_inst_pe_1_0_5_n44) );
  NAND3_X1 npu_inst_pe_1_0_5_U100 ( .A1(npu_inst_pe_1_0_5_n3), .A2(
        npu_inst_pe_1_0_5_n6), .A3(npu_inst_pe_1_0_5_n7), .ZN(
        npu_inst_pe_1_0_5_n40) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_5_n33), .CK(
        npu_inst_pe_1_0_5_net4363), .RN(npu_inst_pe_1_0_5_n8), .Q(
        int_o_data_npu[22]) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_5_n34), .CK(
        npu_inst_pe_1_0_5_net4363), .RN(npu_inst_pe_1_0_5_n8), .Q(
        int_o_data_npu[21]) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_5_n35), .CK(
        npu_inst_pe_1_0_5_net4363), .RN(npu_inst_pe_1_0_5_n8), .Q(
        int_o_data_npu[20]) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_5_n36), .CK(
        npu_inst_pe_1_0_5_net4363), .RN(npu_inst_pe_1_0_5_n8), .Q(
        int_o_data_npu[19]) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_5_n98), .CK(
        npu_inst_pe_1_0_5_net4363), .RN(npu_inst_pe_1_0_5_n8), .Q(
        int_o_data_npu[18]) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_5_n99), .CK(
        npu_inst_pe_1_0_5_net4363), .RN(npu_inst_pe_1_0_5_n8), .Q(
        int_o_data_npu[17]) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_5_n32), .CK(
        npu_inst_pe_1_0_5_net4363), .RN(npu_inst_pe_1_0_5_n8), .Q(
        int_o_data_npu[23]) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_5_n100), 
        .CK(npu_inst_pe_1_0_5_net4363), .RN(npu_inst_pe_1_0_5_n8), .Q(
        int_o_data_npu[16]) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_weight_reg_0_ ( .D(npu_inst_n94), .CK(
        npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n8), .Q(
        npu_inst_pe_1_0_5_int_q_weight_0_), .QN(npu_inst_pe_1_0_5_n27) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_weight_reg_1_ ( .D(npu_inst_n100), .CK(
        npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n8), .Q(
        npu_inst_pe_1_0_5_int_q_weight_1_), .QN(npu_inst_pe_1_0_5_n26) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_5_n112), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n8), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_5_n106), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n8), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_5_n111), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_5_n105), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_5_n110), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_5_n104), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_5_n109), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_5_n103), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_5_n108), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_5_n102), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_5_n107), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_5_n101), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_5_n86), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_5_n87), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n9), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_5_n88), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_5_n89), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_5_n90), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_5_n91), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_5_n92), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_5_n93), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_5_n94), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_5_n95), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_5_n96), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_5_n97), 
        .CK(npu_inst_pe_1_0_5_net4369), .RN(npu_inst_pe_1_0_5_n10), .Q(
        npu_inst_pe_1_0_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_5_net4363) );
  CLKGATETST_X1 npu_inst_pe_1_0_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n48), .SE(1'b0), .GCK(npu_inst_pe_1_0_5_net4369) );
  MUX2_X1 npu_inst_pe_1_0_6_U153 ( .A(npu_inst_pe_1_0_6_n31), .B(
        npu_inst_pe_1_0_6_n28), .S(npu_inst_pe_1_0_6_n7), .Z(
        npu_inst_pe_1_0_6_N93) );
  MUX2_X1 npu_inst_pe_1_0_6_U152 ( .A(npu_inst_pe_1_0_6_n30), .B(
        npu_inst_pe_1_0_6_n29), .S(npu_inst_pe_1_0_6_n5), .Z(
        npu_inst_pe_1_0_6_n31) );
  MUX2_X1 npu_inst_pe_1_0_6_U151 ( .A(npu_inst_pe_1_0_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_6_n3), .Z(
        npu_inst_pe_1_0_6_n30) );
  MUX2_X1 npu_inst_pe_1_0_6_U150 ( .A(npu_inst_pe_1_0_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_6_n3), .Z(
        npu_inst_pe_1_0_6_n29) );
  MUX2_X1 npu_inst_pe_1_0_6_U149 ( .A(npu_inst_pe_1_0_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_6_n3), .Z(
        npu_inst_pe_1_0_6_n28) );
  MUX2_X1 npu_inst_pe_1_0_6_U148 ( .A(npu_inst_pe_1_0_6_n25), .B(
        npu_inst_pe_1_0_6_n22), .S(npu_inst_pe_1_0_6_n7), .Z(
        npu_inst_pe_1_0_6_N94) );
  MUX2_X1 npu_inst_pe_1_0_6_U147 ( .A(npu_inst_pe_1_0_6_n24), .B(
        npu_inst_pe_1_0_6_n23), .S(npu_inst_pe_1_0_6_n5), .Z(
        npu_inst_pe_1_0_6_n25) );
  MUX2_X1 npu_inst_pe_1_0_6_U146 ( .A(npu_inst_pe_1_0_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_6_n3), .Z(
        npu_inst_pe_1_0_6_n24) );
  MUX2_X1 npu_inst_pe_1_0_6_U145 ( .A(npu_inst_pe_1_0_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_6_n3), .Z(
        npu_inst_pe_1_0_6_n23) );
  MUX2_X1 npu_inst_pe_1_0_6_U144 ( .A(npu_inst_pe_1_0_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_6_n3), .Z(
        npu_inst_pe_1_0_6_n22) );
  MUX2_X1 npu_inst_pe_1_0_6_U143 ( .A(npu_inst_pe_1_0_6_n21), .B(
        npu_inst_pe_1_0_6_n18), .S(npu_inst_pe_1_0_6_n7), .Z(
        npu_inst_int_data_x_0__6__1_) );
  MUX2_X1 npu_inst_pe_1_0_6_U142 ( .A(npu_inst_pe_1_0_6_n20), .B(
        npu_inst_pe_1_0_6_n19), .S(npu_inst_pe_1_0_6_n5), .Z(
        npu_inst_pe_1_0_6_n21) );
  MUX2_X1 npu_inst_pe_1_0_6_U141 ( .A(npu_inst_pe_1_0_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_6_n3), .Z(
        npu_inst_pe_1_0_6_n20) );
  MUX2_X1 npu_inst_pe_1_0_6_U140 ( .A(npu_inst_pe_1_0_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_6_n3), .Z(
        npu_inst_pe_1_0_6_n19) );
  MUX2_X1 npu_inst_pe_1_0_6_U139 ( .A(npu_inst_pe_1_0_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_6_n3), .Z(
        npu_inst_pe_1_0_6_n18) );
  MUX2_X1 npu_inst_pe_1_0_6_U138 ( .A(npu_inst_pe_1_0_6_n17), .B(
        npu_inst_pe_1_0_6_n14), .S(npu_inst_pe_1_0_6_n7), .Z(
        npu_inst_int_data_x_0__6__0_) );
  MUX2_X1 npu_inst_pe_1_0_6_U137 ( .A(npu_inst_pe_1_0_6_n16), .B(
        npu_inst_pe_1_0_6_n15), .S(npu_inst_pe_1_0_6_n5), .Z(
        npu_inst_pe_1_0_6_n17) );
  MUX2_X1 npu_inst_pe_1_0_6_U136 ( .A(npu_inst_pe_1_0_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_6_n3), .Z(
        npu_inst_pe_1_0_6_n16) );
  MUX2_X1 npu_inst_pe_1_0_6_U135 ( .A(npu_inst_pe_1_0_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_6_n3), .Z(
        npu_inst_pe_1_0_6_n15) );
  MUX2_X1 npu_inst_pe_1_0_6_U134 ( .A(npu_inst_pe_1_0_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_6_n3), .Z(
        npu_inst_pe_1_0_6_n14) );
  XOR2_X1 npu_inst_pe_1_0_6_U133 ( .A(npu_inst_pe_1_0_6_int_data_0_), .B(
        int_o_data_npu[8]), .Z(npu_inst_pe_1_0_6_N73) );
  AND2_X1 npu_inst_pe_1_0_6_U132 ( .A1(int_o_data_npu[8]), .A2(
        npu_inst_pe_1_0_6_int_data_0_), .ZN(npu_inst_pe_1_0_6_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_6_U131 ( .A(int_o_data_npu[8]), .B(
        npu_inst_pe_1_0_6_n12), .ZN(npu_inst_pe_1_0_6_N65) );
  OR2_X1 npu_inst_pe_1_0_6_U130 ( .A1(npu_inst_pe_1_0_6_n12), .A2(
        int_o_data_npu[8]), .ZN(npu_inst_pe_1_0_6_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_6_U129 ( .A(int_o_data_npu[10]), .B(
        npu_inst_pe_1_0_6_add_79_carry_2_), .Z(npu_inst_pe_1_0_6_N75) );
  AND2_X1 npu_inst_pe_1_0_6_U128 ( .A1(npu_inst_pe_1_0_6_add_79_carry_2_), 
        .A2(int_o_data_npu[10]), .ZN(npu_inst_pe_1_0_6_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_6_U127 ( .A(int_o_data_npu[11]), .B(
        npu_inst_pe_1_0_6_add_79_carry_3_), .Z(npu_inst_pe_1_0_6_N76) );
  AND2_X1 npu_inst_pe_1_0_6_U126 ( .A1(npu_inst_pe_1_0_6_add_79_carry_3_), 
        .A2(int_o_data_npu[11]), .ZN(npu_inst_pe_1_0_6_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_6_U125 ( .A(int_o_data_npu[12]), .B(
        npu_inst_pe_1_0_6_add_79_carry_4_), .Z(npu_inst_pe_1_0_6_N77) );
  AND2_X1 npu_inst_pe_1_0_6_U124 ( .A1(npu_inst_pe_1_0_6_add_79_carry_4_), 
        .A2(int_o_data_npu[12]), .ZN(npu_inst_pe_1_0_6_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_6_U123 ( .A(int_o_data_npu[13]), .B(
        npu_inst_pe_1_0_6_add_79_carry_5_), .Z(npu_inst_pe_1_0_6_N78) );
  AND2_X1 npu_inst_pe_1_0_6_U122 ( .A1(npu_inst_pe_1_0_6_add_79_carry_5_), 
        .A2(int_o_data_npu[13]), .ZN(npu_inst_pe_1_0_6_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_6_U121 ( .A(int_o_data_npu[14]), .B(
        npu_inst_pe_1_0_6_add_79_carry_6_), .Z(npu_inst_pe_1_0_6_N79) );
  AND2_X1 npu_inst_pe_1_0_6_U120 ( .A1(npu_inst_pe_1_0_6_add_79_carry_6_), 
        .A2(int_o_data_npu[14]), .ZN(npu_inst_pe_1_0_6_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_6_U119 ( .A(int_o_data_npu[15]), .B(
        npu_inst_pe_1_0_6_add_79_carry_7_), .Z(npu_inst_pe_1_0_6_N80) );
  XNOR2_X1 npu_inst_pe_1_0_6_U118 ( .A(npu_inst_pe_1_0_6_sub_77_carry_2_), .B(
        int_o_data_npu[10]), .ZN(npu_inst_pe_1_0_6_N67) );
  OR2_X1 npu_inst_pe_1_0_6_U117 ( .A1(int_o_data_npu[10]), .A2(
        npu_inst_pe_1_0_6_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_0_6_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_6_U116 ( .A(npu_inst_pe_1_0_6_sub_77_carry_3_), .B(
        int_o_data_npu[11]), .ZN(npu_inst_pe_1_0_6_N68) );
  OR2_X1 npu_inst_pe_1_0_6_U115 ( .A1(int_o_data_npu[11]), .A2(
        npu_inst_pe_1_0_6_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_0_6_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_6_U114 ( .A(npu_inst_pe_1_0_6_sub_77_carry_4_), .B(
        int_o_data_npu[12]), .ZN(npu_inst_pe_1_0_6_N69) );
  OR2_X1 npu_inst_pe_1_0_6_U113 ( .A1(int_o_data_npu[12]), .A2(
        npu_inst_pe_1_0_6_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_0_6_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_6_U112 ( .A(npu_inst_pe_1_0_6_sub_77_carry_5_), .B(
        int_o_data_npu[13]), .ZN(npu_inst_pe_1_0_6_N70) );
  OR2_X1 npu_inst_pe_1_0_6_U111 ( .A1(int_o_data_npu[13]), .A2(
        npu_inst_pe_1_0_6_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_0_6_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_6_U110 ( .A(npu_inst_pe_1_0_6_sub_77_carry_6_), .B(
        int_o_data_npu[14]), .ZN(npu_inst_pe_1_0_6_N71) );
  OR2_X1 npu_inst_pe_1_0_6_U109 ( .A1(int_o_data_npu[14]), .A2(
        npu_inst_pe_1_0_6_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_0_6_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_6_U108 ( .A(int_o_data_npu[15]), .B(
        npu_inst_pe_1_0_6_sub_77_carry_7_), .ZN(npu_inst_pe_1_0_6_N72) );
  INV_X1 npu_inst_pe_1_0_6_U107 ( .A(npu_inst_n61), .ZN(npu_inst_pe_1_0_6_n6)
         );
  INV_X1 npu_inst_pe_1_0_6_U106 ( .A(npu_inst_pe_1_0_6_n6), .ZN(
        npu_inst_pe_1_0_6_n5) );
  INV_X1 npu_inst_pe_1_0_6_U105 ( .A(npu_inst_n42), .ZN(npu_inst_pe_1_0_6_n2)
         );
  AOI22_X1 npu_inst_pe_1_0_6_U104 ( .A1(npu_inst_int_data_y_1__6__0_), .A2(
        npu_inst_pe_1_0_6_n58), .B1(npu_inst_pe_1_0_6_n118), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_6_n57) );
  INV_X1 npu_inst_pe_1_0_6_U103 ( .A(npu_inst_pe_1_0_6_n57), .ZN(
        npu_inst_pe_1_0_6_n107) );
  AOI22_X1 npu_inst_pe_1_0_6_U102 ( .A1(npu_inst_int_data_y_1__6__0_), .A2(
        npu_inst_pe_1_0_6_n54), .B1(npu_inst_pe_1_0_6_n117), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_6_n53) );
  INV_X1 npu_inst_pe_1_0_6_U99 ( .A(npu_inst_pe_1_0_6_n53), .ZN(
        npu_inst_pe_1_0_6_n108) );
  AOI22_X1 npu_inst_pe_1_0_6_U98 ( .A1(npu_inst_int_data_y_1__6__0_), .A2(
        npu_inst_pe_1_0_6_n50), .B1(npu_inst_pe_1_0_6_n116), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_6_n49) );
  INV_X1 npu_inst_pe_1_0_6_U97 ( .A(npu_inst_pe_1_0_6_n49), .ZN(
        npu_inst_pe_1_0_6_n109) );
  AOI22_X1 npu_inst_pe_1_0_6_U96 ( .A1(npu_inst_int_data_y_1__6__0_), .A2(
        npu_inst_pe_1_0_6_n46), .B1(npu_inst_pe_1_0_6_n115), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_6_n45) );
  INV_X1 npu_inst_pe_1_0_6_U95 ( .A(npu_inst_pe_1_0_6_n45), .ZN(
        npu_inst_pe_1_0_6_n110) );
  AOI22_X1 npu_inst_pe_1_0_6_U94 ( .A1(npu_inst_int_data_y_1__6__0_), .A2(
        npu_inst_pe_1_0_6_n42), .B1(npu_inst_pe_1_0_6_n114), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_6_n41) );
  INV_X1 npu_inst_pe_1_0_6_U93 ( .A(npu_inst_pe_1_0_6_n41), .ZN(
        npu_inst_pe_1_0_6_n111) );
  AOI22_X1 npu_inst_pe_1_0_6_U92 ( .A1(npu_inst_int_data_y_1__6__1_), .A2(
        npu_inst_pe_1_0_6_n58), .B1(npu_inst_pe_1_0_6_n118), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_6_n59) );
  INV_X1 npu_inst_pe_1_0_6_U91 ( .A(npu_inst_pe_1_0_6_n59), .ZN(
        npu_inst_pe_1_0_6_n101) );
  AOI22_X1 npu_inst_pe_1_0_6_U90 ( .A1(npu_inst_int_data_y_1__6__1_), .A2(
        npu_inst_pe_1_0_6_n54), .B1(npu_inst_pe_1_0_6_n117), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_6_n55) );
  INV_X1 npu_inst_pe_1_0_6_U89 ( .A(npu_inst_pe_1_0_6_n55), .ZN(
        npu_inst_pe_1_0_6_n102) );
  AOI22_X1 npu_inst_pe_1_0_6_U88 ( .A1(npu_inst_int_data_y_1__6__1_), .A2(
        npu_inst_pe_1_0_6_n50), .B1(npu_inst_pe_1_0_6_n116), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_6_n51) );
  INV_X1 npu_inst_pe_1_0_6_U87 ( .A(npu_inst_pe_1_0_6_n51), .ZN(
        npu_inst_pe_1_0_6_n103) );
  AOI22_X1 npu_inst_pe_1_0_6_U86 ( .A1(npu_inst_int_data_y_1__6__1_), .A2(
        npu_inst_pe_1_0_6_n46), .B1(npu_inst_pe_1_0_6_n115), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_6_n47) );
  INV_X1 npu_inst_pe_1_0_6_U85 ( .A(npu_inst_pe_1_0_6_n47), .ZN(
        npu_inst_pe_1_0_6_n104) );
  AOI22_X1 npu_inst_pe_1_0_6_U84 ( .A1(npu_inst_int_data_y_1__6__1_), .A2(
        npu_inst_pe_1_0_6_n42), .B1(npu_inst_pe_1_0_6_n114), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_6_n43) );
  INV_X1 npu_inst_pe_1_0_6_U83 ( .A(npu_inst_pe_1_0_6_n43), .ZN(
        npu_inst_pe_1_0_6_n105) );
  AOI22_X1 npu_inst_pe_1_0_6_U82 ( .A1(npu_inst_pe_1_0_6_n38), .A2(
        npu_inst_int_data_y_1__6__1_), .B1(npu_inst_pe_1_0_6_n113), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_6_n39) );
  INV_X1 npu_inst_pe_1_0_6_U81 ( .A(npu_inst_pe_1_0_6_n39), .ZN(
        npu_inst_pe_1_0_6_n106) );
  NAND2_X1 npu_inst_pe_1_0_6_U80 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_6_n60), .ZN(npu_inst_pe_1_0_6_n74) );
  OAI21_X1 npu_inst_pe_1_0_6_U79 ( .B1(npu_inst_pe_1_0_6_n63), .B2(
        npu_inst_pe_1_0_6_n60), .A(npu_inst_pe_1_0_6_n74), .ZN(
        npu_inst_pe_1_0_6_n97) );
  NAND2_X1 npu_inst_pe_1_0_6_U78 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_6_n60), .ZN(npu_inst_pe_1_0_6_n73) );
  OAI21_X1 npu_inst_pe_1_0_6_U77 ( .B1(npu_inst_pe_1_0_6_n61), .B2(
        npu_inst_pe_1_0_6_n60), .A(npu_inst_pe_1_0_6_n73), .ZN(
        npu_inst_pe_1_0_6_n96) );
  NAND2_X1 npu_inst_pe_1_0_6_U76 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_6_n56), .ZN(npu_inst_pe_1_0_6_n72) );
  OAI21_X1 npu_inst_pe_1_0_6_U75 ( .B1(npu_inst_pe_1_0_6_n63), .B2(
        npu_inst_pe_1_0_6_n56), .A(npu_inst_pe_1_0_6_n72), .ZN(
        npu_inst_pe_1_0_6_n95) );
  NAND2_X1 npu_inst_pe_1_0_6_U74 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_6_n56), .ZN(npu_inst_pe_1_0_6_n71) );
  OAI21_X1 npu_inst_pe_1_0_6_U73 ( .B1(npu_inst_pe_1_0_6_n61), .B2(
        npu_inst_pe_1_0_6_n56), .A(npu_inst_pe_1_0_6_n71), .ZN(
        npu_inst_pe_1_0_6_n94) );
  NAND2_X1 npu_inst_pe_1_0_6_U72 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_6_n52), .ZN(npu_inst_pe_1_0_6_n70) );
  OAI21_X1 npu_inst_pe_1_0_6_U71 ( .B1(npu_inst_pe_1_0_6_n63), .B2(
        npu_inst_pe_1_0_6_n52), .A(npu_inst_pe_1_0_6_n70), .ZN(
        npu_inst_pe_1_0_6_n93) );
  NAND2_X1 npu_inst_pe_1_0_6_U70 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_6_n52), .ZN(npu_inst_pe_1_0_6_n69) );
  OAI21_X1 npu_inst_pe_1_0_6_U69 ( .B1(npu_inst_pe_1_0_6_n61), .B2(
        npu_inst_pe_1_0_6_n52), .A(npu_inst_pe_1_0_6_n69), .ZN(
        npu_inst_pe_1_0_6_n92) );
  NAND2_X1 npu_inst_pe_1_0_6_U68 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_6_n48), .ZN(npu_inst_pe_1_0_6_n68) );
  OAI21_X1 npu_inst_pe_1_0_6_U67 ( .B1(npu_inst_pe_1_0_6_n63), .B2(
        npu_inst_pe_1_0_6_n48), .A(npu_inst_pe_1_0_6_n68), .ZN(
        npu_inst_pe_1_0_6_n91) );
  NAND2_X1 npu_inst_pe_1_0_6_U66 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_6_n48), .ZN(npu_inst_pe_1_0_6_n67) );
  OAI21_X1 npu_inst_pe_1_0_6_U65 ( .B1(npu_inst_pe_1_0_6_n61), .B2(
        npu_inst_pe_1_0_6_n48), .A(npu_inst_pe_1_0_6_n67), .ZN(
        npu_inst_pe_1_0_6_n90) );
  NAND2_X1 npu_inst_pe_1_0_6_U64 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_6_n44), .ZN(npu_inst_pe_1_0_6_n66) );
  OAI21_X1 npu_inst_pe_1_0_6_U63 ( .B1(npu_inst_pe_1_0_6_n63), .B2(
        npu_inst_pe_1_0_6_n44), .A(npu_inst_pe_1_0_6_n66), .ZN(
        npu_inst_pe_1_0_6_n89) );
  NAND2_X1 npu_inst_pe_1_0_6_U62 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_6_n44), .ZN(npu_inst_pe_1_0_6_n65) );
  OAI21_X1 npu_inst_pe_1_0_6_U61 ( .B1(npu_inst_pe_1_0_6_n61), .B2(
        npu_inst_pe_1_0_6_n44), .A(npu_inst_pe_1_0_6_n65), .ZN(
        npu_inst_pe_1_0_6_n88) );
  NAND2_X1 npu_inst_pe_1_0_6_U60 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_6_n40), .ZN(npu_inst_pe_1_0_6_n64) );
  OAI21_X1 npu_inst_pe_1_0_6_U59 ( .B1(npu_inst_pe_1_0_6_n63), .B2(
        npu_inst_pe_1_0_6_n40), .A(npu_inst_pe_1_0_6_n64), .ZN(
        npu_inst_pe_1_0_6_n87) );
  NAND2_X1 npu_inst_pe_1_0_6_U58 ( .A1(npu_inst_pe_1_0_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_6_n40), .ZN(npu_inst_pe_1_0_6_n62) );
  OAI21_X1 npu_inst_pe_1_0_6_U57 ( .B1(npu_inst_pe_1_0_6_n61), .B2(
        npu_inst_pe_1_0_6_n40), .A(npu_inst_pe_1_0_6_n62), .ZN(
        npu_inst_pe_1_0_6_n86) );
  AOI22_X1 npu_inst_pe_1_0_6_U56 ( .A1(npu_inst_pe_1_0_6_n38), .A2(
        npu_inst_int_data_y_1__6__0_), .B1(npu_inst_pe_1_0_6_n113), .B2(
        npu_inst_pe_1_0_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_6_n37) );
  INV_X1 npu_inst_pe_1_0_6_U55 ( .A(npu_inst_pe_1_0_6_n37), .ZN(
        npu_inst_pe_1_0_6_n112) );
  AOI222_X1 npu_inst_pe_1_0_6_U54 ( .A1(npu_inst_int_data_res_1__6__0_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N73), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N65), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n84) );
  INV_X1 npu_inst_pe_1_0_6_U53 ( .A(npu_inst_pe_1_0_6_n84), .ZN(
        npu_inst_pe_1_0_6_n100) );
  AOI222_X1 npu_inst_pe_1_0_6_U52 ( .A1(npu_inst_pe_1_0_6_n1), .A2(
        npu_inst_int_data_res_1__6__7_), .B1(npu_inst_pe_1_0_6_N80), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N72), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n75) );
  INV_X1 npu_inst_pe_1_0_6_U51 ( .A(npu_inst_pe_1_0_6_n75), .ZN(
        npu_inst_pe_1_0_6_n32) );
  AOI222_X1 npu_inst_pe_1_0_6_U50 ( .A1(npu_inst_int_data_res_1__6__2_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N75), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N67), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n82) );
  INV_X1 npu_inst_pe_1_0_6_U49 ( .A(npu_inst_pe_1_0_6_n82), .ZN(
        npu_inst_pe_1_0_6_n98) );
  AOI222_X1 npu_inst_pe_1_0_6_U48 ( .A1(npu_inst_int_data_res_1__6__3_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N76), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N68), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n81) );
  INV_X1 npu_inst_pe_1_0_6_U47 ( .A(npu_inst_pe_1_0_6_n81), .ZN(
        npu_inst_pe_1_0_6_n36) );
  AOI222_X1 npu_inst_pe_1_0_6_U46 ( .A1(npu_inst_int_data_res_1__6__4_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N77), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N69), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n80) );
  INV_X1 npu_inst_pe_1_0_6_U45 ( .A(npu_inst_pe_1_0_6_n80), .ZN(
        npu_inst_pe_1_0_6_n35) );
  AOI222_X1 npu_inst_pe_1_0_6_U44 ( .A1(npu_inst_int_data_res_1__6__5_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N78), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N70), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n79) );
  INV_X1 npu_inst_pe_1_0_6_U43 ( .A(npu_inst_pe_1_0_6_n79), .ZN(
        npu_inst_pe_1_0_6_n34) );
  AOI222_X1 npu_inst_pe_1_0_6_U42 ( .A1(npu_inst_int_data_res_1__6__6_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N79), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N71), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n78) );
  INV_X1 npu_inst_pe_1_0_6_U41 ( .A(npu_inst_pe_1_0_6_n78), .ZN(
        npu_inst_pe_1_0_6_n33) );
  AND2_X1 npu_inst_pe_1_0_6_U40 ( .A1(npu_inst_int_data_x_0__6__1_), .A2(
        npu_inst_pe_1_0_6_int_q_weight_1_), .ZN(npu_inst_pe_1_0_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_6_U39 ( .A1(npu_inst_int_data_x_0__6__0_), .A2(
        npu_inst_pe_1_0_6_int_q_weight_1_), .ZN(npu_inst_pe_1_0_6_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_0_6_U38 ( .A(npu_inst_pe_1_0_6_int_data_1_), .ZN(
        npu_inst_pe_1_0_6_n13) );
  NOR3_X1 npu_inst_pe_1_0_6_U37 ( .A1(npu_inst_pe_1_0_6_n26), .A2(npu_inst_n42), .A3(npu_inst_int_ckg[57]), .ZN(npu_inst_pe_1_0_6_n85) );
  OR2_X1 npu_inst_pe_1_0_6_U36 ( .A1(npu_inst_pe_1_0_6_n85), .A2(
        npu_inst_pe_1_0_6_n1), .ZN(npu_inst_pe_1_0_6_N84) );
  AOI222_X1 npu_inst_pe_1_0_6_U35 ( .A1(npu_inst_int_data_res_1__6__1_), .A2(
        npu_inst_pe_1_0_6_n1), .B1(npu_inst_pe_1_0_6_N74), .B2(
        npu_inst_pe_1_0_6_n76), .C1(npu_inst_pe_1_0_6_N66), .C2(
        npu_inst_pe_1_0_6_n77), .ZN(npu_inst_pe_1_0_6_n83) );
  INV_X1 npu_inst_pe_1_0_6_U34 ( .A(npu_inst_pe_1_0_6_n83), .ZN(
        npu_inst_pe_1_0_6_n99) );
  AND2_X1 npu_inst_pe_1_0_6_U33 ( .A1(npu_inst_pe_1_0_6_N93), .A2(npu_inst_n42), .ZN(npu_inst_pe_1_0_6_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_6_U32 ( .A1(npu_inst_n42), .A2(npu_inst_pe_1_0_6_N94), .ZN(npu_inst_pe_1_0_6_o_data_v_1_) );
  AOI22_X1 npu_inst_pe_1_0_6_U31 ( .A1(npu_inst_n42), .A2(
        npu_inst_int_data_y_1__6__1_), .B1(npu_inst_pe_1_0_6_n2), .B2(
        npu_inst_int_data_x_0__7__1_), .ZN(npu_inst_pe_1_0_6_n63) );
  AOI22_X1 npu_inst_pe_1_0_6_U30 ( .A1(npu_inst_n42), .A2(
        npu_inst_int_data_y_1__6__0_), .B1(npu_inst_pe_1_0_6_n2), .B2(
        npu_inst_int_data_x_0__7__0_), .ZN(npu_inst_pe_1_0_6_n61) );
  INV_X1 npu_inst_pe_1_0_6_U29 ( .A(npu_inst_pe_1_0_6_int_data_0_), .ZN(
        npu_inst_pe_1_0_6_n12) );
  INV_X1 npu_inst_pe_1_0_6_U28 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_0_6_n4)
         );
  OR3_X1 npu_inst_pe_1_0_6_U27 ( .A1(npu_inst_pe_1_0_6_n5), .A2(
        npu_inst_pe_1_0_6_n7), .A3(npu_inst_pe_1_0_6_n4), .ZN(
        npu_inst_pe_1_0_6_n56) );
  OR3_X1 npu_inst_pe_1_0_6_U26 ( .A1(npu_inst_pe_1_0_6_n4), .A2(
        npu_inst_pe_1_0_6_n7), .A3(npu_inst_pe_1_0_6_n6), .ZN(
        npu_inst_pe_1_0_6_n48) );
  INV_X1 npu_inst_pe_1_0_6_U25 ( .A(npu_inst_pe_1_0_6_n4), .ZN(
        npu_inst_pe_1_0_6_n3) );
  OR3_X1 npu_inst_pe_1_0_6_U24 ( .A1(npu_inst_pe_1_0_6_n3), .A2(
        npu_inst_pe_1_0_6_n7), .A3(npu_inst_pe_1_0_6_n6), .ZN(
        npu_inst_pe_1_0_6_n52) );
  OR3_X1 npu_inst_pe_1_0_6_U23 ( .A1(npu_inst_pe_1_0_6_n5), .A2(
        npu_inst_pe_1_0_6_n7), .A3(npu_inst_pe_1_0_6_n3), .ZN(
        npu_inst_pe_1_0_6_n60) );
  BUF_X1 npu_inst_pe_1_0_6_U22 ( .A(npu_inst_n30), .Z(npu_inst_pe_1_0_6_n1) );
  NOR2_X1 npu_inst_pe_1_0_6_U21 ( .A1(npu_inst_pe_1_0_6_n60), .A2(
        npu_inst_pe_1_0_6_n2), .ZN(npu_inst_pe_1_0_6_n58) );
  NOR2_X1 npu_inst_pe_1_0_6_U20 ( .A1(npu_inst_pe_1_0_6_n56), .A2(
        npu_inst_pe_1_0_6_n2), .ZN(npu_inst_pe_1_0_6_n54) );
  NOR2_X1 npu_inst_pe_1_0_6_U19 ( .A1(npu_inst_pe_1_0_6_n52), .A2(
        npu_inst_pe_1_0_6_n2), .ZN(npu_inst_pe_1_0_6_n50) );
  NOR2_X1 npu_inst_pe_1_0_6_U18 ( .A1(npu_inst_pe_1_0_6_n48), .A2(
        npu_inst_pe_1_0_6_n2), .ZN(npu_inst_pe_1_0_6_n46) );
  NOR2_X1 npu_inst_pe_1_0_6_U17 ( .A1(npu_inst_pe_1_0_6_n40), .A2(
        npu_inst_pe_1_0_6_n2), .ZN(npu_inst_pe_1_0_6_n38) );
  NOR2_X1 npu_inst_pe_1_0_6_U16 ( .A1(npu_inst_pe_1_0_6_n44), .A2(
        npu_inst_pe_1_0_6_n2), .ZN(npu_inst_pe_1_0_6_n42) );
  BUF_X1 npu_inst_pe_1_0_6_U15 ( .A(npu_inst_n88), .Z(npu_inst_pe_1_0_6_n7) );
  INV_X1 npu_inst_pe_1_0_6_U14 ( .A(npu_inst_n108), .ZN(npu_inst_pe_1_0_6_n11)
         );
  INV_X1 npu_inst_pe_1_0_6_U13 ( .A(npu_inst_pe_1_0_6_n38), .ZN(
        npu_inst_pe_1_0_6_n113) );
  INV_X1 npu_inst_pe_1_0_6_U12 ( .A(npu_inst_pe_1_0_6_n58), .ZN(
        npu_inst_pe_1_0_6_n118) );
  INV_X1 npu_inst_pe_1_0_6_U11 ( .A(npu_inst_pe_1_0_6_n54), .ZN(
        npu_inst_pe_1_0_6_n117) );
  INV_X1 npu_inst_pe_1_0_6_U10 ( .A(npu_inst_pe_1_0_6_n50), .ZN(
        npu_inst_pe_1_0_6_n116) );
  INV_X1 npu_inst_pe_1_0_6_U9 ( .A(npu_inst_pe_1_0_6_n46), .ZN(
        npu_inst_pe_1_0_6_n115) );
  INV_X1 npu_inst_pe_1_0_6_U8 ( .A(npu_inst_pe_1_0_6_n42), .ZN(
        npu_inst_pe_1_0_6_n114) );
  BUF_X1 npu_inst_pe_1_0_6_U7 ( .A(npu_inst_pe_1_0_6_n11), .Z(
        npu_inst_pe_1_0_6_n10) );
  BUF_X1 npu_inst_pe_1_0_6_U6 ( .A(npu_inst_pe_1_0_6_n11), .Z(
        npu_inst_pe_1_0_6_n9) );
  BUF_X1 npu_inst_pe_1_0_6_U5 ( .A(npu_inst_pe_1_0_6_n11), .Z(
        npu_inst_pe_1_0_6_n8) );
  NOR2_X1 npu_inst_pe_1_0_6_U4 ( .A1(npu_inst_pe_1_0_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_6_n1), .ZN(npu_inst_pe_1_0_6_n76) );
  NOR2_X1 npu_inst_pe_1_0_6_U3 ( .A1(npu_inst_pe_1_0_6_n27), .A2(
        npu_inst_pe_1_0_6_n1), .ZN(npu_inst_pe_1_0_6_n77) );
  FA_X1 npu_inst_pe_1_0_6_sub_77_U2_1 ( .A(int_o_data_npu[9]), .B(
        npu_inst_pe_1_0_6_n13), .CI(npu_inst_pe_1_0_6_sub_77_carry_1_), .CO(
        npu_inst_pe_1_0_6_sub_77_carry_2_), .S(npu_inst_pe_1_0_6_N66) );
  FA_X1 npu_inst_pe_1_0_6_add_79_U1_1 ( .A(int_o_data_npu[9]), .B(
        npu_inst_pe_1_0_6_int_data_1_), .CI(npu_inst_pe_1_0_6_add_79_carry_1_), 
        .CO(npu_inst_pe_1_0_6_add_79_carry_2_), .S(npu_inst_pe_1_0_6_N74) );
  NAND3_X1 npu_inst_pe_1_0_6_U101 ( .A1(npu_inst_pe_1_0_6_n4), .A2(
        npu_inst_pe_1_0_6_n6), .A3(npu_inst_pe_1_0_6_n7), .ZN(
        npu_inst_pe_1_0_6_n44) );
  NAND3_X1 npu_inst_pe_1_0_6_U100 ( .A1(npu_inst_pe_1_0_6_n3), .A2(
        npu_inst_pe_1_0_6_n6), .A3(npu_inst_pe_1_0_6_n7), .ZN(
        npu_inst_pe_1_0_6_n40) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_6_n33), .CK(
        npu_inst_pe_1_0_6_net4340), .RN(npu_inst_pe_1_0_6_n8), .Q(
        int_o_data_npu[14]) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_6_n34), .CK(
        npu_inst_pe_1_0_6_net4340), .RN(npu_inst_pe_1_0_6_n8), .Q(
        int_o_data_npu[13]) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_6_n35), .CK(
        npu_inst_pe_1_0_6_net4340), .RN(npu_inst_pe_1_0_6_n8), .Q(
        int_o_data_npu[12]) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_6_n36), .CK(
        npu_inst_pe_1_0_6_net4340), .RN(npu_inst_pe_1_0_6_n8), .Q(
        int_o_data_npu[11]) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_6_n98), .CK(
        npu_inst_pe_1_0_6_net4340), .RN(npu_inst_pe_1_0_6_n8), .Q(
        int_o_data_npu[10]) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_6_n99), .CK(
        npu_inst_pe_1_0_6_net4340), .RN(npu_inst_pe_1_0_6_n8), .Q(
        int_o_data_npu[9]) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_6_n32), .CK(
        npu_inst_pe_1_0_6_net4340), .RN(npu_inst_pe_1_0_6_n8), .Q(
        int_o_data_npu[15]) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_6_n100), 
        .CK(npu_inst_pe_1_0_6_net4340), .RN(npu_inst_pe_1_0_6_n8), .Q(
        int_o_data_npu[8]) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_weight_reg_0_ ( .D(npu_inst_n94), .CK(
        npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n8), .Q(
        npu_inst_pe_1_0_6_int_q_weight_0_), .QN(npu_inst_pe_1_0_6_n27) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_weight_reg_1_ ( .D(npu_inst_n100), .CK(
        npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n8), .Q(
        npu_inst_pe_1_0_6_int_q_weight_1_), .QN(npu_inst_pe_1_0_6_n26) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_6_n112), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n8), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_6_n106), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n8), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_6_n111), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_6_n105), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_6_n110), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_6_n104), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_6_n109), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_6_n103), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_6_n108), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_6_n102), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_6_n107), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_6_n101), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_6_n86), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_6_n87), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n9), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_6_n88), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_6_n89), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_6_n90), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_6_n91), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_6_n92), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_6_n93), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_6_n94), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_6_n95), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_6_n96), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_6_n97), 
        .CK(npu_inst_pe_1_0_6_net4346), .RN(npu_inst_pe_1_0_6_n10), .Q(
        npu_inst_pe_1_0_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_6_net4340) );
  CLKGATETST_X1 npu_inst_pe_1_0_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n48), .SE(1'b0), .GCK(npu_inst_pe_1_0_6_net4346) );
  MUX2_X1 npu_inst_pe_1_0_7_U153 ( .A(npu_inst_pe_1_0_7_n31), .B(
        npu_inst_pe_1_0_7_n28), .S(npu_inst_pe_1_0_7_n7), .Z(
        npu_inst_pe_1_0_7_N93) );
  MUX2_X1 npu_inst_pe_1_0_7_U152 ( .A(npu_inst_pe_1_0_7_n30), .B(
        npu_inst_pe_1_0_7_n29), .S(npu_inst_pe_1_0_7_n5), .Z(
        npu_inst_pe_1_0_7_n31) );
  MUX2_X1 npu_inst_pe_1_0_7_U151 ( .A(npu_inst_pe_1_0_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_0_7_n3), .Z(
        npu_inst_pe_1_0_7_n30) );
  MUX2_X1 npu_inst_pe_1_0_7_U150 ( .A(npu_inst_pe_1_0_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_0_7_n3), .Z(
        npu_inst_pe_1_0_7_n29) );
  MUX2_X1 npu_inst_pe_1_0_7_U149 ( .A(npu_inst_pe_1_0_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_0_7_n3), .Z(
        npu_inst_pe_1_0_7_n28) );
  MUX2_X1 npu_inst_pe_1_0_7_U148 ( .A(npu_inst_pe_1_0_7_n25), .B(
        npu_inst_pe_1_0_7_n22), .S(npu_inst_pe_1_0_7_n7), .Z(
        npu_inst_pe_1_0_7_N94) );
  MUX2_X1 npu_inst_pe_1_0_7_U147 ( .A(npu_inst_pe_1_0_7_n24), .B(
        npu_inst_pe_1_0_7_n23), .S(npu_inst_pe_1_0_7_n5), .Z(
        npu_inst_pe_1_0_7_n25) );
  MUX2_X1 npu_inst_pe_1_0_7_U146 ( .A(npu_inst_pe_1_0_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_0_7_n3), .Z(
        npu_inst_pe_1_0_7_n24) );
  MUX2_X1 npu_inst_pe_1_0_7_U145 ( .A(npu_inst_pe_1_0_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_0_7_n3), .Z(
        npu_inst_pe_1_0_7_n23) );
  MUX2_X1 npu_inst_pe_1_0_7_U144 ( .A(npu_inst_pe_1_0_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_0_7_n3), .Z(
        npu_inst_pe_1_0_7_n22) );
  MUX2_X1 npu_inst_pe_1_0_7_U143 ( .A(npu_inst_pe_1_0_7_n21), .B(
        npu_inst_pe_1_0_7_n18), .S(npu_inst_pe_1_0_7_n7), .Z(
        npu_inst_int_data_x_0__7__1_) );
  MUX2_X1 npu_inst_pe_1_0_7_U142 ( .A(npu_inst_pe_1_0_7_n20), .B(
        npu_inst_pe_1_0_7_n19), .S(npu_inst_pe_1_0_7_n5), .Z(
        npu_inst_pe_1_0_7_n21) );
  MUX2_X1 npu_inst_pe_1_0_7_U141 ( .A(npu_inst_pe_1_0_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_0_7_n3), .Z(
        npu_inst_pe_1_0_7_n20) );
  MUX2_X1 npu_inst_pe_1_0_7_U140 ( .A(npu_inst_pe_1_0_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_0_7_n3), .Z(
        npu_inst_pe_1_0_7_n19) );
  MUX2_X1 npu_inst_pe_1_0_7_U139 ( .A(npu_inst_pe_1_0_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_0_7_n3), .Z(
        npu_inst_pe_1_0_7_n18) );
  MUX2_X1 npu_inst_pe_1_0_7_U138 ( .A(npu_inst_pe_1_0_7_n17), .B(
        npu_inst_pe_1_0_7_n14), .S(npu_inst_pe_1_0_7_n7), .Z(
        npu_inst_int_data_x_0__7__0_) );
  MUX2_X1 npu_inst_pe_1_0_7_U137 ( .A(npu_inst_pe_1_0_7_n16), .B(
        npu_inst_pe_1_0_7_n15), .S(npu_inst_pe_1_0_7_n5), .Z(
        npu_inst_pe_1_0_7_n17) );
  MUX2_X1 npu_inst_pe_1_0_7_U136 ( .A(npu_inst_pe_1_0_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_0_7_n3), .Z(
        npu_inst_pe_1_0_7_n16) );
  MUX2_X1 npu_inst_pe_1_0_7_U135 ( .A(npu_inst_pe_1_0_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_0_7_n3), .Z(
        npu_inst_pe_1_0_7_n15) );
  MUX2_X1 npu_inst_pe_1_0_7_U134 ( .A(npu_inst_pe_1_0_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_0_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_0_7_n3), .Z(
        npu_inst_pe_1_0_7_n14) );
  XOR2_X1 npu_inst_pe_1_0_7_U133 ( .A(npu_inst_pe_1_0_7_int_data_0_), .B(
        int_o_data_npu[0]), .Z(npu_inst_pe_1_0_7_N73) );
  AND2_X1 npu_inst_pe_1_0_7_U132 ( .A1(int_o_data_npu[0]), .A2(
        npu_inst_pe_1_0_7_int_data_0_), .ZN(npu_inst_pe_1_0_7_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_0_7_U131 ( .A(int_o_data_npu[0]), .B(
        npu_inst_pe_1_0_7_n12), .ZN(npu_inst_pe_1_0_7_N65) );
  OR2_X1 npu_inst_pe_1_0_7_U130 ( .A1(npu_inst_pe_1_0_7_n12), .A2(
        int_o_data_npu[0]), .ZN(npu_inst_pe_1_0_7_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_0_7_U129 ( .A(int_o_data_npu[2]), .B(
        npu_inst_pe_1_0_7_add_79_carry_2_), .Z(npu_inst_pe_1_0_7_N75) );
  AND2_X1 npu_inst_pe_1_0_7_U128 ( .A1(npu_inst_pe_1_0_7_add_79_carry_2_), 
        .A2(int_o_data_npu[2]), .ZN(npu_inst_pe_1_0_7_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_0_7_U127 ( .A(int_o_data_npu[3]), .B(
        npu_inst_pe_1_0_7_add_79_carry_3_), .Z(npu_inst_pe_1_0_7_N76) );
  AND2_X1 npu_inst_pe_1_0_7_U126 ( .A1(npu_inst_pe_1_0_7_add_79_carry_3_), 
        .A2(int_o_data_npu[3]), .ZN(npu_inst_pe_1_0_7_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_0_7_U125 ( .A(int_o_data_npu[4]), .B(
        npu_inst_pe_1_0_7_add_79_carry_4_), .Z(npu_inst_pe_1_0_7_N77) );
  AND2_X1 npu_inst_pe_1_0_7_U124 ( .A1(npu_inst_pe_1_0_7_add_79_carry_4_), 
        .A2(int_o_data_npu[4]), .ZN(npu_inst_pe_1_0_7_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_0_7_U123 ( .A(int_o_data_npu[5]), .B(
        npu_inst_pe_1_0_7_add_79_carry_5_), .Z(npu_inst_pe_1_0_7_N78) );
  AND2_X1 npu_inst_pe_1_0_7_U122 ( .A1(npu_inst_pe_1_0_7_add_79_carry_5_), 
        .A2(int_o_data_npu[5]), .ZN(npu_inst_pe_1_0_7_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_0_7_U121 ( .A(int_o_data_npu[6]), .B(
        npu_inst_pe_1_0_7_add_79_carry_6_), .Z(npu_inst_pe_1_0_7_N79) );
  AND2_X1 npu_inst_pe_1_0_7_U120 ( .A1(npu_inst_pe_1_0_7_add_79_carry_6_), 
        .A2(int_o_data_npu[6]), .ZN(npu_inst_pe_1_0_7_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_0_7_U119 ( .A(int_o_data_npu[7]), .B(
        npu_inst_pe_1_0_7_add_79_carry_7_), .Z(npu_inst_pe_1_0_7_N80) );
  XNOR2_X1 npu_inst_pe_1_0_7_U118 ( .A(npu_inst_pe_1_0_7_sub_77_carry_2_), .B(
        int_o_data_npu[2]), .ZN(npu_inst_pe_1_0_7_N67) );
  OR2_X1 npu_inst_pe_1_0_7_U117 ( .A1(int_o_data_npu[2]), .A2(
        npu_inst_pe_1_0_7_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_0_7_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_0_7_U116 ( .A(npu_inst_pe_1_0_7_sub_77_carry_3_), .B(
        int_o_data_npu[3]), .ZN(npu_inst_pe_1_0_7_N68) );
  OR2_X1 npu_inst_pe_1_0_7_U115 ( .A1(int_o_data_npu[3]), .A2(
        npu_inst_pe_1_0_7_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_0_7_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_0_7_U114 ( .A(npu_inst_pe_1_0_7_sub_77_carry_4_), .B(
        int_o_data_npu[4]), .ZN(npu_inst_pe_1_0_7_N69) );
  OR2_X1 npu_inst_pe_1_0_7_U113 ( .A1(int_o_data_npu[4]), .A2(
        npu_inst_pe_1_0_7_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_0_7_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_0_7_U112 ( .A(npu_inst_pe_1_0_7_sub_77_carry_5_), .B(
        int_o_data_npu[5]), .ZN(npu_inst_pe_1_0_7_N70) );
  OR2_X1 npu_inst_pe_1_0_7_U111 ( .A1(int_o_data_npu[5]), .A2(
        npu_inst_pe_1_0_7_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_0_7_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_0_7_U110 ( .A(npu_inst_pe_1_0_7_sub_77_carry_6_), .B(
        int_o_data_npu[6]), .ZN(npu_inst_pe_1_0_7_N71) );
  OR2_X1 npu_inst_pe_1_0_7_U109 ( .A1(int_o_data_npu[6]), .A2(
        npu_inst_pe_1_0_7_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_0_7_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_0_7_U108 ( .A(int_o_data_npu[7]), .B(
        npu_inst_pe_1_0_7_sub_77_carry_7_), .ZN(npu_inst_pe_1_0_7_N72) );
  INV_X1 npu_inst_pe_1_0_7_U107 ( .A(npu_inst_n61), .ZN(npu_inst_pe_1_0_7_n6)
         );
  INV_X1 npu_inst_pe_1_0_7_U106 ( .A(npu_inst_pe_1_0_7_n6), .ZN(
        npu_inst_pe_1_0_7_n5) );
  INV_X1 npu_inst_pe_1_0_7_U105 ( .A(npu_inst_n42), .ZN(npu_inst_pe_1_0_7_n2)
         );
  AOI22_X1 npu_inst_pe_1_0_7_U104 ( .A1(npu_inst_int_data_y_1__7__0_), .A2(
        npu_inst_pe_1_0_7_n58), .B1(npu_inst_pe_1_0_7_n118), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_0_7_n57) );
  INV_X1 npu_inst_pe_1_0_7_U103 ( .A(npu_inst_pe_1_0_7_n57), .ZN(
        npu_inst_pe_1_0_7_n107) );
  AOI22_X1 npu_inst_pe_1_0_7_U102 ( .A1(npu_inst_int_data_y_1__7__0_), .A2(
        npu_inst_pe_1_0_7_n54), .B1(npu_inst_pe_1_0_7_n117), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_0_7_n53) );
  INV_X1 npu_inst_pe_1_0_7_U99 ( .A(npu_inst_pe_1_0_7_n53), .ZN(
        npu_inst_pe_1_0_7_n108) );
  AOI22_X1 npu_inst_pe_1_0_7_U98 ( .A1(npu_inst_int_data_y_1__7__0_), .A2(
        npu_inst_pe_1_0_7_n50), .B1(npu_inst_pe_1_0_7_n116), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_0_7_n49) );
  INV_X1 npu_inst_pe_1_0_7_U97 ( .A(npu_inst_pe_1_0_7_n49), .ZN(
        npu_inst_pe_1_0_7_n109) );
  AOI22_X1 npu_inst_pe_1_0_7_U96 ( .A1(npu_inst_int_data_y_1__7__0_), .A2(
        npu_inst_pe_1_0_7_n46), .B1(npu_inst_pe_1_0_7_n115), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_0_7_n45) );
  INV_X1 npu_inst_pe_1_0_7_U95 ( .A(npu_inst_pe_1_0_7_n45), .ZN(
        npu_inst_pe_1_0_7_n110) );
  AOI22_X1 npu_inst_pe_1_0_7_U94 ( .A1(npu_inst_int_data_y_1__7__0_), .A2(
        npu_inst_pe_1_0_7_n42), .B1(npu_inst_pe_1_0_7_n114), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_0_7_n41) );
  INV_X1 npu_inst_pe_1_0_7_U93 ( .A(npu_inst_pe_1_0_7_n41), .ZN(
        npu_inst_pe_1_0_7_n111) );
  AOI22_X1 npu_inst_pe_1_0_7_U92 ( .A1(npu_inst_int_data_y_1__7__1_), .A2(
        npu_inst_pe_1_0_7_n58), .B1(npu_inst_pe_1_0_7_n118), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_0_7_n59) );
  INV_X1 npu_inst_pe_1_0_7_U91 ( .A(npu_inst_pe_1_0_7_n59), .ZN(
        npu_inst_pe_1_0_7_n101) );
  AOI22_X1 npu_inst_pe_1_0_7_U90 ( .A1(npu_inst_int_data_y_1__7__1_), .A2(
        npu_inst_pe_1_0_7_n54), .B1(npu_inst_pe_1_0_7_n117), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_0_7_n55) );
  INV_X1 npu_inst_pe_1_0_7_U89 ( .A(npu_inst_pe_1_0_7_n55), .ZN(
        npu_inst_pe_1_0_7_n102) );
  AOI22_X1 npu_inst_pe_1_0_7_U88 ( .A1(npu_inst_int_data_y_1__7__1_), .A2(
        npu_inst_pe_1_0_7_n50), .B1(npu_inst_pe_1_0_7_n116), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_0_7_n51) );
  INV_X1 npu_inst_pe_1_0_7_U87 ( .A(npu_inst_pe_1_0_7_n51), .ZN(
        npu_inst_pe_1_0_7_n103) );
  AOI22_X1 npu_inst_pe_1_0_7_U86 ( .A1(npu_inst_int_data_y_1__7__1_), .A2(
        npu_inst_pe_1_0_7_n46), .B1(npu_inst_pe_1_0_7_n115), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_0_7_n47) );
  INV_X1 npu_inst_pe_1_0_7_U85 ( .A(npu_inst_pe_1_0_7_n47), .ZN(
        npu_inst_pe_1_0_7_n104) );
  AOI22_X1 npu_inst_pe_1_0_7_U84 ( .A1(npu_inst_int_data_y_1__7__1_), .A2(
        npu_inst_pe_1_0_7_n42), .B1(npu_inst_pe_1_0_7_n114), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_0_7_n43) );
  INV_X1 npu_inst_pe_1_0_7_U83 ( .A(npu_inst_pe_1_0_7_n43), .ZN(
        npu_inst_pe_1_0_7_n105) );
  AOI22_X1 npu_inst_pe_1_0_7_U82 ( .A1(npu_inst_pe_1_0_7_n38), .A2(
        npu_inst_int_data_y_1__7__1_), .B1(npu_inst_pe_1_0_7_n113), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_0_7_n39) );
  INV_X1 npu_inst_pe_1_0_7_U81 ( .A(npu_inst_pe_1_0_7_n39), .ZN(
        npu_inst_pe_1_0_7_n106) );
  AOI22_X1 npu_inst_pe_1_0_7_U80 ( .A1(npu_inst_pe_1_0_7_n38), .A2(
        npu_inst_int_data_y_1__7__0_), .B1(npu_inst_pe_1_0_7_n113), .B2(
        npu_inst_pe_1_0_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_0_7_n37) );
  INV_X1 npu_inst_pe_1_0_7_U79 ( .A(npu_inst_pe_1_0_7_n37), .ZN(
        npu_inst_pe_1_0_7_n112) );
  AOI222_X1 npu_inst_pe_1_0_7_U78 ( .A1(npu_inst_int_data_res_1__7__0_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N73), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N65), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n84) );
  INV_X1 npu_inst_pe_1_0_7_U77 ( .A(npu_inst_pe_1_0_7_n84), .ZN(
        npu_inst_pe_1_0_7_n100) );
  AOI222_X1 npu_inst_pe_1_0_7_U76 ( .A1(npu_inst_pe_1_0_7_n1), .A2(
        npu_inst_int_data_res_1__7__7_), .B1(npu_inst_pe_1_0_7_N80), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N72), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n75) );
  INV_X1 npu_inst_pe_1_0_7_U75 ( .A(npu_inst_pe_1_0_7_n75), .ZN(
        npu_inst_pe_1_0_7_n32) );
  AOI222_X1 npu_inst_pe_1_0_7_U74 ( .A1(npu_inst_int_data_res_1__7__2_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N75), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N67), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n82) );
  INV_X1 npu_inst_pe_1_0_7_U73 ( .A(npu_inst_pe_1_0_7_n82), .ZN(
        npu_inst_pe_1_0_7_n98) );
  AOI222_X1 npu_inst_pe_1_0_7_U72 ( .A1(npu_inst_int_data_res_1__7__3_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N76), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N68), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n81) );
  INV_X1 npu_inst_pe_1_0_7_U71 ( .A(npu_inst_pe_1_0_7_n81), .ZN(
        npu_inst_pe_1_0_7_n36) );
  AOI222_X1 npu_inst_pe_1_0_7_U70 ( .A1(npu_inst_int_data_res_1__7__4_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N77), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N69), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n80) );
  INV_X1 npu_inst_pe_1_0_7_U69 ( .A(npu_inst_pe_1_0_7_n80), .ZN(
        npu_inst_pe_1_0_7_n35) );
  AOI222_X1 npu_inst_pe_1_0_7_U68 ( .A1(npu_inst_int_data_res_1__7__5_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N78), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N70), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n79) );
  INV_X1 npu_inst_pe_1_0_7_U67 ( .A(npu_inst_pe_1_0_7_n79), .ZN(
        npu_inst_pe_1_0_7_n34) );
  AOI222_X1 npu_inst_pe_1_0_7_U66 ( .A1(npu_inst_int_data_res_1__7__6_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N79), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N71), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n78) );
  INV_X1 npu_inst_pe_1_0_7_U65 ( .A(npu_inst_pe_1_0_7_n78), .ZN(
        npu_inst_pe_1_0_7_n33) );
  NOR3_X1 npu_inst_pe_1_0_7_U64 ( .A1(npu_inst_pe_1_0_7_n26), .A2(npu_inst_n42), .A3(npu_inst_int_ckg[56]), .ZN(npu_inst_pe_1_0_7_n85) );
  OR2_X1 npu_inst_pe_1_0_7_U63 ( .A1(npu_inst_pe_1_0_7_n85), .A2(
        npu_inst_pe_1_0_7_n1), .ZN(npu_inst_pe_1_0_7_N84) );
  AND2_X1 npu_inst_pe_1_0_7_U62 ( .A1(npu_inst_int_data_x_0__7__1_), .A2(
        npu_inst_pe_1_0_7_int_q_weight_1_), .ZN(npu_inst_pe_1_0_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_0_7_U61 ( .A1(npu_inst_int_data_x_0__7__0_), .A2(
        npu_inst_pe_1_0_7_int_q_weight_1_), .ZN(npu_inst_pe_1_0_7_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_0_7_U60 ( .A(npu_inst_pe_1_0_7_int_data_1_), .ZN(
        npu_inst_pe_1_0_7_n13) );
  NAND2_X1 npu_inst_pe_1_0_7_U59 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_0_7_n60), .ZN(npu_inst_pe_1_0_7_n74) );
  OAI21_X1 npu_inst_pe_1_0_7_U58 ( .B1(npu_inst_pe_1_0_7_n63), .B2(
        npu_inst_pe_1_0_7_n60), .A(npu_inst_pe_1_0_7_n74), .ZN(
        npu_inst_pe_1_0_7_n97) );
  NAND2_X1 npu_inst_pe_1_0_7_U57 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_0_7_n60), .ZN(npu_inst_pe_1_0_7_n73) );
  OAI21_X1 npu_inst_pe_1_0_7_U56 ( .B1(npu_inst_pe_1_0_7_n61), .B2(
        npu_inst_pe_1_0_7_n60), .A(npu_inst_pe_1_0_7_n73), .ZN(
        npu_inst_pe_1_0_7_n96) );
  NAND2_X1 npu_inst_pe_1_0_7_U55 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_0_7_n56), .ZN(npu_inst_pe_1_0_7_n72) );
  OAI21_X1 npu_inst_pe_1_0_7_U54 ( .B1(npu_inst_pe_1_0_7_n63), .B2(
        npu_inst_pe_1_0_7_n56), .A(npu_inst_pe_1_0_7_n72), .ZN(
        npu_inst_pe_1_0_7_n95) );
  NAND2_X1 npu_inst_pe_1_0_7_U53 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_0_7_n56), .ZN(npu_inst_pe_1_0_7_n71) );
  OAI21_X1 npu_inst_pe_1_0_7_U52 ( .B1(npu_inst_pe_1_0_7_n61), .B2(
        npu_inst_pe_1_0_7_n56), .A(npu_inst_pe_1_0_7_n71), .ZN(
        npu_inst_pe_1_0_7_n94) );
  NAND2_X1 npu_inst_pe_1_0_7_U51 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_0_7_n52), .ZN(npu_inst_pe_1_0_7_n70) );
  OAI21_X1 npu_inst_pe_1_0_7_U50 ( .B1(npu_inst_pe_1_0_7_n63), .B2(
        npu_inst_pe_1_0_7_n52), .A(npu_inst_pe_1_0_7_n70), .ZN(
        npu_inst_pe_1_0_7_n93) );
  NAND2_X1 npu_inst_pe_1_0_7_U49 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_0_7_n52), .ZN(npu_inst_pe_1_0_7_n69) );
  OAI21_X1 npu_inst_pe_1_0_7_U48 ( .B1(npu_inst_pe_1_0_7_n61), .B2(
        npu_inst_pe_1_0_7_n52), .A(npu_inst_pe_1_0_7_n69), .ZN(
        npu_inst_pe_1_0_7_n92) );
  NAND2_X1 npu_inst_pe_1_0_7_U47 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_0_7_n48), .ZN(npu_inst_pe_1_0_7_n68) );
  OAI21_X1 npu_inst_pe_1_0_7_U46 ( .B1(npu_inst_pe_1_0_7_n63), .B2(
        npu_inst_pe_1_0_7_n48), .A(npu_inst_pe_1_0_7_n68), .ZN(
        npu_inst_pe_1_0_7_n91) );
  NAND2_X1 npu_inst_pe_1_0_7_U45 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_0_7_n48), .ZN(npu_inst_pe_1_0_7_n67) );
  OAI21_X1 npu_inst_pe_1_0_7_U44 ( .B1(npu_inst_pe_1_0_7_n61), .B2(
        npu_inst_pe_1_0_7_n48), .A(npu_inst_pe_1_0_7_n67), .ZN(
        npu_inst_pe_1_0_7_n90) );
  NAND2_X1 npu_inst_pe_1_0_7_U43 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_0_7_n44), .ZN(npu_inst_pe_1_0_7_n66) );
  OAI21_X1 npu_inst_pe_1_0_7_U42 ( .B1(npu_inst_pe_1_0_7_n63), .B2(
        npu_inst_pe_1_0_7_n44), .A(npu_inst_pe_1_0_7_n66), .ZN(
        npu_inst_pe_1_0_7_n89) );
  NAND2_X1 npu_inst_pe_1_0_7_U41 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_0_7_n44), .ZN(npu_inst_pe_1_0_7_n65) );
  OAI21_X1 npu_inst_pe_1_0_7_U40 ( .B1(npu_inst_pe_1_0_7_n61), .B2(
        npu_inst_pe_1_0_7_n44), .A(npu_inst_pe_1_0_7_n65), .ZN(
        npu_inst_pe_1_0_7_n88) );
  NAND2_X1 npu_inst_pe_1_0_7_U39 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_0_7_n40), .ZN(npu_inst_pe_1_0_7_n64) );
  OAI21_X1 npu_inst_pe_1_0_7_U38 ( .B1(npu_inst_pe_1_0_7_n63), .B2(
        npu_inst_pe_1_0_7_n40), .A(npu_inst_pe_1_0_7_n64), .ZN(
        npu_inst_pe_1_0_7_n87) );
  NAND2_X1 npu_inst_pe_1_0_7_U37 ( .A1(npu_inst_pe_1_0_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_0_7_n40), .ZN(npu_inst_pe_1_0_7_n62) );
  OAI21_X1 npu_inst_pe_1_0_7_U36 ( .B1(npu_inst_pe_1_0_7_n61), .B2(
        npu_inst_pe_1_0_7_n40), .A(npu_inst_pe_1_0_7_n62), .ZN(
        npu_inst_pe_1_0_7_n86) );
  AOI222_X1 npu_inst_pe_1_0_7_U35 ( .A1(npu_inst_int_data_res_1__7__1_), .A2(
        npu_inst_pe_1_0_7_n1), .B1(npu_inst_pe_1_0_7_N74), .B2(
        npu_inst_pe_1_0_7_n76), .C1(npu_inst_pe_1_0_7_N66), .C2(
        npu_inst_pe_1_0_7_n77), .ZN(npu_inst_pe_1_0_7_n83) );
  INV_X1 npu_inst_pe_1_0_7_U34 ( .A(npu_inst_pe_1_0_7_n83), .ZN(
        npu_inst_pe_1_0_7_n99) );
  AND2_X1 npu_inst_pe_1_0_7_U33 ( .A1(npu_inst_pe_1_0_7_N93), .A2(npu_inst_n42), .ZN(npu_inst_pe_1_0_7_o_data_v_0_) );
  AND2_X1 npu_inst_pe_1_0_7_U32 ( .A1(npu_inst_n42), .A2(npu_inst_pe_1_0_7_N94), .ZN(npu_inst_pe_1_0_7_o_data_v_1_) );
  INV_X1 npu_inst_pe_1_0_7_U31 ( .A(npu_inst_pe_1_0_7_int_data_0_), .ZN(
        npu_inst_pe_1_0_7_n12) );
  INV_X1 npu_inst_pe_1_0_7_U30 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_0_7_n4)
         );
  AOI22_X1 npu_inst_pe_1_0_7_U29 ( .A1(npu_inst_n42), .A2(
        npu_inst_int_data_y_1__7__1_), .B1(npu_inst_pe_1_0_7_n2), .B2(
        int_i_data_h_npu[15]), .ZN(npu_inst_pe_1_0_7_n63) );
  AOI22_X1 npu_inst_pe_1_0_7_U28 ( .A1(npu_inst_n42), .A2(
        npu_inst_int_data_y_1__7__0_), .B1(npu_inst_pe_1_0_7_n2), .B2(
        int_i_data_h_npu[14]), .ZN(npu_inst_pe_1_0_7_n61) );
  OR3_X1 npu_inst_pe_1_0_7_U27 ( .A1(npu_inst_pe_1_0_7_n5), .A2(
        npu_inst_pe_1_0_7_n7), .A3(npu_inst_pe_1_0_7_n4), .ZN(
        npu_inst_pe_1_0_7_n56) );
  OR3_X1 npu_inst_pe_1_0_7_U26 ( .A1(npu_inst_pe_1_0_7_n4), .A2(
        npu_inst_pe_1_0_7_n7), .A3(npu_inst_pe_1_0_7_n6), .ZN(
        npu_inst_pe_1_0_7_n48) );
  INV_X1 npu_inst_pe_1_0_7_U25 ( .A(npu_inst_pe_1_0_7_n4), .ZN(
        npu_inst_pe_1_0_7_n3) );
  OR3_X1 npu_inst_pe_1_0_7_U24 ( .A1(npu_inst_pe_1_0_7_n3), .A2(
        npu_inst_pe_1_0_7_n7), .A3(npu_inst_pe_1_0_7_n6), .ZN(
        npu_inst_pe_1_0_7_n52) );
  OR3_X1 npu_inst_pe_1_0_7_U23 ( .A1(npu_inst_pe_1_0_7_n5), .A2(
        npu_inst_pe_1_0_7_n7), .A3(npu_inst_pe_1_0_7_n3), .ZN(
        npu_inst_pe_1_0_7_n60) );
  BUF_X1 npu_inst_pe_1_0_7_U22 ( .A(npu_inst_n29), .Z(npu_inst_pe_1_0_7_n1) );
  NOR2_X1 npu_inst_pe_1_0_7_U21 ( .A1(npu_inst_pe_1_0_7_n60), .A2(
        npu_inst_pe_1_0_7_n2), .ZN(npu_inst_pe_1_0_7_n58) );
  NOR2_X1 npu_inst_pe_1_0_7_U20 ( .A1(npu_inst_pe_1_0_7_n56), .A2(
        npu_inst_pe_1_0_7_n2), .ZN(npu_inst_pe_1_0_7_n54) );
  NOR2_X1 npu_inst_pe_1_0_7_U19 ( .A1(npu_inst_pe_1_0_7_n52), .A2(
        npu_inst_pe_1_0_7_n2), .ZN(npu_inst_pe_1_0_7_n50) );
  NOR2_X1 npu_inst_pe_1_0_7_U18 ( .A1(npu_inst_pe_1_0_7_n48), .A2(
        npu_inst_pe_1_0_7_n2), .ZN(npu_inst_pe_1_0_7_n46) );
  NOR2_X1 npu_inst_pe_1_0_7_U17 ( .A1(npu_inst_pe_1_0_7_n40), .A2(
        npu_inst_pe_1_0_7_n2), .ZN(npu_inst_pe_1_0_7_n38) );
  NOR2_X1 npu_inst_pe_1_0_7_U16 ( .A1(npu_inst_pe_1_0_7_n44), .A2(
        npu_inst_pe_1_0_7_n2), .ZN(npu_inst_pe_1_0_7_n42) );
  BUF_X1 npu_inst_pe_1_0_7_U15 ( .A(npu_inst_n88), .Z(npu_inst_pe_1_0_7_n7) );
  INV_X1 npu_inst_pe_1_0_7_U14 ( .A(npu_inst_n108), .ZN(npu_inst_pe_1_0_7_n11)
         );
  INV_X1 npu_inst_pe_1_0_7_U13 ( .A(npu_inst_pe_1_0_7_n38), .ZN(
        npu_inst_pe_1_0_7_n113) );
  INV_X1 npu_inst_pe_1_0_7_U12 ( .A(npu_inst_pe_1_0_7_n58), .ZN(
        npu_inst_pe_1_0_7_n118) );
  INV_X1 npu_inst_pe_1_0_7_U11 ( .A(npu_inst_pe_1_0_7_n54), .ZN(
        npu_inst_pe_1_0_7_n117) );
  INV_X1 npu_inst_pe_1_0_7_U10 ( .A(npu_inst_pe_1_0_7_n50), .ZN(
        npu_inst_pe_1_0_7_n116) );
  INV_X1 npu_inst_pe_1_0_7_U9 ( .A(npu_inst_pe_1_0_7_n46), .ZN(
        npu_inst_pe_1_0_7_n115) );
  INV_X1 npu_inst_pe_1_0_7_U8 ( .A(npu_inst_pe_1_0_7_n42), .ZN(
        npu_inst_pe_1_0_7_n114) );
  BUF_X1 npu_inst_pe_1_0_7_U7 ( .A(npu_inst_pe_1_0_7_n11), .Z(
        npu_inst_pe_1_0_7_n10) );
  BUF_X1 npu_inst_pe_1_0_7_U6 ( .A(npu_inst_pe_1_0_7_n11), .Z(
        npu_inst_pe_1_0_7_n9) );
  BUF_X1 npu_inst_pe_1_0_7_U5 ( .A(npu_inst_pe_1_0_7_n11), .Z(
        npu_inst_pe_1_0_7_n8) );
  NOR2_X1 npu_inst_pe_1_0_7_U4 ( .A1(npu_inst_pe_1_0_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_0_7_n1), .ZN(npu_inst_pe_1_0_7_n76) );
  NOR2_X1 npu_inst_pe_1_0_7_U3 ( .A1(npu_inst_pe_1_0_7_n27), .A2(
        npu_inst_pe_1_0_7_n1), .ZN(npu_inst_pe_1_0_7_n77) );
  FA_X1 npu_inst_pe_1_0_7_sub_77_U2_1 ( .A(int_o_data_npu[1]), .B(
        npu_inst_pe_1_0_7_n13), .CI(npu_inst_pe_1_0_7_sub_77_carry_1_), .CO(
        npu_inst_pe_1_0_7_sub_77_carry_2_), .S(npu_inst_pe_1_0_7_N66) );
  FA_X1 npu_inst_pe_1_0_7_add_79_U1_1 ( .A(int_o_data_npu[1]), .B(
        npu_inst_pe_1_0_7_int_data_1_), .CI(npu_inst_pe_1_0_7_add_79_carry_1_), 
        .CO(npu_inst_pe_1_0_7_add_79_carry_2_), .S(npu_inst_pe_1_0_7_N74) );
  NAND3_X1 npu_inst_pe_1_0_7_U101 ( .A1(npu_inst_pe_1_0_7_n4), .A2(
        npu_inst_pe_1_0_7_n6), .A3(npu_inst_pe_1_0_7_n7), .ZN(
        npu_inst_pe_1_0_7_n44) );
  NAND3_X1 npu_inst_pe_1_0_7_U100 ( .A1(npu_inst_pe_1_0_7_n3), .A2(
        npu_inst_pe_1_0_7_n6), .A3(npu_inst_pe_1_0_7_n7), .ZN(
        npu_inst_pe_1_0_7_n40) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_0_7_n33), .CK(
        npu_inst_pe_1_0_7_net4317), .RN(npu_inst_pe_1_0_7_n8), .Q(
        int_o_data_npu[6]) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_0_7_n34), .CK(
        npu_inst_pe_1_0_7_net4317), .RN(npu_inst_pe_1_0_7_n8), .Q(
        int_o_data_npu[5]) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_0_7_n35), .CK(
        npu_inst_pe_1_0_7_net4317), .RN(npu_inst_pe_1_0_7_n8), .Q(
        int_o_data_npu[4]) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_0_7_n36), .CK(
        npu_inst_pe_1_0_7_net4317), .RN(npu_inst_pe_1_0_7_n8), .Q(
        int_o_data_npu[3]) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_0_7_n98), .CK(
        npu_inst_pe_1_0_7_net4317), .RN(npu_inst_pe_1_0_7_n8), .Q(
        int_o_data_npu[2]) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_0_7_n99), .CK(
        npu_inst_pe_1_0_7_net4317), .RN(npu_inst_pe_1_0_7_n8), .Q(
        int_o_data_npu[1]) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_0_7_n32), .CK(
        npu_inst_pe_1_0_7_net4317), .RN(npu_inst_pe_1_0_7_n8), .Q(
        int_o_data_npu[7]) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_0_7_n100), 
        .CK(npu_inst_pe_1_0_7_net4317), .RN(npu_inst_pe_1_0_7_n8), .Q(
        int_o_data_npu[0]) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_weight_reg_0_ ( .D(npu_inst_n94), .CK(
        npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n8), .Q(
        npu_inst_pe_1_0_7_int_q_weight_0_), .QN(npu_inst_pe_1_0_7_n27) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_weight_reg_1_ ( .D(npu_inst_n100), .CK(
        npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n8), .Q(
        npu_inst_pe_1_0_7_int_q_weight_1_), .QN(npu_inst_pe_1_0_7_n26) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_0_7_n112), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n8), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_0_7_n106), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n8), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_0_7_n111), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_0_7_n105), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_0_7_n110), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_0_7_n104), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_0_7_n109), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_0_7_n103), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_0_7_n108), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_0_7_n102), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_0_7_n107), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_0_7_n101), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_0_7_n86), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_0_7_n87), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n9), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_0_7_n88), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_0_7_n89), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_0_7_n90), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_0_7_n91), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_0_7_n92), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_0_7_n93), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_0_7_n94), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_0_7_n95), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_0_7_n96), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_0_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_0_7_n97), 
        .CK(npu_inst_pe_1_0_7_net4323), .RN(npu_inst_pe_1_0_7_n10), .Q(
        npu_inst_pe_1_0_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_0_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_0_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_0_7_net4317) );
  CLKGATETST_X1 npu_inst_pe_1_0_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n48), .SE(1'b0), .GCK(npu_inst_pe_1_0_7_net4323) );
  MUX2_X1 npu_inst_pe_1_1_0_U153 ( .A(npu_inst_pe_1_1_0_n31), .B(
        npu_inst_pe_1_1_0_n28), .S(npu_inst_pe_1_1_0_n7), .Z(
        npu_inst_pe_1_1_0_N93) );
  MUX2_X1 npu_inst_pe_1_1_0_U152 ( .A(npu_inst_pe_1_1_0_n30), .B(
        npu_inst_pe_1_1_0_n29), .S(npu_inst_pe_1_1_0_n5), .Z(
        npu_inst_pe_1_1_0_n31) );
  MUX2_X1 npu_inst_pe_1_1_0_U151 ( .A(npu_inst_pe_1_1_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_0_n3), .Z(
        npu_inst_pe_1_1_0_n30) );
  MUX2_X1 npu_inst_pe_1_1_0_U150 ( .A(npu_inst_pe_1_1_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_0_n3), .Z(
        npu_inst_pe_1_1_0_n29) );
  MUX2_X1 npu_inst_pe_1_1_0_U149 ( .A(npu_inst_pe_1_1_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_0_n3), .Z(
        npu_inst_pe_1_1_0_n28) );
  MUX2_X1 npu_inst_pe_1_1_0_U148 ( .A(npu_inst_pe_1_1_0_n25), .B(
        npu_inst_pe_1_1_0_n22), .S(npu_inst_pe_1_1_0_n7), .Z(
        npu_inst_pe_1_1_0_N94) );
  MUX2_X1 npu_inst_pe_1_1_0_U147 ( .A(npu_inst_pe_1_1_0_n24), .B(
        npu_inst_pe_1_1_0_n23), .S(npu_inst_pe_1_1_0_n5), .Z(
        npu_inst_pe_1_1_0_n25) );
  MUX2_X1 npu_inst_pe_1_1_0_U146 ( .A(npu_inst_pe_1_1_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_0_n3), .Z(
        npu_inst_pe_1_1_0_n24) );
  MUX2_X1 npu_inst_pe_1_1_0_U145 ( .A(npu_inst_pe_1_1_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_0_n3), .Z(
        npu_inst_pe_1_1_0_n23) );
  MUX2_X1 npu_inst_pe_1_1_0_U144 ( .A(npu_inst_pe_1_1_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_0_n3), .Z(
        npu_inst_pe_1_1_0_n22) );
  MUX2_X1 npu_inst_pe_1_1_0_U143 ( .A(npu_inst_pe_1_1_0_n21), .B(
        npu_inst_pe_1_1_0_n18), .S(npu_inst_pe_1_1_0_n7), .Z(
        npu_inst_pe_1_1_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_1_0_U142 ( .A(npu_inst_pe_1_1_0_n20), .B(
        npu_inst_pe_1_1_0_n19), .S(npu_inst_pe_1_1_0_n5), .Z(
        npu_inst_pe_1_1_0_n21) );
  MUX2_X1 npu_inst_pe_1_1_0_U141 ( .A(npu_inst_pe_1_1_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_0_n3), .Z(
        npu_inst_pe_1_1_0_n20) );
  MUX2_X1 npu_inst_pe_1_1_0_U140 ( .A(npu_inst_pe_1_1_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_0_n3), .Z(
        npu_inst_pe_1_1_0_n19) );
  MUX2_X1 npu_inst_pe_1_1_0_U139 ( .A(npu_inst_pe_1_1_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_0_n3), .Z(
        npu_inst_pe_1_1_0_n18) );
  MUX2_X1 npu_inst_pe_1_1_0_U138 ( .A(npu_inst_pe_1_1_0_n17), .B(
        npu_inst_pe_1_1_0_n14), .S(npu_inst_pe_1_1_0_n7), .Z(
        npu_inst_pe_1_1_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_1_0_U137 ( .A(npu_inst_pe_1_1_0_n16), .B(
        npu_inst_pe_1_1_0_n15), .S(npu_inst_pe_1_1_0_n5), .Z(
        npu_inst_pe_1_1_0_n17) );
  MUX2_X1 npu_inst_pe_1_1_0_U136 ( .A(npu_inst_pe_1_1_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_0_n3), .Z(
        npu_inst_pe_1_1_0_n16) );
  MUX2_X1 npu_inst_pe_1_1_0_U135 ( .A(npu_inst_pe_1_1_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_0_n3), .Z(
        npu_inst_pe_1_1_0_n15) );
  MUX2_X1 npu_inst_pe_1_1_0_U134 ( .A(npu_inst_pe_1_1_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_0_n3), .Z(
        npu_inst_pe_1_1_0_n14) );
  XOR2_X1 npu_inst_pe_1_1_0_U133 ( .A(npu_inst_pe_1_1_0_int_data_0_), .B(
        npu_inst_int_data_res_1__0__0_), .Z(npu_inst_pe_1_1_0_N73) );
  AND2_X1 npu_inst_pe_1_1_0_U132 ( .A1(npu_inst_int_data_res_1__0__0_), .A2(
        npu_inst_pe_1_1_0_int_data_0_), .ZN(npu_inst_pe_1_1_0_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_0_U131 ( .A(npu_inst_int_data_res_1__0__0_), .B(
        npu_inst_pe_1_1_0_n12), .ZN(npu_inst_pe_1_1_0_N65) );
  OR2_X1 npu_inst_pe_1_1_0_U130 ( .A1(npu_inst_pe_1_1_0_n12), .A2(
        npu_inst_int_data_res_1__0__0_), .ZN(npu_inst_pe_1_1_0_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_0_U129 ( .A(npu_inst_int_data_res_1__0__2_), .B(
        npu_inst_pe_1_1_0_add_79_carry_2_), .Z(npu_inst_pe_1_1_0_N75) );
  AND2_X1 npu_inst_pe_1_1_0_U128 ( .A1(npu_inst_pe_1_1_0_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_1__0__2_), .ZN(
        npu_inst_pe_1_1_0_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_0_U127 ( .A(npu_inst_int_data_res_1__0__3_), .B(
        npu_inst_pe_1_1_0_add_79_carry_3_), .Z(npu_inst_pe_1_1_0_N76) );
  AND2_X1 npu_inst_pe_1_1_0_U126 ( .A1(npu_inst_pe_1_1_0_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_1__0__3_), .ZN(
        npu_inst_pe_1_1_0_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_0_U125 ( .A(npu_inst_int_data_res_1__0__4_), .B(
        npu_inst_pe_1_1_0_add_79_carry_4_), .Z(npu_inst_pe_1_1_0_N77) );
  AND2_X1 npu_inst_pe_1_1_0_U124 ( .A1(npu_inst_pe_1_1_0_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_1__0__4_), .ZN(
        npu_inst_pe_1_1_0_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_0_U123 ( .A(npu_inst_int_data_res_1__0__5_), .B(
        npu_inst_pe_1_1_0_add_79_carry_5_), .Z(npu_inst_pe_1_1_0_N78) );
  AND2_X1 npu_inst_pe_1_1_0_U122 ( .A1(npu_inst_pe_1_1_0_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_1__0__5_), .ZN(
        npu_inst_pe_1_1_0_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_0_U121 ( .A(npu_inst_int_data_res_1__0__6_), .B(
        npu_inst_pe_1_1_0_add_79_carry_6_), .Z(npu_inst_pe_1_1_0_N79) );
  AND2_X1 npu_inst_pe_1_1_0_U120 ( .A1(npu_inst_pe_1_1_0_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_1__0__6_), .ZN(
        npu_inst_pe_1_1_0_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_0_U119 ( .A(npu_inst_int_data_res_1__0__7_), .B(
        npu_inst_pe_1_1_0_add_79_carry_7_), .Z(npu_inst_pe_1_1_0_N80) );
  XNOR2_X1 npu_inst_pe_1_1_0_U118 ( .A(npu_inst_pe_1_1_0_sub_77_carry_2_), .B(
        npu_inst_int_data_res_1__0__2_), .ZN(npu_inst_pe_1_1_0_N67) );
  OR2_X1 npu_inst_pe_1_1_0_U117 ( .A1(npu_inst_int_data_res_1__0__2_), .A2(
        npu_inst_pe_1_1_0_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_1_0_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_0_U116 ( .A(npu_inst_pe_1_1_0_sub_77_carry_3_), .B(
        npu_inst_int_data_res_1__0__3_), .ZN(npu_inst_pe_1_1_0_N68) );
  OR2_X1 npu_inst_pe_1_1_0_U115 ( .A1(npu_inst_int_data_res_1__0__3_), .A2(
        npu_inst_pe_1_1_0_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_1_0_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_0_U114 ( .A(npu_inst_pe_1_1_0_sub_77_carry_4_), .B(
        npu_inst_int_data_res_1__0__4_), .ZN(npu_inst_pe_1_1_0_N69) );
  OR2_X1 npu_inst_pe_1_1_0_U113 ( .A1(npu_inst_int_data_res_1__0__4_), .A2(
        npu_inst_pe_1_1_0_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_1_0_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_0_U112 ( .A(npu_inst_pe_1_1_0_sub_77_carry_5_), .B(
        npu_inst_int_data_res_1__0__5_), .ZN(npu_inst_pe_1_1_0_N70) );
  OR2_X1 npu_inst_pe_1_1_0_U111 ( .A1(npu_inst_int_data_res_1__0__5_), .A2(
        npu_inst_pe_1_1_0_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_1_0_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_0_U110 ( .A(npu_inst_pe_1_1_0_sub_77_carry_6_), .B(
        npu_inst_int_data_res_1__0__6_), .ZN(npu_inst_pe_1_1_0_N71) );
  OR2_X1 npu_inst_pe_1_1_0_U109 ( .A1(npu_inst_int_data_res_1__0__6_), .A2(
        npu_inst_pe_1_1_0_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_1_0_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_0_U108 ( .A(npu_inst_int_data_res_1__0__7_), .B(
        npu_inst_pe_1_1_0_sub_77_carry_7_), .ZN(npu_inst_pe_1_1_0_N72) );
  INV_X1 npu_inst_pe_1_1_0_U107 ( .A(npu_inst_n61), .ZN(npu_inst_pe_1_1_0_n6)
         );
  INV_X1 npu_inst_pe_1_1_0_U106 ( .A(npu_inst_pe_1_1_0_n6), .ZN(
        npu_inst_pe_1_1_0_n5) );
  INV_X1 npu_inst_pe_1_1_0_U105 ( .A(npu_inst_n41), .ZN(npu_inst_pe_1_1_0_n2)
         );
  AOI22_X1 npu_inst_pe_1_1_0_U104 ( .A1(npu_inst_int_data_y_2__0__0_), .A2(
        npu_inst_pe_1_1_0_n58), .B1(npu_inst_pe_1_1_0_n118), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_0_n57) );
  INV_X1 npu_inst_pe_1_1_0_U103 ( .A(npu_inst_pe_1_1_0_n57), .ZN(
        npu_inst_pe_1_1_0_n107) );
  AOI22_X1 npu_inst_pe_1_1_0_U102 ( .A1(npu_inst_int_data_y_2__0__0_), .A2(
        npu_inst_pe_1_1_0_n54), .B1(npu_inst_pe_1_1_0_n117), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_0_n53) );
  INV_X1 npu_inst_pe_1_1_0_U99 ( .A(npu_inst_pe_1_1_0_n53), .ZN(
        npu_inst_pe_1_1_0_n108) );
  AOI22_X1 npu_inst_pe_1_1_0_U98 ( .A1(npu_inst_int_data_y_2__0__0_), .A2(
        npu_inst_pe_1_1_0_n50), .B1(npu_inst_pe_1_1_0_n116), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_0_n49) );
  INV_X1 npu_inst_pe_1_1_0_U97 ( .A(npu_inst_pe_1_1_0_n49), .ZN(
        npu_inst_pe_1_1_0_n109) );
  AOI22_X1 npu_inst_pe_1_1_0_U96 ( .A1(npu_inst_int_data_y_2__0__0_), .A2(
        npu_inst_pe_1_1_0_n46), .B1(npu_inst_pe_1_1_0_n115), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_0_n45) );
  INV_X1 npu_inst_pe_1_1_0_U95 ( .A(npu_inst_pe_1_1_0_n45), .ZN(
        npu_inst_pe_1_1_0_n110) );
  AOI22_X1 npu_inst_pe_1_1_0_U94 ( .A1(npu_inst_int_data_y_2__0__0_), .A2(
        npu_inst_pe_1_1_0_n42), .B1(npu_inst_pe_1_1_0_n114), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_0_n41) );
  INV_X1 npu_inst_pe_1_1_0_U93 ( .A(npu_inst_pe_1_1_0_n41), .ZN(
        npu_inst_pe_1_1_0_n111) );
  AOI22_X1 npu_inst_pe_1_1_0_U92 ( .A1(npu_inst_int_data_y_2__0__1_), .A2(
        npu_inst_pe_1_1_0_n58), .B1(npu_inst_pe_1_1_0_n118), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_0_n59) );
  INV_X1 npu_inst_pe_1_1_0_U91 ( .A(npu_inst_pe_1_1_0_n59), .ZN(
        npu_inst_pe_1_1_0_n101) );
  AOI22_X1 npu_inst_pe_1_1_0_U90 ( .A1(npu_inst_int_data_y_2__0__1_), .A2(
        npu_inst_pe_1_1_0_n54), .B1(npu_inst_pe_1_1_0_n117), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_0_n55) );
  INV_X1 npu_inst_pe_1_1_0_U89 ( .A(npu_inst_pe_1_1_0_n55), .ZN(
        npu_inst_pe_1_1_0_n102) );
  AOI22_X1 npu_inst_pe_1_1_0_U88 ( .A1(npu_inst_int_data_y_2__0__1_), .A2(
        npu_inst_pe_1_1_0_n50), .B1(npu_inst_pe_1_1_0_n116), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_0_n51) );
  INV_X1 npu_inst_pe_1_1_0_U87 ( .A(npu_inst_pe_1_1_0_n51), .ZN(
        npu_inst_pe_1_1_0_n103) );
  AOI22_X1 npu_inst_pe_1_1_0_U86 ( .A1(npu_inst_int_data_y_2__0__1_), .A2(
        npu_inst_pe_1_1_0_n46), .B1(npu_inst_pe_1_1_0_n115), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_0_n47) );
  INV_X1 npu_inst_pe_1_1_0_U85 ( .A(npu_inst_pe_1_1_0_n47), .ZN(
        npu_inst_pe_1_1_0_n104) );
  AOI22_X1 npu_inst_pe_1_1_0_U84 ( .A1(npu_inst_int_data_y_2__0__1_), .A2(
        npu_inst_pe_1_1_0_n42), .B1(npu_inst_pe_1_1_0_n114), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_0_n43) );
  INV_X1 npu_inst_pe_1_1_0_U83 ( .A(npu_inst_pe_1_1_0_n43), .ZN(
        npu_inst_pe_1_1_0_n105) );
  AOI22_X1 npu_inst_pe_1_1_0_U82 ( .A1(npu_inst_pe_1_1_0_n38), .A2(
        npu_inst_int_data_y_2__0__1_), .B1(npu_inst_pe_1_1_0_n113), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_0_n39) );
  INV_X1 npu_inst_pe_1_1_0_U81 ( .A(npu_inst_pe_1_1_0_n39), .ZN(
        npu_inst_pe_1_1_0_n106) );
  NAND2_X1 npu_inst_pe_1_1_0_U80 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_0_n60), .ZN(npu_inst_pe_1_1_0_n74) );
  OAI21_X1 npu_inst_pe_1_1_0_U79 ( .B1(npu_inst_pe_1_1_0_n63), .B2(
        npu_inst_pe_1_1_0_n60), .A(npu_inst_pe_1_1_0_n74), .ZN(
        npu_inst_pe_1_1_0_n97) );
  NAND2_X1 npu_inst_pe_1_1_0_U78 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_0_n60), .ZN(npu_inst_pe_1_1_0_n73) );
  OAI21_X1 npu_inst_pe_1_1_0_U77 ( .B1(npu_inst_pe_1_1_0_n61), .B2(
        npu_inst_pe_1_1_0_n60), .A(npu_inst_pe_1_1_0_n73), .ZN(
        npu_inst_pe_1_1_0_n96) );
  NAND2_X1 npu_inst_pe_1_1_0_U76 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_0_n56), .ZN(npu_inst_pe_1_1_0_n72) );
  OAI21_X1 npu_inst_pe_1_1_0_U75 ( .B1(npu_inst_pe_1_1_0_n63), .B2(
        npu_inst_pe_1_1_0_n56), .A(npu_inst_pe_1_1_0_n72), .ZN(
        npu_inst_pe_1_1_0_n95) );
  NAND2_X1 npu_inst_pe_1_1_0_U74 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_0_n56), .ZN(npu_inst_pe_1_1_0_n71) );
  OAI21_X1 npu_inst_pe_1_1_0_U73 ( .B1(npu_inst_pe_1_1_0_n61), .B2(
        npu_inst_pe_1_1_0_n56), .A(npu_inst_pe_1_1_0_n71), .ZN(
        npu_inst_pe_1_1_0_n94) );
  NAND2_X1 npu_inst_pe_1_1_0_U72 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_0_n52), .ZN(npu_inst_pe_1_1_0_n70) );
  OAI21_X1 npu_inst_pe_1_1_0_U71 ( .B1(npu_inst_pe_1_1_0_n63), .B2(
        npu_inst_pe_1_1_0_n52), .A(npu_inst_pe_1_1_0_n70), .ZN(
        npu_inst_pe_1_1_0_n93) );
  NAND2_X1 npu_inst_pe_1_1_0_U70 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_0_n52), .ZN(npu_inst_pe_1_1_0_n69) );
  OAI21_X1 npu_inst_pe_1_1_0_U69 ( .B1(npu_inst_pe_1_1_0_n61), .B2(
        npu_inst_pe_1_1_0_n52), .A(npu_inst_pe_1_1_0_n69), .ZN(
        npu_inst_pe_1_1_0_n92) );
  NAND2_X1 npu_inst_pe_1_1_0_U68 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_0_n48), .ZN(npu_inst_pe_1_1_0_n68) );
  OAI21_X1 npu_inst_pe_1_1_0_U67 ( .B1(npu_inst_pe_1_1_0_n63), .B2(
        npu_inst_pe_1_1_0_n48), .A(npu_inst_pe_1_1_0_n68), .ZN(
        npu_inst_pe_1_1_0_n91) );
  NAND2_X1 npu_inst_pe_1_1_0_U66 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_0_n48), .ZN(npu_inst_pe_1_1_0_n67) );
  OAI21_X1 npu_inst_pe_1_1_0_U65 ( .B1(npu_inst_pe_1_1_0_n61), .B2(
        npu_inst_pe_1_1_0_n48), .A(npu_inst_pe_1_1_0_n67), .ZN(
        npu_inst_pe_1_1_0_n90) );
  NAND2_X1 npu_inst_pe_1_1_0_U64 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_0_n44), .ZN(npu_inst_pe_1_1_0_n66) );
  OAI21_X1 npu_inst_pe_1_1_0_U63 ( .B1(npu_inst_pe_1_1_0_n63), .B2(
        npu_inst_pe_1_1_0_n44), .A(npu_inst_pe_1_1_0_n66), .ZN(
        npu_inst_pe_1_1_0_n89) );
  NAND2_X1 npu_inst_pe_1_1_0_U62 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_0_n44), .ZN(npu_inst_pe_1_1_0_n65) );
  OAI21_X1 npu_inst_pe_1_1_0_U61 ( .B1(npu_inst_pe_1_1_0_n61), .B2(
        npu_inst_pe_1_1_0_n44), .A(npu_inst_pe_1_1_0_n65), .ZN(
        npu_inst_pe_1_1_0_n88) );
  NAND2_X1 npu_inst_pe_1_1_0_U60 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_0_n40), .ZN(npu_inst_pe_1_1_0_n64) );
  OAI21_X1 npu_inst_pe_1_1_0_U59 ( .B1(npu_inst_pe_1_1_0_n63), .B2(
        npu_inst_pe_1_1_0_n40), .A(npu_inst_pe_1_1_0_n64), .ZN(
        npu_inst_pe_1_1_0_n87) );
  NAND2_X1 npu_inst_pe_1_1_0_U58 ( .A1(npu_inst_pe_1_1_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_0_n40), .ZN(npu_inst_pe_1_1_0_n62) );
  OAI21_X1 npu_inst_pe_1_1_0_U57 ( .B1(npu_inst_pe_1_1_0_n61), .B2(
        npu_inst_pe_1_1_0_n40), .A(npu_inst_pe_1_1_0_n62), .ZN(
        npu_inst_pe_1_1_0_n86) );
  AOI22_X1 npu_inst_pe_1_1_0_U56 ( .A1(npu_inst_pe_1_1_0_n38), .A2(
        npu_inst_int_data_y_2__0__0_), .B1(npu_inst_pe_1_1_0_n113), .B2(
        npu_inst_pe_1_1_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_0_n37) );
  INV_X1 npu_inst_pe_1_1_0_U55 ( .A(npu_inst_pe_1_1_0_n37), .ZN(
        npu_inst_pe_1_1_0_n112) );
  AND2_X1 npu_inst_pe_1_1_0_U54 ( .A1(npu_inst_pe_1_1_0_N93), .A2(npu_inst_n41), .ZN(npu_inst_int_data_y_1__0__0_) );
  AND2_X1 npu_inst_pe_1_1_0_U53 ( .A1(npu_inst_n41), .A2(npu_inst_pe_1_1_0_N94), .ZN(npu_inst_int_data_y_1__0__1_) );
  AOI222_X1 npu_inst_pe_1_1_0_U52 ( .A1(npu_inst_int_data_res_2__0__0_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N73), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N65), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n84) );
  INV_X1 npu_inst_pe_1_1_0_U51 ( .A(npu_inst_pe_1_1_0_n84), .ZN(
        npu_inst_pe_1_1_0_n100) );
  AOI222_X1 npu_inst_pe_1_1_0_U50 ( .A1(npu_inst_pe_1_1_0_n1), .A2(
        npu_inst_int_data_res_2__0__7_), .B1(npu_inst_pe_1_1_0_N80), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N72), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n75) );
  INV_X1 npu_inst_pe_1_1_0_U49 ( .A(npu_inst_pe_1_1_0_n75), .ZN(
        npu_inst_pe_1_1_0_n32) );
  AOI222_X1 npu_inst_pe_1_1_0_U48 ( .A1(npu_inst_int_data_res_2__0__1_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N74), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N66), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n83) );
  INV_X1 npu_inst_pe_1_1_0_U47 ( .A(npu_inst_pe_1_1_0_n83), .ZN(
        npu_inst_pe_1_1_0_n99) );
  AOI222_X1 npu_inst_pe_1_1_0_U46 ( .A1(npu_inst_int_data_res_2__0__3_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N76), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N68), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n81) );
  INV_X1 npu_inst_pe_1_1_0_U45 ( .A(npu_inst_pe_1_1_0_n81), .ZN(
        npu_inst_pe_1_1_0_n36) );
  AOI222_X1 npu_inst_pe_1_1_0_U44 ( .A1(npu_inst_int_data_res_2__0__4_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N77), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N69), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n80) );
  INV_X1 npu_inst_pe_1_1_0_U43 ( .A(npu_inst_pe_1_1_0_n80), .ZN(
        npu_inst_pe_1_1_0_n35) );
  AOI222_X1 npu_inst_pe_1_1_0_U42 ( .A1(npu_inst_int_data_res_2__0__5_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N78), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N70), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n79) );
  INV_X1 npu_inst_pe_1_1_0_U41 ( .A(npu_inst_pe_1_1_0_n79), .ZN(
        npu_inst_pe_1_1_0_n34) );
  AOI222_X1 npu_inst_pe_1_1_0_U40 ( .A1(npu_inst_int_data_res_2__0__6_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N79), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N71), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n78) );
  INV_X1 npu_inst_pe_1_1_0_U39 ( .A(npu_inst_pe_1_1_0_n78), .ZN(
        npu_inst_pe_1_1_0_n33) );
  AND2_X1 npu_inst_pe_1_1_0_U38 ( .A1(npu_inst_pe_1_1_0_o_data_h_1_), .A2(
        npu_inst_pe_1_1_0_int_q_weight_1_), .ZN(npu_inst_pe_1_1_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_0_U37 ( .A1(npu_inst_pe_1_1_0_o_data_h_0_), .A2(
        npu_inst_pe_1_1_0_int_q_weight_1_), .ZN(npu_inst_pe_1_1_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_1_0_U36 ( .A(npu_inst_pe_1_1_0_int_data_1_), .ZN(
        npu_inst_pe_1_1_0_n13) );
  NOR3_X1 npu_inst_pe_1_1_0_U35 ( .A1(npu_inst_pe_1_1_0_n26), .A2(npu_inst_n41), .A3(npu_inst_int_ckg[55]), .ZN(npu_inst_pe_1_1_0_n85) );
  OR2_X1 npu_inst_pe_1_1_0_U34 ( .A1(npu_inst_pe_1_1_0_n85), .A2(
        npu_inst_pe_1_1_0_n1), .ZN(npu_inst_pe_1_1_0_N84) );
  AOI222_X1 npu_inst_pe_1_1_0_U33 ( .A1(npu_inst_int_data_res_2__0__2_), .A2(
        npu_inst_pe_1_1_0_n1), .B1(npu_inst_pe_1_1_0_N75), .B2(
        npu_inst_pe_1_1_0_n76), .C1(npu_inst_pe_1_1_0_N67), .C2(
        npu_inst_pe_1_1_0_n77), .ZN(npu_inst_pe_1_1_0_n82) );
  INV_X1 npu_inst_pe_1_1_0_U32 ( .A(npu_inst_pe_1_1_0_n82), .ZN(
        npu_inst_pe_1_1_0_n98) );
  AOI22_X1 npu_inst_pe_1_1_0_U31 ( .A1(npu_inst_n41), .A2(
        npu_inst_int_data_y_2__0__1_), .B1(npu_inst_pe_1_1_0_n2), .B2(
        npu_inst_int_data_x_1__1__1_), .ZN(npu_inst_pe_1_1_0_n63) );
  AOI22_X1 npu_inst_pe_1_1_0_U30 ( .A1(npu_inst_n41), .A2(
        npu_inst_int_data_y_2__0__0_), .B1(npu_inst_pe_1_1_0_n2), .B2(
        npu_inst_int_data_x_1__1__0_), .ZN(npu_inst_pe_1_1_0_n61) );
  INV_X1 npu_inst_pe_1_1_0_U29 ( .A(npu_inst_pe_1_1_0_int_data_0_), .ZN(
        npu_inst_pe_1_1_0_n12) );
  INV_X1 npu_inst_pe_1_1_0_U28 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_1_0_n4)
         );
  OR3_X1 npu_inst_pe_1_1_0_U27 ( .A1(npu_inst_pe_1_1_0_n5), .A2(
        npu_inst_pe_1_1_0_n7), .A3(npu_inst_pe_1_1_0_n4), .ZN(
        npu_inst_pe_1_1_0_n56) );
  OR3_X1 npu_inst_pe_1_1_0_U26 ( .A1(npu_inst_pe_1_1_0_n4), .A2(
        npu_inst_pe_1_1_0_n7), .A3(npu_inst_pe_1_1_0_n6), .ZN(
        npu_inst_pe_1_1_0_n48) );
  INV_X1 npu_inst_pe_1_1_0_U25 ( .A(npu_inst_pe_1_1_0_n4), .ZN(
        npu_inst_pe_1_1_0_n3) );
  OR3_X1 npu_inst_pe_1_1_0_U24 ( .A1(npu_inst_pe_1_1_0_n3), .A2(
        npu_inst_pe_1_1_0_n7), .A3(npu_inst_pe_1_1_0_n6), .ZN(
        npu_inst_pe_1_1_0_n52) );
  OR3_X1 npu_inst_pe_1_1_0_U23 ( .A1(npu_inst_pe_1_1_0_n5), .A2(
        npu_inst_pe_1_1_0_n7), .A3(npu_inst_pe_1_1_0_n3), .ZN(
        npu_inst_pe_1_1_0_n60) );
  BUF_X1 npu_inst_pe_1_1_0_U22 ( .A(npu_inst_n29), .Z(npu_inst_pe_1_1_0_n1) );
  NOR2_X1 npu_inst_pe_1_1_0_U21 ( .A1(npu_inst_pe_1_1_0_n60), .A2(
        npu_inst_pe_1_1_0_n2), .ZN(npu_inst_pe_1_1_0_n58) );
  NOR2_X1 npu_inst_pe_1_1_0_U20 ( .A1(npu_inst_pe_1_1_0_n56), .A2(
        npu_inst_pe_1_1_0_n2), .ZN(npu_inst_pe_1_1_0_n54) );
  NOR2_X1 npu_inst_pe_1_1_0_U19 ( .A1(npu_inst_pe_1_1_0_n52), .A2(
        npu_inst_pe_1_1_0_n2), .ZN(npu_inst_pe_1_1_0_n50) );
  NOR2_X1 npu_inst_pe_1_1_0_U18 ( .A1(npu_inst_pe_1_1_0_n48), .A2(
        npu_inst_pe_1_1_0_n2), .ZN(npu_inst_pe_1_1_0_n46) );
  NOR2_X1 npu_inst_pe_1_1_0_U17 ( .A1(npu_inst_pe_1_1_0_n40), .A2(
        npu_inst_pe_1_1_0_n2), .ZN(npu_inst_pe_1_1_0_n38) );
  NOR2_X1 npu_inst_pe_1_1_0_U16 ( .A1(npu_inst_pe_1_1_0_n44), .A2(
        npu_inst_pe_1_1_0_n2), .ZN(npu_inst_pe_1_1_0_n42) );
  BUF_X1 npu_inst_pe_1_1_0_U15 ( .A(npu_inst_n87), .Z(npu_inst_pe_1_1_0_n7) );
  INV_X1 npu_inst_pe_1_1_0_U14 ( .A(npu_inst_n108), .ZN(npu_inst_pe_1_1_0_n11)
         );
  INV_X1 npu_inst_pe_1_1_0_U13 ( .A(npu_inst_pe_1_1_0_n38), .ZN(
        npu_inst_pe_1_1_0_n113) );
  INV_X1 npu_inst_pe_1_1_0_U12 ( .A(npu_inst_pe_1_1_0_n58), .ZN(
        npu_inst_pe_1_1_0_n118) );
  INV_X1 npu_inst_pe_1_1_0_U11 ( .A(npu_inst_pe_1_1_0_n54), .ZN(
        npu_inst_pe_1_1_0_n117) );
  INV_X1 npu_inst_pe_1_1_0_U10 ( .A(npu_inst_pe_1_1_0_n50), .ZN(
        npu_inst_pe_1_1_0_n116) );
  INV_X1 npu_inst_pe_1_1_0_U9 ( .A(npu_inst_pe_1_1_0_n46), .ZN(
        npu_inst_pe_1_1_0_n115) );
  INV_X1 npu_inst_pe_1_1_0_U8 ( .A(npu_inst_pe_1_1_0_n42), .ZN(
        npu_inst_pe_1_1_0_n114) );
  BUF_X1 npu_inst_pe_1_1_0_U7 ( .A(npu_inst_pe_1_1_0_n11), .Z(
        npu_inst_pe_1_1_0_n10) );
  BUF_X1 npu_inst_pe_1_1_0_U6 ( .A(npu_inst_pe_1_1_0_n11), .Z(
        npu_inst_pe_1_1_0_n9) );
  BUF_X1 npu_inst_pe_1_1_0_U5 ( .A(npu_inst_pe_1_1_0_n11), .Z(
        npu_inst_pe_1_1_0_n8) );
  NOR2_X1 npu_inst_pe_1_1_0_U4 ( .A1(npu_inst_pe_1_1_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_0_n1), .ZN(npu_inst_pe_1_1_0_n76) );
  NOR2_X1 npu_inst_pe_1_1_0_U3 ( .A1(npu_inst_pe_1_1_0_n27), .A2(
        npu_inst_pe_1_1_0_n1), .ZN(npu_inst_pe_1_1_0_n77) );
  FA_X1 npu_inst_pe_1_1_0_sub_77_U2_1 ( .A(npu_inst_int_data_res_1__0__1_), 
        .B(npu_inst_pe_1_1_0_n13), .CI(npu_inst_pe_1_1_0_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_1_0_sub_77_carry_2_), .S(npu_inst_pe_1_1_0_N66) );
  FA_X1 npu_inst_pe_1_1_0_add_79_U1_1 ( .A(npu_inst_int_data_res_1__0__1_), 
        .B(npu_inst_pe_1_1_0_int_data_1_), .CI(
        npu_inst_pe_1_1_0_add_79_carry_1_), .CO(
        npu_inst_pe_1_1_0_add_79_carry_2_), .S(npu_inst_pe_1_1_0_N74) );
  NAND3_X1 npu_inst_pe_1_1_0_U101 ( .A1(npu_inst_pe_1_1_0_n4), .A2(
        npu_inst_pe_1_1_0_n6), .A3(npu_inst_pe_1_1_0_n7), .ZN(
        npu_inst_pe_1_1_0_n44) );
  NAND3_X1 npu_inst_pe_1_1_0_U100 ( .A1(npu_inst_pe_1_1_0_n3), .A2(
        npu_inst_pe_1_1_0_n6), .A3(npu_inst_pe_1_1_0_n7), .ZN(
        npu_inst_pe_1_1_0_n40) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_0_n33), .CK(
        npu_inst_pe_1_1_0_net4294), .RN(npu_inst_pe_1_1_0_n8), .Q(
        npu_inst_int_data_res_1__0__6_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_0_n34), .CK(
        npu_inst_pe_1_1_0_net4294), .RN(npu_inst_pe_1_1_0_n8), .Q(
        npu_inst_int_data_res_1__0__5_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_0_n35), .CK(
        npu_inst_pe_1_1_0_net4294), .RN(npu_inst_pe_1_1_0_n8), .Q(
        npu_inst_int_data_res_1__0__4_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_0_n36), .CK(
        npu_inst_pe_1_1_0_net4294), .RN(npu_inst_pe_1_1_0_n8), .Q(
        npu_inst_int_data_res_1__0__3_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_0_n98), .CK(
        npu_inst_pe_1_1_0_net4294), .RN(npu_inst_pe_1_1_0_n8), .Q(
        npu_inst_int_data_res_1__0__2_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_0_n99), .CK(
        npu_inst_pe_1_1_0_net4294), .RN(npu_inst_pe_1_1_0_n8), .Q(
        npu_inst_int_data_res_1__0__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_0_n32), .CK(
        npu_inst_pe_1_1_0_net4294), .RN(npu_inst_pe_1_1_0_n8), .Q(
        npu_inst_int_data_res_1__0__7_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_0_n100), 
        .CK(npu_inst_pe_1_1_0_net4294), .RN(npu_inst_pe_1_1_0_n8), .Q(
        npu_inst_int_data_res_1__0__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_weight_reg_0_ ( .D(npu_inst_n94), .CK(
        npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n8), .Q(
        npu_inst_pe_1_1_0_int_q_weight_0_), .QN(npu_inst_pe_1_1_0_n27) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_weight_reg_1_ ( .D(npu_inst_n100), .CK(
        npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n8), .Q(
        npu_inst_pe_1_1_0_int_q_weight_1_), .QN(npu_inst_pe_1_1_0_n26) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_0_n112), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n8), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_0_n106), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n8), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_0_n111), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_0_n105), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_0_n110), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_0_n104), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_0_n109), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_0_n103), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_0_n108), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_0_n102), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_0_n107), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_0_n101), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_0_n86), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_0_n87), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n9), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_0_n88), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_0_n89), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_0_n90), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_0_n91), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_0_n92), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_0_n93), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_0_n94), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_0_n95), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_0_n96), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_0_n97), 
        .CK(npu_inst_pe_1_1_0_net4300), .RN(npu_inst_pe_1_1_0_n10), .Q(
        npu_inst_pe_1_1_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_0_net4294) );
  CLKGATETST_X1 npu_inst_pe_1_1_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n48), .SE(1'b0), .GCK(npu_inst_pe_1_1_0_net4300) );
  MUX2_X1 npu_inst_pe_1_1_1_U153 ( .A(npu_inst_pe_1_1_1_n31), .B(
        npu_inst_pe_1_1_1_n28), .S(npu_inst_pe_1_1_1_n7), .Z(
        npu_inst_pe_1_1_1_N93) );
  MUX2_X1 npu_inst_pe_1_1_1_U152 ( .A(npu_inst_pe_1_1_1_n30), .B(
        npu_inst_pe_1_1_1_n29), .S(npu_inst_pe_1_1_1_n5), .Z(
        npu_inst_pe_1_1_1_n31) );
  MUX2_X1 npu_inst_pe_1_1_1_U151 ( .A(npu_inst_pe_1_1_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_1_n3), .Z(
        npu_inst_pe_1_1_1_n30) );
  MUX2_X1 npu_inst_pe_1_1_1_U150 ( .A(npu_inst_pe_1_1_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_1_n3), .Z(
        npu_inst_pe_1_1_1_n29) );
  MUX2_X1 npu_inst_pe_1_1_1_U149 ( .A(npu_inst_pe_1_1_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_1_n3), .Z(
        npu_inst_pe_1_1_1_n28) );
  MUX2_X1 npu_inst_pe_1_1_1_U148 ( .A(npu_inst_pe_1_1_1_n25), .B(
        npu_inst_pe_1_1_1_n22), .S(npu_inst_pe_1_1_1_n7), .Z(
        npu_inst_pe_1_1_1_N94) );
  MUX2_X1 npu_inst_pe_1_1_1_U147 ( .A(npu_inst_pe_1_1_1_n24), .B(
        npu_inst_pe_1_1_1_n23), .S(npu_inst_pe_1_1_1_n5), .Z(
        npu_inst_pe_1_1_1_n25) );
  MUX2_X1 npu_inst_pe_1_1_1_U146 ( .A(npu_inst_pe_1_1_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_1_n3), .Z(
        npu_inst_pe_1_1_1_n24) );
  MUX2_X1 npu_inst_pe_1_1_1_U145 ( .A(npu_inst_pe_1_1_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_1_n3), .Z(
        npu_inst_pe_1_1_1_n23) );
  MUX2_X1 npu_inst_pe_1_1_1_U144 ( .A(npu_inst_pe_1_1_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_1_n3), .Z(
        npu_inst_pe_1_1_1_n22) );
  MUX2_X1 npu_inst_pe_1_1_1_U143 ( .A(npu_inst_pe_1_1_1_n21), .B(
        npu_inst_pe_1_1_1_n18), .S(npu_inst_pe_1_1_1_n7), .Z(
        npu_inst_int_data_x_1__1__1_) );
  MUX2_X1 npu_inst_pe_1_1_1_U142 ( .A(npu_inst_pe_1_1_1_n20), .B(
        npu_inst_pe_1_1_1_n19), .S(npu_inst_pe_1_1_1_n5), .Z(
        npu_inst_pe_1_1_1_n21) );
  MUX2_X1 npu_inst_pe_1_1_1_U141 ( .A(npu_inst_pe_1_1_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_1_n3), .Z(
        npu_inst_pe_1_1_1_n20) );
  MUX2_X1 npu_inst_pe_1_1_1_U140 ( .A(npu_inst_pe_1_1_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_1_n3), .Z(
        npu_inst_pe_1_1_1_n19) );
  MUX2_X1 npu_inst_pe_1_1_1_U139 ( .A(npu_inst_pe_1_1_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_1_n3), .Z(
        npu_inst_pe_1_1_1_n18) );
  MUX2_X1 npu_inst_pe_1_1_1_U138 ( .A(npu_inst_pe_1_1_1_n17), .B(
        npu_inst_pe_1_1_1_n14), .S(npu_inst_pe_1_1_1_n7), .Z(
        npu_inst_int_data_x_1__1__0_) );
  MUX2_X1 npu_inst_pe_1_1_1_U137 ( .A(npu_inst_pe_1_1_1_n16), .B(
        npu_inst_pe_1_1_1_n15), .S(npu_inst_pe_1_1_1_n5), .Z(
        npu_inst_pe_1_1_1_n17) );
  MUX2_X1 npu_inst_pe_1_1_1_U136 ( .A(npu_inst_pe_1_1_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_1_n3), .Z(
        npu_inst_pe_1_1_1_n16) );
  MUX2_X1 npu_inst_pe_1_1_1_U135 ( .A(npu_inst_pe_1_1_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_1_n3), .Z(
        npu_inst_pe_1_1_1_n15) );
  MUX2_X1 npu_inst_pe_1_1_1_U134 ( .A(npu_inst_pe_1_1_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_1_n3), .Z(
        npu_inst_pe_1_1_1_n14) );
  XOR2_X1 npu_inst_pe_1_1_1_U133 ( .A(npu_inst_pe_1_1_1_int_data_0_), .B(
        npu_inst_int_data_res_1__1__0_), .Z(npu_inst_pe_1_1_1_N73) );
  AND2_X1 npu_inst_pe_1_1_1_U132 ( .A1(npu_inst_int_data_res_1__1__0_), .A2(
        npu_inst_pe_1_1_1_int_data_0_), .ZN(npu_inst_pe_1_1_1_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_1_U131 ( .A(npu_inst_int_data_res_1__1__0_), .B(
        npu_inst_pe_1_1_1_n12), .ZN(npu_inst_pe_1_1_1_N65) );
  OR2_X1 npu_inst_pe_1_1_1_U130 ( .A1(npu_inst_pe_1_1_1_n12), .A2(
        npu_inst_int_data_res_1__1__0_), .ZN(npu_inst_pe_1_1_1_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_1_U129 ( .A(npu_inst_int_data_res_1__1__2_), .B(
        npu_inst_pe_1_1_1_add_79_carry_2_), .Z(npu_inst_pe_1_1_1_N75) );
  AND2_X1 npu_inst_pe_1_1_1_U128 ( .A1(npu_inst_pe_1_1_1_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_1__1__2_), .ZN(
        npu_inst_pe_1_1_1_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_1_U127 ( .A(npu_inst_int_data_res_1__1__3_), .B(
        npu_inst_pe_1_1_1_add_79_carry_3_), .Z(npu_inst_pe_1_1_1_N76) );
  AND2_X1 npu_inst_pe_1_1_1_U126 ( .A1(npu_inst_pe_1_1_1_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_1__1__3_), .ZN(
        npu_inst_pe_1_1_1_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_1_U125 ( .A(npu_inst_int_data_res_1__1__4_), .B(
        npu_inst_pe_1_1_1_add_79_carry_4_), .Z(npu_inst_pe_1_1_1_N77) );
  AND2_X1 npu_inst_pe_1_1_1_U124 ( .A1(npu_inst_pe_1_1_1_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_1__1__4_), .ZN(
        npu_inst_pe_1_1_1_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_1_U123 ( .A(npu_inst_int_data_res_1__1__5_), .B(
        npu_inst_pe_1_1_1_add_79_carry_5_), .Z(npu_inst_pe_1_1_1_N78) );
  AND2_X1 npu_inst_pe_1_1_1_U122 ( .A1(npu_inst_pe_1_1_1_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_1__1__5_), .ZN(
        npu_inst_pe_1_1_1_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_1_U121 ( .A(npu_inst_int_data_res_1__1__6_), .B(
        npu_inst_pe_1_1_1_add_79_carry_6_), .Z(npu_inst_pe_1_1_1_N79) );
  AND2_X1 npu_inst_pe_1_1_1_U120 ( .A1(npu_inst_pe_1_1_1_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_1__1__6_), .ZN(
        npu_inst_pe_1_1_1_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_1_U119 ( .A(npu_inst_int_data_res_1__1__7_), .B(
        npu_inst_pe_1_1_1_add_79_carry_7_), .Z(npu_inst_pe_1_1_1_N80) );
  XNOR2_X1 npu_inst_pe_1_1_1_U118 ( .A(npu_inst_pe_1_1_1_sub_77_carry_2_), .B(
        npu_inst_int_data_res_1__1__2_), .ZN(npu_inst_pe_1_1_1_N67) );
  OR2_X1 npu_inst_pe_1_1_1_U117 ( .A1(npu_inst_int_data_res_1__1__2_), .A2(
        npu_inst_pe_1_1_1_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_1_1_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_1_U116 ( .A(npu_inst_pe_1_1_1_sub_77_carry_3_), .B(
        npu_inst_int_data_res_1__1__3_), .ZN(npu_inst_pe_1_1_1_N68) );
  OR2_X1 npu_inst_pe_1_1_1_U115 ( .A1(npu_inst_int_data_res_1__1__3_), .A2(
        npu_inst_pe_1_1_1_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_1_1_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_1_U114 ( .A(npu_inst_pe_1_1_1_sub_77_carry_4_), .B(
        npu_inst_int_data_res_1__1__4_), .ZN(npu_inst_pe_1_1_1_N69) );
  OR2_X1 npu_inst_pe_1_1_1_U113 ( .A1(npu_inst_int_data_res_1__1__4_), .A2(
        npu_inst_pe_1_1_1_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_1_1_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_1_U112 ( .A(npu_inst_pe_1_1_1_sub_77_carry_5_), .B(
        npu_inst_int_data_res_1__1__5_), .ZN(npu_inst_pe_1_1_1_N70) );
  OR2_X1 npu_inst_pe_1_1_1_U111 ( .A1(npu_inst_int_data_res_1__1__5_), .A2(
        npu_inst_pe_1_1_1_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_1_1_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_1_U110 ( .A(npu_inst_pe_1_1_1_sub_77_carry_6_), .B(
        npu_inst_int_data_res_1__1__6_), .ZN(npu_inst_pe_1_1_1_N71) );
  OR2_X1 npu_inst_pe_1_1_1_U109 ( .A1(npu_inst_int_data_res_1__1__6_), .A2(
        npu_inst_pe_1_1_1_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_1_1_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_1_U108 ( .A(npu_inst_int_data_res_1__1__7_), .B(
        npu_inst_pe_1_1_1_sub_77_carry_7_), .ZN(npu_inst_pe_1_1_1_N72) );
  INV_X1 npu_inst_pe_1_1_1_U107 ( .A(npu_inst_n61), .ZN(npu_inst_pe_1_1_1_n6)
         );
  INV_X1 npu_inst_pe_1_1_1_U106 ( .A(npu_inst_pe_1_1_1_n6), .ZN(
        npu_inst_pe_1_1_1_n5) );
  INV_X1 npu_inst_pe_1_1_1_U105 ( .A(npu_inst_n41), .ZN(npu_inst_pe_1_1_1_n2)
         );
  AOI22_X1 npu_inst_pe_1_1_1_U104 ( .A1(npu_inst_int_data_y_2__1__0_), .A2(
        npu_inst_pe_1_1_1_n58), .B1(npu_inst_pe_1_1_1_n118), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_1_n57) );
  INV_X1 npu_inst_pe_1_1_1_U103 ( .A(npu_inst_pe_1_1_1_n57), .ZN(
        npu_inst_pe_1_1_1_n107) );
  AOI22_X1 npu_inst_pe_1_1_1_U102 ( .A1(npu_inst_int_data_y_2__1__0_), .A2(
        npu_inst_pe_1_1_1_n54), .B1(npu_inst_pe_1_1_1_n117), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_1_n53) );
  INV_X1 npu_inst_pe_1_1_1_U99 ( .A(npu_inst_pe_1_1_1_n53), .ZN(
        npu_inst_pe_1_1_1_n108) );
  AOI22_X1 npu_inst_pe_1_1_1_U98 ( .A1(npu_inst_int_data_y_2__1__0_), .A2(
        npu_inst_pe_1_1_1_n50), .B1(npu_inst_pe_1_1_1_n116), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_1_n49) );
  INV_X1 npu_inst_pe_1_1_1_U97 ( .A(npu_inst_pe_1_1_1_n49), .ZN(
        npu_inst_pe_1_1_1_n109) );
  AOI22_X1 npu_inst_pe_1_1_1_U96 ( .A1(npu_inst_int_data_y_2__1__0_), .A2(
        npu_inst_pe_1_1_1_n46), .B1(npu_inst_pe_1_1_1_n115), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_1_n45) );
  INV_X1 npu_inst_pe_1_1_1_U95 ( .A(npu_inst_pe_1_1_1_n45), .ZN(
        npu_inst_pe_1_1_1_n110) );
  AOI22_X1 npu_inst_pe_1_1_1_U94 ( .A1(npu_inst_int_data_y_2__1__0_), .A2(
        npu_inst_pe_1_1_1_n42), .B1(npu_inst_pe_1_1_1_n114), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_1_n41) );
  INV_X1 npu_inst_pe_1_1_1_U93 ( .A(npu_inst_pe_1_1_1_n41), .ZN(
        npu_inst_pe_1_1_1_n111) );
  AOI22_X1 npu_inst_pe_1_1_1_U92 ( .A1(npu_inst_int_data_y_2__1__1_), .A2(
        npu_inst_pe_1_1_1_n58), .B1(npu_inst_pe_1_1_1_n118), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_1_n59) );
  INV_X1 npu_inst_pe_1_1_1_U91 ( .A(npu_inst_pe_1_1_1_n59), .ZN(
        npu_inst_pe_1_1_1_n101) );
  AOI22_X1 npu_inst_pe_1_1_1_U90 ( .A1(npu_inst_int_data_y_2__1__1_), .A2(
        npu_inst_pe_1_1_1_n54), .B1(npu_inst_pe_1_1_1_n117), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_1_n55) );
  INV_X1 npu_inst_pe_1_1_1_U89 ( .A(npu_inst_pe_1_1_1_n55), .ZN(
        npu_inst_pe_1_1_1_n102) );
  AOI22_X1 npu_inst_pe_1_1_1_U88 ( .A1(npu_inst_int_data_y_2__1__1_), .A2(
        npu_inst_pe_1_1_1_n50), .B1(npu_inst_pe_1_1_1_n116), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_1_n51) );
  INV_X1 npu_inst_pe_1_1_1_U87 ( .A(npu_inst_pe_1_1_1_n51), .ZN(
        npu_inst_pe_1_1_1_n103) );
  AOI22_X1 npu_inst_pe_1_1_1_U86 ( .A1(npu_inst_int_data_y_2__1__1_), .A2(
        npu_inst_pe_1_1_1_n46), .B1(npu_inst_pe_1_1_1_n115), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_1_n47) );
  INV_X1 npu_inst_pe_1_1_1_U85 ( .A(npu_inst_pe_1_1_1_n47), .ZN(
        npu_inst_pe_1_1_1_n104) );
  AOI22_X1 npu_inst_pe_1_1_1_U84 ( .A1(npu_inst_int_data_y_2__1__1_), .A2(
        npu_inst_pe_1_1_1_n42), .B1(npu_inst_pe_1_1_1_n114), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_1_n43) );
  INV_X1 npu_inst_pe_1_1_1_U83 ( .A(npu_inst_pe_1_1_1_n43), .ZN(
        npu_inst_pe_1_1_1_n105) );
  AOI22_X1 npu_inst_pe_1_1_1_U82 ( .A1(npu_inst_pe_1_1_1_n38), .A2(
        npu_inst_int_data_y_2__1__1_), .B1(npu_inst_pe_1_1_1_n113), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_1_n39) );
  INV_X1 npu_inst_pe_1_1_1_U81 ( .A(npu_inst_pe_1_1_1_n39), .ZN(
        npu_inst_pe_1_1_1_n106) );
  AND2_X1 npu_inst_pe_1_1_1_U80 ( .A1(npu_inst_pe_1_1_1_N93), .A2(npu_inst_n41), .ZN(npu_inst_int_data_y_1__1__0_) );
  NAND2_X1 npu_inst_pe_1_1_1_U79 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_1_n60), .ZN(npu_inst_pe_1_1_1_n74) );
  OAI21_X1 npu_inst_pe_1_1_1_U78 ( .B1(npu_inst_pe_1_1_1_n63), .B2(
        npu_inst_pe_1_1_1_n60), .A(npu_inst_pe_1_1_1_n74), .ZN(
        npu_inst_pe_1_1_1_n97) );
  NAND2_X1 npu_inst_pe_1_1_1_U77 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_1_n60), .ZN(npu_inst_pe_1_1_1_n73) );
  OAI21_X1 npu_inst_pe_1_1_1_U76 ( .B1(npu_inst_pe_1_1_1_n61), .B2(
        npu_inst_pe_1_1_1_n60), .A(npu_inst_pe_1_1_1_n73), .ZN(
        npu_inst_pe_1_1_1_n96) );
  NAND2_X1 npu_inst_pe_1_1_1_U75 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_1_n56), .ZN(npu_inst_pe_1_1_1_n72) );
  OAI21_X1 npu_inst_pe_1_1_1_U74 ( .B1(npu_inst_pe_1_1_1_n63), .B2(
        npu_inst_pe_1_1_1_n56), .A(npu_inst_pe_1_1_1_n72), .ZN(
        npu_inst_pe_1_1_1_n95) );
  NAND2_X1 npu_inst_pe_1_1_1_U73 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_1_n56), .ZN(npu_inst_pe_1_1_1_n71) );
  OAI21_X1 npu_inst_pe_1_1_1_U72 ( .B1(npu_inst_pe_1_1_1_n61), .B2(
        npu_inst_pe_1_1_1_n56), .A(npu_inst_pe_1_1_1_n71), .ZN(
        npu_inst_pe_1_1_1_n94) );
  NAND2_X1 npu_inst_pe_1_1_1_U71 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_1_n52), .ZN(npu_inst_pe_1_1_1_n70) );
  OAI21_X1 npu_inst_pe_1_1_1_U70 ( .B1(npu_inst_pe_1_1_1_n63), .B2(
        npu_inst_pe_1_1_1_n52), .A(npu_inst_pe_1_1_1_n70), .ZN(
        npu_inst_pe_1_1_1_n93) );
  NAND2_X1 npu_inst_pe_1_1_1_U69 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_1_n52), .ZN(npu_inst_pe_1_1_1_n69) );
  OAI21_X1 npu_inst_pe_1_1_1_U68 ( .B1(npu_inst_pe_1_1_1_n61), .B2(
        npu_inst_pe_1_1_1_n52), .A(npu_inst_pe_1_1_1_n69), .ZN(
        npu_inst_pe_1_1_1_n92) );
  NAND2_X1 npu_inst_pe_1_1_1_U67 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_1_n48), .ZN(npu_inst_pe_1_1_1_n68) );
  OAI21_X1 npu_inst_pe_1_1_1_U66 ( .B1(npu_inst_pe_1_1_1_n63), .B2(
        npu_inst_pe_1_1_1_n48), .A(npu_inst_pe_1_1_1_n68), .ZN(
        npu_inst_pe_1_1_1_n91) );
  NAND2_X1 npu_inst_pe_1_1_1_U65 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_1_n48), .ZN(npu_inst_pe_1_1_1_n67) );
  OAI21_X1 npu_inst_pe_1_1_1_U64 ( .B1(npu_inst_pe_1_1_1_n61), .B2(
        npu_inst_pe_1_1_1_n48), .A(npu_inst_pe_1_1_1_n67), .ZN(
        npu_inst_pe_1_1_1_n90) );
  NAND2_X1 npu_inst_pe_1_1_1_U63 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_1_n44), .ZN(npu_inst_pe_1_1_1_n66) );
  OAI21_X1 npu_inst_pe_1_1_1_U62 ( .B1(npu_inst_pe_1_1_1_n63), .B2(
        npu_inst_pe_1_1_1_n44), .A(npu_inst_pe_1_1_1_n66), .ZN(
        npu_inst_pe_1_1_1_n89) );
  NAND2_X1 npu_inst_pe_1_1_1_U61 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_1_n44), .ZN(npu_inst_pe_1_1_1_n65) );
  OAI21_X1 npu_inst_pe_1_1_1_U60 ( .B1(npu_inst_pe_1_1_1_n61), .B2(
        npu_inst_pe_1_1_1_n44), .A(npu_inst_pe_1_1_1_n65), .ZN(
        npu_inst_pe_1_1_1_n88) );
  NAND2_X1 npu_inst_pe_1_1_1_U59 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_1_n40), .ZN(npu_inst_pe_1_1_1_n64) );
  OAI21_X1 npu_inst_pe_1_1_1_U58 ( .B1(npu_inst_pe_1_1_1_n63), .B2(
        npu_inst_pe_1_1_1_n40), .A(npu_inst_pe_1_1_1_n64), .ZN(
        npu_inst_pe_1_1_1_n87) );
  NAND2_X1 npu_inst_pe_1_1_1_U57 ( .A1(npu_inst_pe_1_1_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_1_n40), .ZN(npu_inst_pe_1_1_1_n62) );
  OAI21_X1 npu_inst_pe_1_1_1_U56 ( .B1(npu_inst_pe_1_1_1_n61), .B2(
        npu_inst_pe_1_1_1_n40), .A(npu_inst_pe_1_1_1_n62), .ZN(
        npu_inst_pe_1_1_1_n86) );
  AOI22_X1 npu_inst_pe_1_1_1_U55 ( .A1(npu_inst_pe_1_1_1_n38), .A2(
        npu_inst_int_data_y_2__1__0_), .B1(npu_inst_pe_1_1_1_n113), .B2(
        npu_inst_pe_1_1_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_1_n37) );
  INV_X1 npu_inst_pe_1_1_1_U54 ( .A(npu_inst_pe_1_1_1_n37), .ZN(
        npu_inst_pe_1_1_1_n112) );
  AND2_X1 npu_inst_pe_1_1_1_U53 ( .A1(npu_inst_n41), .A2(npu_inst_pe_1_1_1_N94), .ZN(npu_inst_int_data_y_1__1__1_) );
  AOI222_X1 npu_inst_pe_1_1_1_U52 ( .A1(npu_inst_int_data_res_2__1__0_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N73), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N65), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n84) );
  INV_X1 npu_inst_pe_1_1_1_U51 ( .A(npu_inst_pe_1_1_1_n84), .ZN(
        npu_inst_pe_1_1_1_n100) );
  AOI222_X1 npu_inst_pe_1_1_1_U50 ( .A1(npu_inst_pe_1_1_1_n1), .A2(
        npu_inst_int_data_res_2__1__7_), .B1(npu_inst_pe_1_1_1_N80), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N72), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n75) );
  INV_X1 npu_inst_pe_1_1_1_U49 ( .A(npu_inst_pe_1_1_1_n75), .ZN(
        npu_inst_pe_1_1_1_n32) );
  AOI222_X1 npu_inst_pe_1_1_1_U48 ( .A1(npu_inst_int_data_res_2__1__1_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N74), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N66), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n83) );
  INV_X1 npu_inst_pe_1_1_1_U47 ( .A(npu_inst_pe_1_1_1_n83), .ZN(
        npu_inst_pe_1_1_1_n99) );
  AOI222_X1 npu_inst_pe_1_1_1_U46 ( .A1(npu_inst_int_data_res_2__1__3_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N76), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N68), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n81) );
  INV_X1 npu_inst_pe_1_1_1_U45 ( .A(npu_inst_pe_1_1_1_n81), .ZN(
        npu_inst_pe_1_1_1_n36) );
  AOI222_X1 npu_inst_pe_1_1_1_U44 ( .A1(npu_inst_int_data_res_2__1__4_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N77), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N69), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n80) );
  INV_X1 npu_inst_pe_1_1_1_U43 ( .A(npu_inst_pe_1_1_1_n80), .ZN(
        npu_inst_pe_1_1_1_n35) );
  AOI222_X1 npu_inst_pe_1_1_1_U42 ( .A1(npu_inst_int_data_res_2__1__5_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N78), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N70), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n79) );
  INV_X1 npu_inst_pe_1_1_1_U41 ( .A(npu_inst_pe_1_1_1_n79), .ZN(
        npu_inst_pe_1_1_1_n34) );
  AOI222_X1 npu_inst_pe_1_1_1_U40 ( .A1(npu_inst_int_data_res_2__1__6_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N79), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N71), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n78) );
  INV_X1 npu_inst_pe_1_1_1_U39 ( .A(npu_inst_pe_1_1_1_n78), .ZN(
        npu_inst_pe_1_1_1_n33) );
  AND2_X1 npu_inst_pe_1_1_1_U38 ( .A1(npu_inst_int_data_x_1__1__1_), .A2(
        npu_inst_pe_1_1_1_int_q_weight_1_), .ZN(npu_inst_pe_1_1_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_1_U37 ( .A1(npu_inst_int_data_x_1__1__0_), .A2(
        npu_inst_pe_1_1_1_int_q_weight_1_), .ZN(npu_inst_pe_1_1_1_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_1_1_U36 ( .A(npu_inst_pe_1_1_1_int_data_1_), .ZN(
        npu_inst_pe_1_1_1_n13) );
  NOR3_X1 npu_inst_pe_1_1_1_U35 ( .A1(npu_inst_pe_1_1_1_n26), .A2(npu_inst_n41), .A3(npu_inst_int_ckg[54]), .ZN(npu_inst_pe_1_1_1_n85) );
  OR2_X1 npu_inst_pe_1_1_1_U34 ( .A1(npu_inst_pe_1_1_1_n85), .A2(
        npu_inst_pe_1_1_1_n1), .ZN(npu_inst_pe_1_1_1_N84) );
  AOI222_X1 npu_inst_pe_1_1_1_U33 ( .A1(npu_inst_int_data_res_2__1__2_), .A2(
        npu_inst_pe_1_1_1_n1), .B1(npu_inst_pe_1_1_1_N75), .B2(
        npu_inst_pe_1_1_1_n76), .C1(npu_inst_pe_1_1_1_N67), .C2(
        npu_inst_pe_1_1_1_n77), .ZN(npu_inst_pe_1_1_1_n82) );
  INV_X1 npu_inst_pe_1_1_1_U32 ( .A(npu_inst_pe_1_1_1_n82), .ZN(
        npu_inst_pe_1_1_1_n98) );
  AOI22_X1 npu_inst_pe_1_1_1_U31 ( .A1(npu_inst_n41), .A2(
        npu_inst_int_data_y_2__1__1_), .B1(npu_inst_pe_1_1_1_n2), .B2(
        npu_inst_int_data_x_1__2__1_), .ZN(npu_inst_pe_1_1_1_n63) );
  AOI22_X1 npu_inst_pe_1_1_1_U30 ( .A1(npu_inst_n41), .A2(
        npu_inst_int_data_y_2__1__0_), .B1(npu_inst_pe_1_1_1_n2), .B2(
        npu_inst_int_data_x_1__2__0_), .ZN(npu_inst_pe_1_1_1_n61) );
  INV_X1 npu_inst_pe_1_1_1_U29 ( .A(npu_inst_pe_1_1_1_int_data_0_), .ZN(
        npu_inst_pe_1_1_1_n12) );
  INV_X1 npu_inst_pe_1_1_1_U28 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_1_1_n4)
         );
  OR3_X1 npu_inst_pe_1_1_1_U27 ( .A1(npu_inst_pe_1_1_1_n5), .A2(
        npu_inst_pe_1_1_1_n7), .A3(npu_inst_pe_1_1_1_n4), .ZN(
        npu_inst_pe_1_1_1_n56) );
  OR3_X1 npu_inst_pe_1_1_1_U26 ( .A1(npu_inst_pe_1_1_1_n4), .A2(
        npu_inst_pe_1_1_1_n7), .A3(npu_inst_pe_1_1_1_n6), .ZN(
        npu_inst_pe_1_1_1_n48) );
  INV_X1 npu_inst_pe_1_1_1_U25 ( .A(npu_inst_pe_1_1_1_n4), .ZN(
        npu_inst_pe_1_1_1_n3) );
  OR3_X1 npu_inst_pe_1_1_1_U24 ( .A1(npu_inst_pe_1_1_1_n3), .A2(
        npu_inst_pe_1_1_1_n7), .A3(npu_inst_pe_1_1_1_n6), .ZN(
        npu_inst_pe_1_1_1_n52) );
  OR3_X1 npu_inst_pe_1_1_1_U23 ( .A1(npu_inst_pe_1_1_1_n5), .A2(
        npu_inst_pe_1_1_1_n7), .A3(npu_inst_pe_1_1_1_n3), .ZN(
        npu_inst_pe_1_1_1_n60) );
  BUF_X1 npu_inst_pe_1_1_1_U22 ( .A(npu_inst_n29), .Z(npu_inst_pe_1_1_1_n1) );
  NOR2_X1 npu_inst_pe_1_1_1_U21 ( .A1(npu_inst_pe_1_1_1_n60), .A2(
        npu_inst_pe_1_1_1_n2), .ZN(npu_inst_pe_1_1_1_n58) );
  NOR2_X1 npu_inst_pe_1_1_1_U20 ( .A1(npu_inst_pe_1_1_1_n56), .A2(
        npu_inst_pe_1_1_1_n2), .ZN(npu_inst_pe_1_1_1_n54) );
  NOR2_X1 npu_inst_pe_1_1_1_U19 ( .A1(npu_inst_pe_1_1_1_n52), .A2(
        npu_inst_pe_1_1_1_n2), .ZN(npu_inst_pe_1_1_1_n50) );
  NOR2_X1 npu_inst_pe_1_1_1_U18 ( .A1(npu_inst_pe_1_1_1_n48), .A2(
        npu_inst_pe_1_1_1_n2), .ZN(npu_inst_pe_1_1_1_n46) );
  NOR2_X1 npu_inst_pe_1_1_1_U17 ( .A1(npu_inst_pe_1_1_1_n40), .A2(
        npu_inst_pe_1_1_1_n2), .ZN(npu_inst_pe_1_1_1_n38) );
  NOR2_X1 npu_inst_pe_1_1_1_U16 ( .A1(npu_inst_pe_1_1_1_n44), .A2(
        npu_inst_pe_1_1_1_n2), .ZN(npu_inst_pe_1_1_1_n42) );
  BUF_X1 npu_inst_pe_1_1_1_U15 ( .A(npu_inst_n87), .Z(npu_inst_pe_1_1_1_n7) );
  INV_X1 npu_inst_pe_1_1_1_U14 ( .A(npu_inst_n108), .ZN(npu_inst_pe_1_1_1_n11)
         );
  INV_X1 npu_inst_pe_1_1_1_U13 ( .A(npu_inst_pe_1_1_1_n38), .ZN(
        npu_inst_pe_1_1_1_n113) );
  INV_X1 npu_inst_pe_1_1_1_U12 ( .A(npu_inst_pe_1_1_1_n58), .ZN(
        npu_inst_pe_1_1_1_n118) );
  INV_X1 npu_inst_pe_1_1_1_U11 ( .A(npu_inst_pe_1_1_1_n54), .ZN(
        npu_inst_pe_1_1_1_n117) );
  INV_X1 npu_inst_pe_1_1_1_U10 ( .A(npu_inst_pe_1_1_1_n50), .ZN(
        npu_inst_pe_1_1_1_n116) );
  INV_X1 npu_inst_pe_1_1_1_U9 ( .A(npu_inst_pe_1_1_1_n46), .ZN(
        npu_inst_pe_1_1_1_n115) );
  INV_X1 npu_inst_pe_1_1_1_U8 ( .A(npu_inst_pe_1_1_1_n42), .ZN(
        npu_inst_pe_1_1_1_n114) );
  BUF_X1 npu_inst_pe_1_1_1_U7 ( .A(npu_inst_pe_1_1_1_n11), .Z(
        npu_inst_pe_1_1_1_n10) );
  BUF_X1 npu_inst_pe_1_1_1_U6 ( .A(npu_inst_pe_1_1_1_n11), .Z(
        npu_inst_pe_1_1_1_n9) );
  BUF_X1 npu_inst_pe_1_1_1_U5 ( .A(npu_inst_pe_1_1_1_n11), .Z(
        npu_inst_pe_1_1_1_n8) );
  NOR2_X1 npu_inst_pe_1_1_1_U4 ( .A1(npu_inst_pe_1_1_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_1_n1), .ZN(npu_inst_pe_1_1_1_n76) );
  NOR2_X1 npu_inst_pe_1_1_1_U3 ( .A1(npu_inst_pe_1_1_1_n27), .A2(
        npu_inst_pe_1_1_1_n1), .ZN(npu_inst_pe_1_1_1_n77) );
  FA_X1 npu_inst_pe_1_1_1_sub_77_U2_1 ( .A(npu_inst_int_data_res_1__1__1_), 
        .B(npu_inst_pe_1_1_1_n13), .CI(npu_inst_pe_1_1_1_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_1_1_sub_77_carry_2_), .S(npu_inst_pe_1_1_1_N66) );
  FA_X1 npu_inst_pe_1_1_1_add_79_U1_1 ( .A(npu_inst_int_data_res_1__1__1_), 
        .B(npu_inst_pe_1_1_1_int_data_1_), .CI(
        npu_inst_pe_1_1_1_add_79_carry_1_), .CO(
        npu_inst_pe_1_1_1_add_79_carry_2_), .S(npu_inst_pe_1_1_1_N74) );
  NAND3_X1 npu_inst_pe_1_1_1_U101 ( .A1(npu_inst_pe_1_1_1_n4), .A2(
        npu_inst_pe_1_1_1_n6), .A3(npu_inst_pe_1_1_1_n7), .ZN(
        npu_inst_pe_1_1_1_n44) );
  NAND3_X1 npu_inst_pe_1_1_1_U100 ( .A1(npu_inst_pe_1_1_1_n3), .A2(
        npu_inst_pe_1_1_1_n6), .A3(npu_inst_pe_1_1_1_n7), .ZN(
        npu_inst_pe_1_1_1_n40) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_1_n33), .CK(
        npu_inst_pe_1_1_1_net4271), .RN(npu_inst_pe_1_1_1_n8), .Q(
        npu_inst_int_data_res_1__1__6_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_1_n34), .CK(
        npu_inst_pe_1_1_1_net4271), .RN(npu_inst_pe_1_1_1_n8), .Q(
        npu_inst_int_data_res_1__1__5_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_1_n35), .CK(
        npu_inst_pe_1_1_1_net4271), .RN(npu_inst_pe_1_1_1_n8), .Q(
        npu_inst_int_data_res_1__1__4_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_1_n36), .CK(
        npu_inst_pe_1_1_1_net4271), .RN(npu_inst_pe_1_1_1_n8), .Q(
        npu_inst_int_data_res_1__1__3_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_1_n98), .CK(
        npu_inst_pe_1_1_1_net4271), .RN(npu_inst_pe_1_1_1_n8), .Q(
        npu_inst_int_data_res_1__1__2_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_1_n99), .CK(
        npu_inst_pe_1_1_1_net4271), .RN(npu_inst_pe_1_1_1_n8), .Q(
        npu_inst_int_data_res_1__1__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_1_n32), .CK(
        npu_inst_pe_1_1_1_net4271), .RN(npu_inst_pe_1_1_1_n8), .Q(
        npu_inst_int_data_res_1__1__7_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_1_n100), 
        .CK(npu_inst_pe_1_1_1_net4271), .RN(npu_inst_pe_1_1_1_n8), .Q(
        npu_inst_int_data_res_1__1__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_weight_reg_0_ ( .D(npu_inst_n94), .CK(
        npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n8), .Q(
        npu_inst_pe_1_1_1_int_q_weight_0_), .QN(npu_inst_pe_1_1_1_n27) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_weight_reg_1_ ( .D(npu_inst_n100), .CK(
        npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n8), .Q(
        npu_inst_pe_1_1_1_int_q_weight_1_), .QN(npu_inst_pe_1_1_1_n26) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_1_n112), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n8), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_1_n106), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n8), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_1_n111), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_1_n105), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_1_n110), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_1_n104), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_1_n109), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_1_n103), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_1_n108), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_1_n102), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_1_n107), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_1_n101), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_1_n86), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_1_n87), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n9), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_1_n88), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_1_n89), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_1_n90), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_1_n91), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_1_n92), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_1_n93), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_1_n94), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_1_n95), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_1_n96), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_1_n97), 
        .CK(npu_inst_pe_1_1_1_net4277), .RN(npu_inst_pe_1_1_1_n10), .Q(
        npu_inst_pe_1_1_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_1_net4271) );
  CLKGATETST_X1 npu_inst_pe_1_1_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n47), .SE(1'b0), .GCK(npu_inst_pe_1_1_1_net4277) );
  MUX2_X1 npu_inst_pe_1_1_2_U153 ( .A(npu_inst_pe_1_1_2_n31), .B(
        npu_inst_pe_1_1_2_n28), .S(npu_inst_pe_1_1_2_n7), .Z(
        npu_inst_pe_1_1_2_N93) );
  MUX2_X1 npu_inst_pe_1_1_2_U152 ( .A(npu_inst_pe_1_1_2_n30), .B(
        npu_inst_pe_1_1_2_n29), .S(npu_inst_pe_1_1_2_n5), .Z(
        npu_inst_pe_1_1_2_n31) );
  MUX2_X1 npu_inst_pe_1_1_2_U151 ( .A(npu_inst_pe_1_1_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_2_n3), .Z(
        npu_inst_pe_1_1_2_n30) );
  MUX2_X1 npu_inst_pe_1_1_2_U150 ( .A(npu_inst_pe_1_1_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_2_n3), .Z(
        npu_inst_pe_1_1_2_n29) );
  MUX2_X1 npu_inst_pe_1_1_2_U149 ( .A(npu_inst_pe_1_1_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_2_n3), .Z(
        npu_inst_pe_1_1_2_n28) );
  MUX2_X1 npu_inst_pe_1_1_2_U148 ( .A(npu_inst_pe_1_1_2_n25), .B(
        npu_inst_pe_1_1_2_n22), .S(npu_inst_pe_1_1_2_n7), .Z(
        npu_inst_pe_1_1_2_N94) );
  MUX2_X1 npu_inst_pe_1_1_2_U147 ( .A(npu_inst_pe_1_1_2_n24), .B(
        npu_inst_pe_1_1_2_n23), .S(npu_inst_pe_1_1_2_n5), .Z(
        npu_inst_pe_1_1_2_n25) );
  MUX2_X1 npu_inst_pe_1_1_2_U146 ( .A(npu_inst_pe_1_1_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_2_n3), .Z(
        npu_inst_pe_1_1_2_n24) );
  MUX2_X1 npu_inst_pe_1_1_2_U145 ( .A(npu_inst_pe_1_1_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_2_n3), .Z(
        npu_inst_pe_1_1_2_n23) );
  MUX2_X1 npu_inst_pe_1_1_2_U144 ( .A(npu_inst_pe_1_1_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_2_n3), .Z(
        npu_inst_pe_1_1_2_n22) );
  MUX2_X1 npu_inst_pe_1_1_2_U143 ( .A(npu_inst_pe_1_1_2_n21), .B(
        npu_inst_pe_1_1_2_n18), .S(npu_inst_pe_1_1_2_n7), .Z(
        npu_inst_int_data_x_1__2__1_) );
  MUX2_X1 npu_inst_pe_1_1_2_U142 ( .A(npu_inst_pe_1_1_2_n20), .B(
        npu_inst_pe_1_1_2_n19), .S(npu_inst_pe_1_1_2_n5), .Z(
        npu_inst_pe_1_1_2_n21) );
  MUX2_X1 npu_inst_pe_1_1_2_U141 ( .A(npu_inst_pe_1_1_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_2_n3), .Z(
        npu_inst_pe_1_1_2_n20) );
  MUX2_X1 npu_inst_pe_1_1_2_U140 ( .A(npu_inst_pe_1_1_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_2_n3), .Z(
        npu_inst_pe_1_1_2_n19) );
  MUX2_X1 npu_inst_pe_1_1_2_U139 ( .A(npu_inst_pe_1_1_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_2_n3), .Z(
        npu_inst_pe_1_1_2_n18) );
  MUX2_X1 npu_inst_pe_1_1_2_U138 ( .A(npu_inst_pe_1_1_2_n17), .B(
        npu_inst_pe_1_1_2_n14), .S(npu_inst_pe_1_1_2_n7), .Z(
        npu_inst_int_data_x_1__2__0_) );
  MUX2_X1 npu_inst_pe_1_1_2_U137 ( .A(npu_inst_pe_1_1_2_n16), .B(
        npu_inst_pe_1_1_2_n15), .S(npu_inst_pe_1_1_2_n5), .Z(
        npu_inst_pe_1_1_2_n17) );
  MUX2_X1 npu_inst_pe_1_1_2_U136 ( .A(npu_inst_pe_1_1_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_2_n3), .Z(
        npu_inst_pe_1_1_2_n16) );
  MUX2_X1 npu_inst_pe_1_1_2_U135 ( .A(npu_inst_pe_1_1_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_2_n3), .Z(
        npu_inst_pe_1_1_2_n15) );
  MUX2_X1 npu_inst_pe_1_1_2_U134 ( .A(npu_inst_pe_1_1_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_2_n3), .Z(
        npu_inst_pe_1_1_2_n14) );
  XOR2_X1 npu_inst_pe_1_1_2_U133 ( .A(npu_inst_pe_1_1_2_int_data_0_), .B(
        npu_inst_int_data_res_1__2__0_), .Z(npu_inst_pe_1_1_2_N73) );
  AND2_X1 npu_inst_pe_1_1_2_U132 ( .A1(npu_inst_int_data_res_1__2__0_), .A2(
        npu_inst_pe_1_1_2_int_data_0_), .ZN(npu_inst_pe_1_1_2_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_2_U131 ( .A(npu_inst_int_data_res_1__2__0_), .B(
        npu_inst_pe_1_1_2_n12), .ZN(npu_inst_pe_1_1_2_N65) );
  OR2_X1 npu_inst_pe_1_1_2_U130 ( .A1(npu_inst_pe_1_1_2_n12), .A2(
        npu_inst_int_data_res_1__2__0_), .ZN(npu_inst_pe_1_1_2_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_2_U129 ( .A(npu_inst_int_data_res_1__2__2_), .B(
        npu_inst_pe_1_1_2_add_79_carry_2_), .Z(npu_inst_pe_1_1_2_N75) );
  AND2_X1 npu_inst_pe_1_1_2_U128 ( .A1(npu_inst_pe_1_1_2_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_1__2__2_), .ZN(
        npu_inst_pe_1_1_2_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_2_U127 ( .A(npu_inst_int_data_res_1__2__3_), .B(
        npu_inst_pe_1_1_2_add_79_carry_3_), .Z(npu_inst_pe_1_1_2_N76) );
  AND2_X1 npu_inst_pe_1_1_2_U126 ( .A1(npu_inst_pe_1_1_2_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_1__2__3_), .ZN(
        npu_inst_pe_1_1_2_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_2_U125 ( .A(npu_inst_int_data_res_1__2__4_), .B(
        npu_inst_pe_1_1_2_add_79_carry_4_), .Z(npu_inst_pe_1_1_2_N77) );
  AND2_X1 npu_inst_pe_1_1_2_U124 ( .A1(npu_inst_pe_1_1_2_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_1__2__4_), .ZN(
        npu_inst_pe_1_1_2_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_2_U123 ( .A(npu_inst_int_data_res_1__2__5_), .B(
        npu_inst_pe_1_1_2_add_79_carry_5_), .Z(npu_inst_pe_1_1_2_N78) );
  AND2_X1 npu_inst_pe_1_1_2_U122 ( .A1(npu_inst_pe_1_1_2_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_1__2__5_), .ZN(
        npu_inst_pe_1_1_2_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_2_U121 ( .A(npu_inst_int_data_res_1__2__6_), .B(
        npu_inst_pe_1_1_2_add_79_carry_6_), .Z(npu_inst_pe_1_1_2_N79) );
  AND2_X1 npu_inst_pe_1_1_2_U120 ( .A1(npu_inst_pe_1_1_2_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_1__2__6_), .ZN(
        npu_inst_pe_1_1_2_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_2_U119 ( .A(npu_inst_int_data_res_1__2__7_), .B(
        npu_inst_pe_1_1_2_add_79_carry_7_), .Z(npu_inst_pe_1_1_2_N80) );
  XNOR2_X1 npu_inst_pe_1_1_2_U118 ( .A(npu_inst_pe_1_1_2_sub_77_carry_2_), .B(
        npu_inst_int_data_res_1__2__2_), .ZN(npu_inst_pe_1_1_2_N67) );
  OR2_X1 npu_inst_pe_1_1_2_U117 ( .A1(npu_inst_int_data_res_1__2__2_), .A2(
        npu_inst_pe_1_1_2_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_1_2_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_2_U116 ( .A(npu_inst_pe_1_1_2_sub_77_carry_3_), .B(
        npu_inst_int_data_res_1__2__3_), .ZN(npu_inst_pe_1_1_2_N68) );
  OR2_X1 npu_inst_pe_1_1_2_U115 ( .A1(npu_inst_int_data_res_1__2__3_), .A2(
        npu_inst_pe_1_1_2_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_1_2_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_2_U114 ( .A(npu_inst_pe_1_1_2_sub_77_carry_4_), .B(
        npu_inst_int_data_res_1__2__4_), .ZN(npu_inst_pe_1_1_2_N69) );
  OR2_X1 npu_inst_pe_1_1_2_U113 ( .A1(npu_inst_int_data_res_1__2__4_), .A2(
        npu_inst_pe_1_1_2_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_1_2_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_2_U112 ( .A(npu_inst_pe_1_1_2_sub_77_carry_5_), .B(
        npu_inst_int_data_res_1__2__5_), .ZN(npu_inst_pe_1_1_2_N70) );
  OR2_X1 npu_inst_pe_1_1_2_U111 ( .A1(npu_inst_int_data_res_1__2__5_), .A2(
        npu_inst_pe_1_1_2_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_1_2_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_2_U110 ( .A(npu_inst_pe_1_1_2_sub_77_carry_6_), .B(
        npu_inst_int_data_res_1__2__6_), .ZN(npu_inst_pe_1_1_2_N71) );
  OR2_X1 npu_inst_pe_1_1_2_U109 ( .A1(npu_inst_int_data_res_1__2__6_), .A2(
        npu_inst_pe_1_1_2_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_1_2_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_2_U108 ( .A(npu_inst_int_data_res_1__2__7_), .B(
        npu_inst_pe_1_1_2_sub_77_carry_7_), .ZN(npu_inst_pe_1_1_2_N72) );
  INV_X1 npu_inst_pe_1_1_2_U107 ( .A(npu_inst_n61), .ZN(npu_inst_pe_1_1_2_n6)
         );
  INV_X1 npu_inst_pe_1_1_2_U106 ( .A(npu_inst_pe_1_1_2_n6), .ZN(
        npu_inst_pe_1_1_2_n5) );
  INV_X1 npu_inst_pe_1_1_2_U105 ( .A(npu_inst_n41), .ZN(npu_inst_pe_1_1_2_n2)
         );
  AOI22_X1 npu_inst_pe_1_1_2_U104 ( .A1(npu_inst_int_data_y_2__2__0_), .A2(
        npu_inst_pe_1_1_2_n58), .B1(npu_inst_pe_1_1_2_n118), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_2_n57) );
  INV_X1 npu_inst_pe_1_1_2_U103 ( .A(npu_inst_pe_1_1_2_n57), .ZN(
        npu_inst_pe_1_1_2_n107) );
  AOI22_X1 npu_inst_pe_1_1_2_U102 ( .A1(npu_inst_int_data_y_2__2__0_), .A2(
        npu_inst_pe_1_1_2_n54), .B1(npu_inst_pe_1_1_2_n117), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_2_n53) );
  INV_X1 npu_inst_pe_1_1_2_U99 ( .A(npu_inst_pe_1_1_2_n53), .ZN(
        npu_inst_pe_1_1_2_n108) );
  AOI22_X1 npu_inst_pe_1_1_2_U98 ( .A1(npu_inst_int_data_y_2__2__0_), .A2(
        npu_inst_pe_1_1_2_n50), .B1(npu_inst_pe_1_1_2_n116), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_2_n49) );
  INV_X1 npu_inst_pe_1_1_2_U97 ( .A(npu_inst_pe_1_1_2_n49), .ZN(
        npu_inst_pe_1_1_2_n109) );
  AOI22_X1 npu_inst_pe_1_1_2_U96 ( .A1(npu_inst_int_data_y_2__2__0_), .A2(
        npu_inst_pe_1_1_2_n46), .B1(npu_inst_pe_1_1_2_n115), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_2_n45) );
  INV_X1 npu_inst_pe_1_1_2_U95 ( .A(npu_inst_pe_1_1_2_n45), .ZN(
        npu_inst_pe_1_1_2_n110) );
  AOI22_X1 npu_inst_pe_1_1_2_U94 ( .A1(npu_inst_int_data_y_2__2__0_), .A2(
        npu_inst_pe_1_1_2_n42), .B1(npu_inst_pe_1_1_2_n114), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_2_n41) );
  INV_X1 npu_inst_pe_1_1_2_U93 ( .A(npu_inst_pe_1_1_2_n41), .ZN(
        npu_inst_pe_1_1_2_n111) );
  AOI22_X1 npu_inst_pe_1_1_2_U92 ( .A1(npu_inst_int_data_y_2__2__1_), .A2(
        npu_inst_pe_1_1_2_n58), .B1(npu_inst_pe_1_1_2_n118), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_2_n59) );
  INV_X1 npu_inst_pe_1_1_2_U91 ( .A(npu_inst_pe_1_1_2_n59), .ZN(
        npu_inst_pe_1_1_2_n101) );
  AOI22_X1 npu_inst_pe_1_1_2_U90 ( .A1(npu_inst_int_data_y_2__2__1_), .A2(
        npu_inst_pe_1_1_2_n54), .B1(npu_inst_pe_1_1_2_n117), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_2_n55) );
  INV_X1 npu_inst_pe_1_1_2_U89 ( .A(npu_inst_pe_1_1_2_n55), .ZN(
        npu_inst_pe_1_1_2_n102) );
  AOI22_X1 npu_inst_pe_1_1_2_U88 ( .A1(npu_inst_int_data_y_2__2__1_), .A2(
        npu_inst_pe_1_1_2_n50), .B1(npu_inst_pe_1_1_2_n116), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_2_n51) );
  INV_X1 npu_inst_pe_1_1_2_U87 ( .A(npu_inst_pe_1_1_2_n51), .ZN(
        npu_inst_pe_1_1_2_n103) );
  AOI22_X1 npu_inst_pe_1_1_2_U86 ( .A1(npu_inst_int_data_y_2__2__1_), .A2(
        npu_inst_pe_1_1_2_n46), .B1(npu_inst_pe_1_1_2_n115), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_2_n47) );
  INV_X1 npu_inst_pe_1_1_2_U85 ( .A(npu_inst_pe_1_1_2_n47), .ZN(
        npu_inst_pe_1_1_2_n104) );
  AOI22_X1 npu_inst_pe_1_1_2_U84 ( .A1(npu_inst_int_data_y_2__2__1_), .A2(
        npu_inst_pe_1_1_2_n42), .B1(npu_inst_pe_1_1_2_n114), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_2_n43) );
  INV_X1 npu_inst_pe_1_1_2_U83 ( .A(npu_inst_pe_1_1_2_n43), .ZN(
        npu_inst_pe_1_1_2_n105) );
  AOI22_X1 npu_inst_pe_1_1_2_U82 ( .A1(npu_inst_pe_1_1_2_n38), .A2(
        npu_inst_int_data_y_2__2__1_), .B1(npu_inst_pe_1_1_2_n113), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_2_n39) );
  INV_X1 npu_inst_pe_1_1_2_U81 ( .A(npu_inst_pe_1_1_2_n39), .ZN(
        npu_inst_pe_1_1_2_n106) );
  AND2_X1 npu_inst_pe_1_1_2_U80 ( .A1(npu_inst_pe_1_1_2_N93), .A2(npu_inst_n41), .ZN(npu_inst_int_data_y_1__2__0_) );
  NAND2_X1 npu_inst_pe_1_1_2_U79 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_2_n60), .ZN(npu_inst_pe_1_1_2_n74) );
  OAI21_X1 npu_inst_pe_1_1_2_U78 ( .B1(npu_inst_pe_1_1_2_n63), .B2(
        npu_inst_pe_1_1_2_n60), .A(npu_inst_pe_1_1_2_n74), .ZN(
        npu_inst_pe_1_1_2_n97) );
  NAND2_X1 npu_inst_pe_1_1_2_U77 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_2_n60), .ZN(npu_inst_pe_1_1_2_n73) );
  OAI21_X1 npu_inst_pe_1_1_2_U76 ( .B1(npu_inst_pe_1_1_2_n61), .B2(
        npu_inst_pe_1_1_2_n60), .A(npu_inst_pe_1_1_2_n73), .ZN(
        npu_inst_pe_1_1_2_n96) );
  NAND2_X1 npu_inst_pe_1_1_2_U75 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_2_n56), .ZN(npu_inst_pe_1_1_2_n72) );
  OAI21_X1 npu_inst_pe_1_1_2_U74 ( .B1(npu_inst_pe_1_1_2_n63), .B2(
        npu_inst_pe_1_1_2_n56), .A(npu_inst_pe_1_1_2_n72), .ZN(
        npu_inst_pe_1_1_2_n95) );
  NAND2_X1 npu_inst_pe_1_1_2_U73 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_2_n56), .ZN(npu_inst_pe_1_1_2_n71) );
  OAI21_X1 npu_inst_pe_1_1_2_U72 ( .B1(npu_inst_pe_1_1_2_n61), .B2(
        npu_inst_pe_1_1_2_n56), .A(npu_inst_pe_1_1_2_n71), .ZN(
        npu_inst_pe_1_1_2_n94) );
  NAND2_X1 npu_inst_pe_1_1_2_U71 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_2_n52), .ZN(npu_inst_pe_1_1_2_n70) );
  OAI21_X1 npu_inst_pe_1_1_2_U70 ( .B1(npu_inst_pe_1_1_2_n63), .B2(
        npu_inst_pe_1_1_2_n52), .A(npu_inst_pe_1_1_2_n70), .ZN(
        npu_inst_pe_1_1_2_n93) );
  NAND2_X1 npu_inst_pe_1_1_2_U69 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_2_n52), .ZN(npu_inst_pe_1_1_2_n69) );
  OAI21_X1 npu_inst_pe_1_1_2_U68 ( .B1(npu_inst_pe_1_1_2_n61), .B2(
        npu_inst_pe_1_1_2_n52), .A(npu_inst_pe_1_1_2_n69), .ZN(
        npu_inst_pe_1_1_2_n92) );
  NAND2_X1 npu_inst_pe_1_1_2_U67 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_2_n48), .ZN(npu_inst_pe_1_1_2_n68) );
  OAI21_X1 npu_inst_pe_1_1_2_U66 ( .B1(npu_inst_pe_1_1_2_n63), .B2(
        npu_inst_pe_1_1_2_n48), .A(npu_inst_pe_1_1_2_n68), .ZN(
        npu_inst_pe_1_1_2_n91) );
  NAND2_X1 npu_inst_pe_1_1_2_U65 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_2_n48), .ZN(npu_inst_pe_1_1_2_n67) );
  OAI21_X1 npu_inst_pe_1_1_2_U64 ( .B1(npu_inst_pe_1_1_2_n61), .B2(
        npu_inst_pe_1_1_2_n48), .A(npu_inst_pe_1_1_2_n67), .ZN(
        npu_inst_pe_1_1_2_n90) );
  NAND2_X1 npu_inst_pe_1_1_2_U63 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_2_n44), .ZN(npu_inst_pe_1_1_2_n66) );
  OAI21_X1 npu_inst_pe_1_1_2_U62 ( .B1(npu_inst_pe_1_1_2_n63), .B2(
        npu_inst_pe_1_1_2_n44), .A(npu_inst_pe_1_1_2_n66), .ZN(
        npu_inst_pe_1_1_2_n89) );
  NAND2_X1 npu_inst_pe_1_1_2_U61 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_2_n44), .ZN(npu_inst_pe_1_1_2_n65) );
  OAI21_X1 npu_inst_pe_1_1_2_U60 ( .B1(npu_inst_pe_1_1_2_n61), .B2(
        npu_inst_pe_1_1_2_n44), .A(npu_inst_pe_1_1_2_n65), .ZN(
        npu_inst_pe_1_1_2_n88) );
  NAND2_X1 npu_inst_pe_1_1_2_U59 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_2_n40), .ZN(npu_inst_pe_1_1_2_n64) );
  OAI21_X1 npu_inst_pe_1_1_2_U58 ( .B1(npu_inst_pe_1_1_2_n63), .B2(
        npu_inst_pe_1_1_2_n40), .A(npu_inst_pe_1_1_2_n64), .ZN(
        npu_inst_pe_1_1_2_n87) );
  NAND2_X1 npu_inst_pe_1_1_2_U57 ( .A1(npu_inst_pe_1_1_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_2_n40), .ZN(npu_inst_pe_1_1_2_n62) );
  OAI21_X1 npu_inst_pe_1_1_2_U56 ( .B1(npu_inst_pe_1_1_2_n61), .B2(
        npu_inst_pe_1_1_2_n40), .A(npu_inst_pe_1_1_2_n62), .ZN(
        npu_inst_pe_1_1_2_n86) );
  AOI22_X1 npu_inst_pe_1_1_2_U55 ( .A1(npu_inst_pe_1_1_2_n38), .A2(
        npu_inst_int_data_y_2__2__0_), .B1(npu_inst_pe_1_1_2_n113), .B2(
        npu_inst_pe_1_1_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_2_n37) );
  INV_X1 npu_inst_pe_1_1_2_U54 ( .A(npu_inst_pe_1_1_2_n37), .ZN(
        npu_inst_pe_1_1_2_n112) );
  AND2_X1 npu_inst_pe_1_1_2_U53 ( .A1(npu_inst_n41), .A2(npu_inst_pe_1_1_2_N94), .ZN(npu_inst_int_data_y_1__2__1_) );
  AOI222_X1 npu_inst_pe_1_1_2_U52 ( .A1(npu_inst_int_data_res_2__2__0_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N73), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N65), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n84) );
  INV_X1 npu_inst_pe_1_1_2_U51 ( .A(npu_inst_pe_1_1_2_n84), .ZN(
        npu_inst_pe_1_1_2_n100) );
  AOI222_X1 npu_inst_pe_1_1_2_U50 ( .A1(npu_inst_pe_1_1_2_n1), .A2(
        npu_inst_int_data_res_2__2__7_), .B1(npu_inst_pe_1_1_2_N80), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N72), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n75) );
  INV_X1 npu_inst_pe_1_1_2_U49 ( .A(npu_inst_pe_1_1_2_n75), .ZN(
        npu_inst_pe_1_1_2_n32) );
  AOI222_X1 npu_inst_pe_1_1_2_U48 ( .A1(npu_inst_int_data_res_2__2__1_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N74), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N66), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n83) );
  INV_X1 npu_inst_pe_1_1_2_U47 ( .A(npu_inst_pe_1_1_2_n83), .ZN(
        npu_inst_pe_1_1_2_n99) );
  AOI222_X1 npu_inst_pe_1_1_2_U46 ( .A1(npu_inst_int_data_res_2__2__3_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N76), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N68), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n81) );
  INV_X1 npu_inst_pe_1_1_2_U45 ( .A(npu_inst_pe_1_1_2_n81), .ZN(
        npu_inst_pe_1_1_2_n36) );
  AOI222_X1 npu_inst_pe_1_1_2_U44 ( .A1(npu_inst_int_data_res_2__2__4_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N77), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N69), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n80) );
  INV_X1 npu_inst_pe_1_1_2_U43 ( .A(npu_inst_pe_1_1_2_n80), .ZN(
        npu_inst_pe_1_1_2_n35) );
  AOI222_X1 npu_inst_pe_1_1_2_U42 ( .A1(npu_inst_int_data_res_2__2__5_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N78), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N70), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n79) );
  INV_X1 npu_inst_pe_1_1_2_U41 ( .A(npu_inst_pe_1_1_2_n79), .ZN(
        npu_inst_pe_1_1_2_n34) );
  AOI222_X1 npu_inst_pe_1_1_2_U40 ( .A1(npu_inst_int_data_res_2__2__6_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N79), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N71), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n78) );
  INV_X1 npu_inst_pe_1_1_2_U39 ( .A(npu_inst_pe_1_1_2_n78), .ZN(
        npu_inst_pe_1_1_2_n33) );
  AND2_X1 npu_inst_pe_1_1_2_U38 ( .A1(npu_inst_int_data_x_1__2__1_), .A2(
        npu_inst_pe_1_1_2_int_q_weight_1_), .ZN(npu_inst_pe_1_1_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_2_U37 ( .A1(npu_inst_int_data_x_1__2__0_), .A2(
        npu_inst_pe_1_1_2_int_q_weight_1_), .ZN(npu_inst_pe_1_1_2_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_1_2_U36 ( .A(npu_inst_pe_1_1_2_int_data_1_), .ZN(
        npu_inst_pe_1_1_2_n13) );
  NOR3_X1 npu_inst_pe_1_1_2_U35 ( .A1(npu_inst_pe_1_1_2_n26), .A2(npu_inst_n41), .A3(npu_inst_int_ckg[53]), .ZN(npu_inst_pe_1_1_2_n85) );
  OR2_X1 npu_inst_pe_1_1_2_U34 ( .A1(npu_inst_pe_1_1_2_n85), .A2(
        npu_inst_pe_1_1_2_n1), .ZN(npu_inst_pe_1_1_2_N84) );
  AOI222_X1 npu_inst_pe_1_1_2_U33 ( .A1(npu_inst_int_data_res_2__2__2_), .A2(
        npu_inst_pe_1_1_2_n1), .B1(npu_inst_pe_1_1_2_N75), .B2(
        npu_inst_pe_1_1_2_n76), .C1(npu_inst_pe_1_1_2_N67), .C2(
        npu_inst_pe_1_1_2_n77), .ZN(npu_inst_pe_1_1_2_n82) );
  INV_X1 npu_inst_pe_1_1_2_U32 ( .A(npu_inst_pe_1_1_2_n82), .ZN(
        npu_inst_pe_1_1_2_n98) );
  AOI22_X1 npu_inst_pe_1_1_2_U31 ( .A1(npu_inst_n41), .A2(
        npu_inst_int_data_y_2__2__1_), .B1(npu_inst_pe_1_1_2_n2), .B2(
        npu_inst_int_data_x_1__3__1_), .ZN(npu_inst_pe_1_1_2_n63) );
  AOI22_X1 npu_inst_pe_1_1_2_U30 ( .A1(npu_inst_n41), .A2(
        npu_inst_int_data_y_2__2__0_), .B1(npu_inst_pe_1_1_2_n2), .B2(
        npu_inst_int_data_x_1__3__0_), .ZN(npu_inst_pe_1_1_2_n61) );
  INV_X1 npu_inst_pe_1_1_2_U29 ( .A(npu_inst_pe_1_1_2_int_data_0_), .ZN(
        npu_inst_pe_1_1_2_n12) );
  INV_X1 npu_inst_pe_1_1_2_U28 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_1_2_n4)
         );
  OR3_X1 npu_inst_pe_1_1_2_U27 ( .A1(npu_inst_pe_1_1_2_n5), .A2(
        npu_inst_pe_1_1_2_n7), .A3(npu_inst_pe_1_1_2_n4), .ZN(
        npu_inst_pe_1_1_2_n56) );
  OR3_X1 npu_inst_pe_1_1_2_U26 ( .A1(npu_inst_pe_1_1_2_n4), .A2(
        npu_inst_pe_1_1_2_n7), .A3(npu_inst_pe_1_1_2_n6), .ZN(
        npu_inst_pe_1_1_2_n48) );
  INV_X1 npu_inst_pe_1_1_2_U25 ( .A(npu_inst_pe_1_1_2_n4), .ZN(
        npu_inst_pe_1_1_2_n3) );
  OR3_X1 npu_inst_pe_1_1_2_U24 ( .A1(npu_inst_pe_1_1_2_n3), .A2(
        npu_inst_pe_1_1_2_n7), .A3(npu_inst_pe_1_1_2_n6), .ZN(
        npu_inst_pe_1_1_2_n52) );
  OR3_X1 npu_inst_pe_1_1_2_U23 ( .A1(npu_inst_pe_1_1_2_n5), .A2(
        npu_inst_pe_1_1_2_n7), .A3(npu_inst_pe_1_1_2_n3), .ZN(
        npu_inst_pe_1_1_2_n60) );
  BUF_X1 npu_inst_pe_1_1_2_U22 ( .A(npu_inst_n28), .Z(npu_inst_pe_1_1_2_n1) );
  NOR2_X1 npu_inst_pe_1_1_2_U21 ( .A1(npu_inst_pe_1_1_2_n60), .A2(
        npu_inst_pe_1_1_2_n2), .ZN(npu_inst_pe_1_1_2_n58) );
  NOR2_X1 npu_inst_pe_1_1_2_U20 ( .A1(npu_inst_pe_1_1_2_n56), .A2(
        npu_inst_pe_1_1_2_n2), .ZN(npu_inst_pe_1_1_2_n54) );
  NOR2_X1 npu_inst_pe_1_1_2_U19 ( .A1(npu_inst_pe_1_1_2_n52), .A2(
        npu_inst_pe_1_1_2_n2), .ZN(npu_inst_pe_1_1_2_n50) );
  NOR2_X1 npu_inst_pe_1_1_2_U18 ( .A1(npu_inst_pe_1_1_2_n48), .A2(
        npu_inst_pe_1_1_2_n2), .ZN(npu_inst_pe_1_1_2_n46) );
  NOR2_X1 npu_inst_pe_1_1_2_U17 ( .A1(npu_inst_pe_1_1_2_n40), .A2(
        npu_inst_pe_1_1_2_n2), .ZN(npu_inst_pe_1_1_2_n38) );
  NOR2_X1 npu_inst_pe_1_1_2_U16 ( .A1(npu_inst_pe_1_1_2_n44), .A2(
        npu_inst_pe_1_1_2_n2), .ZN(npu_inst_pe_1_1_2_n42) );
  BUF_X1 npu_inst_pe_1_1_2_U15 ( .A(npu_inst_n87), .Z(npu_inst_pe_1_1_2_n7) );
  INV_X1 npu_inst_pe_1_1_2_U14 ( .A(npu_inst_n108), .ZN(npu_inst_pe_1_1_2_n11)
         );
  INV_X1 npu_inst_pe_1_1_2_U13 ( .A(npu_inst_pe_1_1_2_n38), .ZN(
        npu_inst_pe_1_1_2_n113) );
  INV_X1 npu_inst_pe_1_1_2_U12 ( .A(npu_inst_pe_1_1_2_n58), .ZN(
        npu_inst_pe_1_1_2_n118) );
  INV_X1 npu_inst_pe_1_1_2_U11 ( .A(npu_inst_pe_1_1_2_n54), .ZN(
        npu_inst_pe_1_1_2_n117) );
  INV_X1 npu_inst_pe_1_1_2_U10 ( .A(npu_inst_pe_1_1_2_n50), .ZN(
        npu_inst_pe_1_1_2_n116) );
  INV_X1 npu_inst_pe_1_1_2_U9 ( .A(npu_inst_pe_1_1_2_n46), .ZN(
        npu_inst_pe_1_1_2_n115) );
  INV_X1 npu_inst_pe_1_1_2_U8 ( .A(npu_inst_pe_1_1_2_n42), .ZN(
        npu_inst_pe_1_1_2_n114) );
  BUF_X1 npu_inst_pe_1_1_2_U7 ( .A(npu_inst_pe_1_1_2_n11), .Z(
        npu_inst_pe_1_1_2_n10) );
  BUF_X1 npu_inst_pe_1_1_2_U6 ( .A(npu_inst_pe_1_1_2_n11), .Z(
        npu_inst_pe_1_1_2_n9) );
  BUF_X1 npu_inst_pe_1_1_2_U5 ( .A(npu_inst_pe_1_1_2_n11), .Z(
        npu_inst_pe_1_1_2_n8) );
  NOR2_X1 npu_inst_pe_1_1_2_U4 ( .A1(npu_inst_pe_1_1_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_2_n1), .ZN(npu_inst_pe_1_1_2_n76) );
  NOR2_X1 npu_inst_pe_1_1_2_U3 ( .A1(npu_inst_pe_1_1_2_n27), .A2(
        npu_inst_pe_1_1_2_n1), .ZN(npu_inst_pe_1_1_2_n77) );
  FA_X1 npu_inst_pe_1_1_2_sub_77_U2_1 ( .A(npu_inst_int_data_res_1__2__1_), 
        .B(npu_inst_pe_1_1_2_n13), .CI(npu_inst_pe_1_1_2_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_1_2_sub_77_carry_2_), .S(npu_inst_pe_1_1_2_N66) );
  FA_X1 npu_inst_pe_1_1_2_add_79_U1_1 ( .A(npu_inst_int_data_res_1__2__1_), 
        .B(npu_inst_pe_1_1_2_int_data_1_), .CI(
        npu_inst_pe_1_1_2_add_79_carry_1_), .CO(
        npu_inst_pe_1_1_2_add_79_carry_2_), .S(npu_inst_pe_1_1_2_N74) );
  NAND3_X1 npu_inst_pe_1_1_2_U101 ( .A1(npu_inst_pe_1_1_2_n4), .A2(
        npu_inst_pe_1_1_2_n6), .A3(npu_inst_pe_1_1_2_n7), .ZN(
        npu_inst_pe_1_1_2_n44) );
  NAND3_X1 npu_inst_pe_1_1_2_U100 ( .A1(npu_inst_pe_1_1_2_n3), .A2(
        npu_inst_pe_1_1_2_n6), .A3(npu_inst_pe_1_1_2_n7), .ZN(
        npu_inst_pe_1_1_2_n40) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_2_n33), .CK(
        npu_inst_pe_1_1_2_net4248), .RN(npu_inst_pe_1_1_2_n8), .Q(
        npu_inst_int_data_res_1__2__6_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_2_n34), .CK(
        npu_inst_pe_1_1_2_net4248), .RN(npu_inst_pe_1_1_2_n8), .Q(
        npu_inst_int_data_res_1__2__5_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_2_n35), .CK(
        npu_inst_pe_1_1_2_net4248), .RN(npu_inst_pe_1_1_2_n8), .Q(
        npu_inst_int_data_res_1__2__4_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_2_n36), .CK(
        npu_inst_pe_1_1_2_net4248), .RN(npu_inst_pe_1_1_2_n8), .Q(
        npu_inst_int_data_res_1__2__3_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_2_n98), .CK(
        npu_inst_pe_1_1_2_net4248), .RN(npu_inst_pe_1_1_2_n8), .Q(
        npu_inst_int_data_res_1__2__2_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_2_n99), .CK(
        npu_inst_pe_1_1_2_net4248), .RN(npu_inst_pe_1_1_2_n8), .Q(
        npu_inst_int_data_res_1__2__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_2_n32), .CK(
        npu_inst_pe_1_1_2_net4248), .RN(npu_inst_pe_1_1_2_n8), .Q(
        npu_inst_int_data_res_1__2__7_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_2_n100), 
        .CK(npu_inst_pe_1_1_2_net4248), .RN(npu_inst_pe_1_1_2_n8), .Q(
        npu_inst_int_data_res_1__2__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_weight_reg_0_ ( .D(npu_inst_n94), .CK(
        npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n8), .Q(
        npu_inst_pe_1_1_2_int_q_weight_0_), .QN(npu_inst_pe_1_1_2_n27) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_weight_reg_1_ ( .D(npu_inst_n100), .CK(
        npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n8), .Q(
        npu_inst_pe_1_1_2_int_q_weight_1_), .QN(npu_inst_pe_1_1_2_n26) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_2_n112), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n8), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_2_n106), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n8), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_2_n111), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_2_n105), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_2_n110), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_2_n104), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_2_n109), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_2_n103), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_2_n108), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_2_n102), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_2_n107), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_2_n101), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_2_n86), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_2_n87), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n9), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_2_n88), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_2_n89), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_2_n90), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_2_n91), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_2_n92), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_2_n93), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_2_n94), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_2_n95), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_2_n96), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_2_n97), 
        .CK(npu_inst_pe_1_1_2_net4254), .RN(npu_inst_pe_1_1_2_n10), .Q(
        npu_inst_pe_1_1_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_2_net4248) );
  CLKGATETST_X1 npu_inst_pe_1_1_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n47), .SE(1'b0), .GCK(npu_inst_pe_1_1_2_net4254) );
  MUX2_X1 npu_inst_pe_1_1_3_U153 ( .A(npu_inst_pe_1_1_3_n31), .B(
        npu_inst_pe_1_1_3_n28), .S(npu_inst_pe_1_1_3_n7), .Z(
        npu_inst_pe_1_1_3_N93) );
  MUX2_X1 npu_inst_pe_1_1_3_U152 ( .A(npu_inst_pe_1_1_3_n30), .B(
        npu_inst_pe_1_1_3_n29), .S(npu_inst_pe_1_1_3_n5), .Z(
        npu_inst_pe_1_1_3_n31) );
  MUX2_X1 npu_inst_pe_1_1_3_U151 ( .A(npu_inst_pe_1_1_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_3_n3), .Z(
        npu_inst_pe_1_1_3_n30) );
  MUX2_X1 npu_inst_pe_1_1_3_U150 ( .A(npu_inst_pe_1_1_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_3_n3), .Z(
        npu_inst_pe_1_1_3_n29) );
  MUX2_X1 npu_inst_pe_1_1_3_U149 ( .A(npu_inst_pe_1_1_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_3_n3), .Z(
        npu_inst_pe_1_1_3_n28) );
  MUX2_X1 npu_inst_pe_1_1_3_U148 ( .A(npu_inst_pe_1_1_3_n25), .B(
        npu_inst_pe_1_1_3_n22), .S(npu_inst_pe_1_1_3_n7), .Z(
        npu_inst_pe_1_1_3_N94) );
  MUX2_X1 npu_inst_pe_1_1_3_U147 ( .A(npu_inst_pe_1_1_3_n24), .B(
        npu_inst_pe_1_1_3_n23), .S(npu_inst_pe_1_1_3_n5), .Z(
        npu_inst_pe_1_1_3_n25) );
  MUX2_X1 npu_inst_pe_1_1_3_U146 ( .A(npu_inst_pe_1_1_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_3_n3), .Z(
        npu_inst_pe_1_1_3_n24) );
  MUX2_X1 npu_inst_pe_1_1_3_U145 ( .A(npu_inst_pe_1_1_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_3_n3), .Z(
        npu_inst_pe_1_1_3_n23) );
  MUX2_X1 npu_inst_pe_1_1_3_U144 ( .A(npu_inst_pe_1_1_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_3_n3), .Z(
        npu_inst_pe_1_1_3_n22) );
  MUX2_X1 npu_inst_pe_1_1_3_U143 ( .A(npu_inst_pe_1_1_3_n21), .B(
        npu_inst_pe_1_1_3_n18), .S(npu_inst_pe_1_1_3_n7), .Z(
        npu_inst_int_data_x_1__3__1_) );
  MUX2_X1 npu_inst_pe_1_1_3_U142 ( .A(npu_inst_pe_1_1_3_n20), .B(
        npu_inst_pe_1_1_3_n19), .S(npu_inst_pe_1_1_3_n5), .Z(
        npu_inst_pe_1_1_3_n21) );
  MUX2_X1 npu_inst_pe_1_1_3_U141 ( .A(npu_inst_pe_1_1_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_3_n3), .Z(
        npu_inst_pe_1_1_3_n20) );
  MUX2_X1 npu_inst_pe_1_1_3_U140 ( .A(npu_inst_pe_1_1_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_3_n3), .Z(
        npu_inst_pe_1_1_3_n19) );
  MUX2_X1 npu_inst_pe_1_1_3_U139 ( .A(npu_inst_pe_1_1_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_3_n3), .Z(
        npu_inst_pe_1_1_3_n18) );
  MUX2_X1 npu_inst_pe_1_1_3_U138 ( .A(npu_inst_pe_1_1_3_n17), .B(
        npu_inst_pe_1_1_3_n14), .S(npu_inst_pe_1_1_3_n7), .Z(
        npu_inst_int_data_x_1__3__0_) );
  MUX2_X1 npu_inst_pe_1_1_3_U137 ( .A(npu_inst_pe_1_1_3_n16), .B(
        npu_inst_pe_1_1_3_n15), .S(npu_inst_pe_1_1_3_n5), .Z(
        npu_inst_pe_1_1_3_n17) );
  MUX2_X1 npu_inst_pe_1_1_3_U136 ( .A(npu_inst_pe_1_1_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_3_n3), .Z(
        npu_inst_pe_1_1_3_n16) );
  MUX2_X1 npu_inst_pe_1_1_3_U135 ( .A(npu_inst_pe_1_1_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_3_n3), .Z(
        npu_inst_pe_1_1_3_n15) );
  MUX2_X1 npu_inst_pe_1_1_3_U134 ( .A(npu_inst_pe_1_1_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_3_n3), .Z(
        npu_inst_pe_1_1_3_n14) );
  XOR2_X1 npu_inst_pe_1_1_3_U133 ( .A(npu_inst_pe_1_1_3_int_data_0_), .B(
        npu_inst_int_data_res_1__3__0_), .Z(npu_inst_pe_1_1_3_N73) );
  AND2_X1 npu_inst_pe_1_1_3_U132 ( .A1(npu_inst_int_data_res_1__3__0_), .A2(
        npu_inst_pe_1_1_3_int_data_0_), .ZN(npu_inst_pe_1_1_3_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_3_U131 ( .A(npu_inst_int_data_res_1__3__0_), .B(
        npu_inst_pe_1_1_3_n12), .ZN(npu_inst_pe_1_1_3_N65) );
  OR2_X1 npu_inst_pe_1_1_3_U130 ( .A1(npu_inst_pe_1_1_3_n12), .A2(
        npu_inst_int_data_res_1__3__0_), .ZN(npu_inst_pe_1_1_3_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_3_U129 ( .A(npu_inst_int_data_res_1__3__2_), .B(
        npu_inst_pe_1_1_3_add_79_carry_2_), .Z(npu_inst_pe_1_1_3_N75) );
  AND2_X1 npu_inst_pe_1_1_3_U128 ( .A1(npu_inst_pe_1_1_3_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_1__3__2_), .ZN(
        npu_inst_pe_1_1_3_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_3_U127 ( .A(npu_inst_int_data_res_1__3__3_), .B(
        npu_inst_pe_1_1_3_add_79_carry_3_), .Z(npu_inst_pe_1_1_3_N76) );
  AND2_X1 npu_inst_pe_1_1_3_U126 ( .A1(npu_inst_pe_1_1_3_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_1__3__3_), .ZN(
        npu_inst_pe_1_1_3_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_3_U125 ( .A(npu_inst_int_data_res_1__3__4_), .B(
        npu_inst_pe_1_1_3_add_79_carry_4_), .Z(npu_inst_pe_1_1_3_N77) );
  AND2_X1 npu_inst_pe_1_1_3_U124 ( .A1(npu_inst_pe_1_1_3_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_1__3__4_), .ZN(
        npu_inst_pe_1_1_3_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_3_U123 ( .A(npu_inst_int_data_res_1__3__5_), .B(
        npu_inst_pe_1_1_3_add_79_carry_5_), .Z(npu_inst_pe_1_1_3_N78) );
  AND2_X1 npu_inst_pe_1_1_3_U122 ( .A1(npu_inst_pe_1_1_3_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_1__3__5_), .ZN(
        npu_inst_pe_1_1_3_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_3_U121 ( .A(npu_inst_int_data_res_1__3__6_), .B(
        npu_inst_pe_1_1_3_add_79_carry_6_), .Z(npu_inst_pe_1_1_3_N79) );
  AND2_X1 npu_inst_pe_1_1_3_U120 ( .A1(npu_inst_pe_1_1_3_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_1__3__6_), .ZN(
        npu_inst_pe_1_1_3_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_3_U119 ( .A(npu_inst_int_data_res_1__3__7_), .B(
        npu_inst_pe_1_1_3_add_79_carry_7_), .Z(npu_inst_pe_1_1_3_N80) );
  XNOR2_X1 npu_inst_pe_1_1_3_U118 ( .A(npu_inst_pe_1_1_3_sub_77_carry_2_), .B(
        npu_inst_int_data_res_1__3__2_), .ZN(npu_inst_pe_1_1_3_N67) );
  OR2_X1 npu_inst_pe_1_1_3_U117 ( .A1(npu_inst_int_data_res_1__3__2_), .A2(
        npu_inst_pe_1_1_3_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_1_3_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_3_U116 ( .A(npu_inst_pe_1_1_3_sub_77_carry_3_), .B(
        npu_inst_int_data_res_1__3__3_), .ZN(npu_inst_pe_1_1_3_N68) );
  OR2_X1 npu_inst_pe_1_1_3_U115 ( .A1(npu_inst_int_data_res_1__3__3_), .A2(
        npu_inst_pe_1_1_3_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_1_3_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_3_U114 ( .A(npu_inst_pe_1_1_3_sub_77_carry_4_), .B(
        npu_inst_int_data_res_1__3__4_), .ZN(npu_inst_pe_1_1_3_N69) );
  OR2_X1 npu_inst_pe_1_1_3_U113 ( .A1(npu_inst_int_data_res_1__3__4_), .A2(
        npu_inst_pe_1_1_3_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_1_3_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_3_U112 ( .A(npu_inst_pe_1_1_3_sub_77_carry_5_), .B(
        npu_inst_int_data_res_1__3__5_), .ZN(npu_inst_pe_1_1_3_N70) );
  OR2_X1 npu_inst_pe_1_1_3_U111 ( .A1(npu_inst_int_data_res_1__3__5_), .A2(
        npu_inst_pe_1_1_3_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_1_3_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_3_U110 ( .A(npu_inst_pe_1_1_3_sub_77_carry_6_), .B(
        npu_inst_int_data_res_1__3__6_), .ZN(npu_inst_pe_1_1_3_N71) );
  OR2_X1 npu_inst_pe_1_1_3_U109 ( .A1(npu_inst_int_data_res_1__3__6_), .A2(
        npu_inst_pe_1_1_3_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_1_3_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_3_U108 ( .A(npu_inst_int_data_res_1__3__7_), .B(
        npu_inst_pe_1_1_3_sub_77_carry_7_), .ZN(npu_inst_pe_1_1_3_N72) );
  INV_X1 npu_inst_pe_1_1_3_U107 ( .A(npu_inst_n61), .ZN(npu_inst_pe_1_1_3_n6)
         );
  INV_X1 npu_inst_pe_1_1_3_U106 ( .A(npu_inst_pe_1_1_3_n6), .ZN(
        npu_inst_pe_1_1_3_n5) );
  INV_X1 npu_inst_pe_1_1_3_U105 ( .A(npu_inst_n41), .ZN(npu_inst_pe_1_1_3_n2)
         );
  AOI22_X1 npu_inst_pe_1_1_3_U104 ( .A1(npu_inst_int_data_y_2__3__0_), .A2(
        npu_inst_pe_1_1_3_n58), .B1(npu_inst_pe_1_1_3_n118), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_3_n57) );
  INV_X1 npu_inst_pe_1_1_3_U103 ( .A(npu_inst_pe_1_1_3_n57), .ZN(
        npu_inst_pe_1_1_3_n107) );
  AOI22_X1 npu_inst_pe_1_1_3_U102 ( .A1(npu_inst_int_data_y_2__3__0_), .A2(
        npu_inst_pe_1_1_3_n54), .B1(npu_inst_pe_1_1_3_n117), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_3_n53) );
  INV_X1 npu_inst_pe_1_1_3_U99 ( .A(npu_inst_pe_1_1_3_n53), .ZN(
        npu_inst_pe_1_1_3_n108) );
  AOI22_X1 npu_inst_pe_1_1_3_U98 ( .A1(npu_inst_int_data_y_2__3__0_), .A2(
        npu_inst_pe_1_1_3_n50), .B1(npu_inst_pe_1_1_3_n116), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_3_n49) );
  INV_X1 npu_inst_pe_1_1_3_U97 ( .A(npu_inst_pe_1_1_3_n49), .ZN(
        npu_inst_pe_1_1_3_n109) );
  AOI22_X1 npu_inst_pe_1_1_3_U96 ( .A1(npu_inst_int_data_y_2__3__0_), .A2(
        npu_inst_pe_1_1_3_n46), .B1(npu_inst_pe_1_1_3_n115), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_3_n45) );
  INV_X1 npu_inst_pe_1_1_3_U95 ( .A(npu_inst_pe_1_1_3_n45), .ZN(
        npu_inst_pe_1_1_3_n110) );
  AOI22_X1 npu_inst_pe_1_1_3_U94 ( .A1(npu_inst_int_data_y_2__3__0_), .A2(
        npu_inst_pe_1_1_3_n42), .B1(npu_inst_pe_1_1_3_n114), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_3_n41) );
  INV_X1 npu_inst_pe_1_1_3_U93 ( .A(npu_inst_pe_1_1_3_n41), .ZN(
        npu_inst_pe_1_1_3_n111) );
  AOI22_X1 npu_inst_pe_1_1_3_U92 ( .A1(npu_inst_int_data_y_2__3__1_), .A2(
        npu_inst_pe_1_1_3_n58), .B1(npu_inst_pe_1_1_3_n118), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_3_n59) );
  INV_X1 npu_inst_pe_1_1_3_U91 ( .A(npu_inst_pe_1_1_3_n59), .ZN(
        npu_inst_pe_1_1_3_n101) );
  AOI22_X1 npu_inst_pe_1_1_3_U90 ( .A1(npu_inst_int_data_y_2__3__1_), .A2(
        npu_inst_pe_1_1_3_n54), .B1(npu_inst_pe_1_1_3_n117), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_3_n55) );
  INV_X1 npu_inst_pe_1_1_3_U89 ( .A(npu_inst_pe_1_1_3_n55), .ZN(
        npu_inst_pe_1_1_3_n102) );
  AOI22_X1 npu_inst_pe_1_1_3_U88 ( .A1(npu_inst_int_data_y_2__3__1_), .A2(
        npu_inst_pe_1_1_3_n50), .B1(npu_inst_pe_1_1_3_n116), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_3_n51) );
  INV_X1 npu_inst_pe_1_1_3_U87 ( .A(npu_inst_pe_1_1_3_n51), .ZN(
        npu_inst_pe_1_1_3_n103) );
  AOI22_X1 npu_inst_pe_1_1_3_U86 ( .A1(npu_inst_int_data_y_2__3__1_), .A2(
        npu_inst_pe_1_1_3_n46), .B1(npu_inst_pe_1_1_3_n115), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_3_n47) );
  INV_X1 npu_inst_pe_1_1_3_U85 ( .A(npu_inst_pe_1_1_3_n47), .ZN(
        npu_inst_pe_1_1_3_n104) );
  AOI22_X1 npu_inst_pe_1_1_3_U84 ( .A1(npu_inst_int_data_y_2__3__1_), .A2(
        npu_inst_pe_1_1_3_n42), .B1(npu_inst_pe_1_1_3_n114), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_3_n43) );
  INV_X1 npu_inst_pe_1_1_3_U83 ( .A(npu_inst_pe_1_1_3_n43), .ZN(
        npu_inst_pe_1_1_3_n105) );
  AOI22_X1 npu_inst_pe_1_1_3_U82 ( .A1(npu_inst_pe_1_1_3_n38), .A2(
        npu_inst_int_data_y_2__3__1_), .B1(npu_inst_pe_1_1_3_n113), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_3_n39) );
  INV_X1 npu_inst_pe_1_1_3_U81 ( .A(npu_inst_pe_1_1_3_n39), .ZN(
        npu_inst_pe_1_1_3_n106) );
  AND2_X1 npu_inst_pe_1_1_3_U80 ( .A1(npu_inst_pe_1_1_3_N93), .A2(npu_inst_n41), .ZN(npu_inst_int_data_y_1__3__0_) );
  NAND2_X1 npu_inst_pe_1_1_3_U79 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_3_n60), .ZN(npu_inst_pe_1_1_3_n74) );
  OAI21_X1 npu_inst_pe_1_1_3_U78 ( .B1(npu_inst_pe_1_1_3_n63), .B2(
        npu_inst_pe_1_1_3_n60), .A(npu_inst_pe_1_1_3_n74), .ZN(
        npu_inst_pe_1_1_3_n97) );
  NAND2_X1 npu_inst_pe_1_1_3_U77 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_3_n60), .ZN(npu_inst_pe_1_1_3_n73) );
  OAI21_X1 npu_inst_pe_1_1_3_U76 ( .B1(npu_inst_pe_1_1_3_n61), .B2(
        npu_inst_pe_1_1_3_n60), .A(npu_inst_pe_1_1_3_n73), .ZN(
        npu_inst_pe_1_1_3_n96) );
  NAND2_X1 npu_inst_pe_1_1_3_U75 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_3_n56), .ZN(npu_inst_pe_1_1_3_n72) );
  OAI21_X1 npu_inst_pe_1_1_3_U74 ( .B1(npu_inst_pe_1_1_3_n63), .B2(
        npu_inst_pe_1_1_3_n56), .A(npu_inst_pe_1_1_3_n72), .ZN(
        npu_inst_pe_1_1_3_n95) );
  NAND2_X1 npu_inst_pe_1_1_3_U73 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_3_n56), .ZN(npu_inst_pe_1_1_3_n71) );
  OAI21_X1 npu_inst_pe_1_1_3_U72 ( .B1(npu_inst_pe_1_1_3_n61), .B2(
        npu_inst_pe_1_1_3_n56), .A(npu_inst_pe_1_1_3_n71), .ZN(
        npu_inst_pe_1_1_3_n94) );
  NAND2_X1 npu_inst_pe_1_1_3_U71 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_3_n52), .ZN(npu_inst_pe_1_1_3_n70) );
  OAI21_X1 npu_inst_pe_1_1_3_U70 ( .B1(npu_inst_pe_1_1_3_n63), .B2(
        npu_inst_pe_1_1_3_n52), .A(npu_inst_pe_1_1_3_n70), .ZN(
        npu_inst_pe_1_1_3_n93) );
  NAND2_X1 npu_inst_pe_1_1_3_U69 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_3_n52), .ZN(npu_inst_pe_1_1_3_n69) );
  OAI21_X1 npu_inst_pe_1_1_3_U68 ( .B1(npu_inst_pe_1_1_3_n61), .B2(
        npu_inst_pe_1_1_3_n52), .A(npu_inst_pe_1_1_3_n69), .ZN(
        npu_inst_pe_1_1_3_n92) );
  NAND2_X1 npu_inst_pe_1_1_3_U67 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_3_n48), .ZN(npu_inst_pe_1_1_3_n68) );
  OAI21_X1 npu_inst_pe_1_1_3_U66 ( .B1(npu_inst_pe_1_1_3_n63), .B2(
        npu_inst_pe_1_1_3_n48), .A(npu_inst_pe_1_1_3_n68), .ZN(
        npu_inst_pe_1_1_3_n91) );
  NAND2_X1 npu_inst_pe_1_1_3_U65 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_3_n48), .ZN(npu_inst_pe_1_1_3_n67) );
  OAI21_X1 npu_inst_pe_1_1_3_U64 ( .B1(npu_inst_pe_1_1_3_n61), .B2(
        npu_inst_pe_1_1_3_n48), .A(npu_inst_pe_1_1_3_n67), .ZN(
        npu_inst_pe_1_1_3_n90) );
  NAND2_X1 npu_inst_pe_1_1_3_U63 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_3_n44), .ZN(npu_inst_pe_1_1_3_n66) );
  OAI21_X1 npu_inst_pe_1_1_3_U62 ( .B1(npu_inst_pe_1_1_3_n63), .B2(
        npu_inst_pe_1_1_3_n44), .A(npu_inst_pe_1_1_3_n66), .ZN(
        npu_inst_pe_1_1_3_n89) );
  NAND2_X1 npu_inst_pe_1_1_3_U61 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_3_n44), .ZN(npu_inst_pe_1_1_3_n65) );
  OAI21_X1 npu_inst_pe_1_1_3_U60 ( .B1(npu_inst_pe_1_1_3_n61), .B2(
        npu_inst_pe_1_1_3_n44), .A(npu_inst_pe_1_1_3_n65), .ZN(
        npu_inst_pe_1_1_3_n88) );
  NAND2_X1 npu_inst_pe_1_1_3_U59 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_3_n40), .ZN(npu_inst_pe_1_1_3_n64) );
  OAI21_X1 npu_inst_pe_1_1_3_U58 ( .B1(npu_inst_pe_1_1_3_n63), .B2(
        npu_inst_pe_1_1_3_n40), .A(npu_inst_pe_1_1_3_n64), .ZN(
        npu_inst_pe_1_1_3_n87) );
  NAND2_X1 npu_inst_pe_1_1_3_U57 ( .A1(npu_inst_pe_1_1_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_3_n40), .ZN(npu_inst_pe_1_1_3_n62) );
  OAI21_X1 npu_inst_pe_1_1_3_U56 ( .B1(npu_inst_pe_1_1_3_n61), .B2(
        npu_inst_pe_1_1_3_n40), .A(npu_inst_pe_1_1_3_n62), .ZN(
        npu_inst_pe_1_1_3_n86) );
  AOI22_X1 npu_inst_pe_1_1_3_U55 ( .A1(npu_inst_pe_1_1_3_n38), .A2(
        npu_inst_int_data_y_2__3__0_), .B1(npu_inst_pe_1_1_3_n113), .B2(
        npu_inst_pe_1_1_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_3_n37) );
  INV_X1 npu_inst_pe_1_1_3_U54 ( .A(npu_inst_pe_1_1_3_n37), .ZN(
        npu_inst_pe_1_1_3_n112) );
  AND2_X1 npu_inst_pe_1_1_3_U53 ( .A1(npu_inst_n41), .A2(npu_inst_pe_1_1_3_N94), .ZN(npu_inst_int_data_y_1__3__1_) );
  AOI222_X1 npu_inst_pe_1_1_3_U52 ( .A1(npu_inst_int_data_res_2__3__0_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N73), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N65), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n84) );
  INV_X1 npu_inst_pe_1_1_3_U51 ( .A(npu_inst_pe_1_1_3_n84), .ZN(
        npu_inst_pe_1_1_3_n100) );
  AOI222_X1 npu_inst_pe_1_1_3_U50 ( .A1(npu_inst_pe_1_1_3_n1), .A2(
        npu_inst_int_data_res_2__3__7_), .B1(npu_inst_pe_1_1_3_N80), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N72), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n75) );
  INV_X1 npu_inst_pe_1_1_3_U49 ( .A(npu_inst_pe_1_1_3_n75), .ZN(
        npu_inst_pe_1_1_3_n32) );
  AOI222_X1 npu_inst_pe_1_1_3_U48 ( .A1(npu_inst_int_data_res_2__3__1_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N74), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N66), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n83) );
  INV_X1 npu_inst_pe_1_1_3_U47 ( .A(npu_inst_pe_1_1_3_n83), .ZN(
        npu_inst_pe_1_1_3_n99) );
  AOI222_X1 npu_inst_pe_1_1_3_U46 ( .A1(npu_inst_int_data_res_2__3__3_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N76), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N68), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n81) );
  INV_X1 npu_inst_pe_1_1_3_U45 ( .A(npu_inst_pe_1_1_3_n81), .ZN(
        npu_inst_pe_1_1_3_n36) );
  AOI222_X1 npu_inst_pe_1_1_3_U44 ( .A1(npu_inst_int_data_res_2__3__4_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N77), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N69), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n80) );
  INV_X1 npu_inst_pe_1_1_3_U43 ( .A(npu_inst_pe_1_1_3_n80), .ZN(
        npu_inst_pe_1_1_3_n35) );
  AOI222_X1 npu_inst_pe_1_1_3_U42 ( .A1(npu_inst_int_data_res_2__3__5_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N78), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N70), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n79) );
  INV_X1 npu_inst_pe_1_1_3_U41 ( .A(npu_inst_pe_1_1_3_n79), .ZN(
        npu_inst_pe_1_1_3_n34) );
  AOI222_X1 npu_inst_pe_1_1_3_U40 ( .A1(npu_inst_int_data_res_2__3__6_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N79), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N71), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n78) );
  INV_X1 npu_inst_pe_1_1_3_U39 ( .A(npu_inst_pe_1_1_3_n78), .ZN(
        npu_inst_pe_1_1_3_n33) );
  AND2_X1 npu_inst_pe_1_1_3_U38 ( .A1(npu_inst_int_data_x_1__3__1_), .A2(
        npu_inst_pe_1_1_3_int_q_weight_1_), .ZN(npu_inst_pe_1_1_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_3_U37 ( .A1(npu_inst_int_data_x_1__3__0_), .A2(
        npu_inst_pe_1_1_3_int_q_weight_1_), .ZN(npu_inst_pe_1_1_3_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_1_3_U36 ( .A(npu_inst_pe_1_1_3_int_data_1_), .ZN(
        npu_inst_pe_1_1_3_n13) );
  NOR3_X1 npu_inst_pe_1_1_3_U35 ( .A1(npu_inst_pe_1_1_3_n26), .A2(npu_inst_n41), .A3(npu_inst_int_ckg[52]), .ZN(npu_inst_pe_1_1_3_n85) );
  OR2_X1 npu_inst_pe_1_1_3_U34 ( .A1(npu_inst_pe_1_1_3_n85), .A2(
        npu_inst_pe_1_1_3_n1), .ZN(npu_inst_pe_1_1_3_N84) );
  AOI222_X1 npu_inst_pe_1_1_3_U33 ( .A1(npu_inst_int_data_res_2__3__2_), .A2(
        npu_inst_pe_1_1_3_n1), .B1(npu_inst_pe_1_1_3_N75), .B2(
        npu_inst_pe_1_1_3_n76), .C1(npu_inst_pe_1_1_3_N67), .C2(
        npu_inst_pe_1_1_3_n77), .ZN(npu_inst_pe_1_1_3_n82) );
  INV_X1 npu_inst_pe_1_1_3_U32 ( .A(npu_inst_pe_1_1_3_n82), .ZN(
        npu_inst_pe_1_1_3_n98) );
  AOI22_X1 npu_inst_pe_1_1_3_U31 ( .A1(npu_inst_n41), .A2(
        npu_inst_int_data_y_2__3__1_), .B1(npu_inst_pe_1_1_3_n2), .B2(
        npu_inst_int_data_x_1__4__1_), .ZN(npu_inst_pe_1_1_3_n63) );
  AOI22_X1 npu_inst_pe_1_1_3_U30 ( .A1(npu_inst_n41), .A2(
        npu_inst_int_data_y_2__3__0_), .B1(npu_inst_pe_1_1_3_n2), .B2(
        npu_inst_int_data_x_1__4__0_), .ZN(npu_inst_pe_1_1_3_n61) );
  INV_X1 npu_inst_pe_1_1_3_U29 ( .A(npu_inst_pe_1_1_3_int_data_0_), .ZN(
        npu_inst_pe_1_1_3_n12) );
  INV_X1 npu_inst_pe_1_1_3_U28 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_1_3_n4)
         );
  OR3_X1 npu_inst_pe_1_1_3_U27 ( .A1(npu_inst_pe_1_1_3_n5), .A2(
        npu_inst_pe_1_1_3_n7), .A3(npu_inst_pe_1_1_3_n4), .ZN(
        npu_inst_pe_1_1_3_n56) );
  OR3_X1 npu_inst_pe_1_1_3_U26 ( .A1(npu_inst_pe_1_1_3_n4), .A2(
        npu_inst_pe_1_1_3_n7), .A3(npu_inst_pe_1_1_3_n6), .ZN(
        npu_inst_pe_1_1_3_n48) );
  INV_X1 npu_inst_pe_1_1_3_U25 ( .A(npu_inst_pe_1_1_3_n4), .ZN(
        npu_inst_pe_1_1_3_n3) );
  OR3_X1 npu_inst_pe_1_1_3_U24 ( .A1(npu_inst_pe_1_1_3_n3), .A2(
        npu_inst_pe_1_1_3_n7), .A3(npu_inst_pe_1_1_3_n6), .ZN(
        npu_inst_pe_1_1_3_n52) );
  OR3_X1 npu_inst_pe_1_1_3_U23 ( .A1(npu_inst_pe_1_1_3_n5), .A2(
        npu_inst_pe_1_1_3_n7), .A3(npu_inst_pe_1_1_3_n3), .ZN(
        npu_inst_pe_1_1_3_n60) );
  BUF_X1 npu_inst_pe_1_1_3_U22 ( .A(npu_inst_n28), .Z(npu_inst_pe_1_1_3_n1) );
  NOR2_X1 npu_inst_pe_1_1_3_U21 ( .A1(npu_inst_pe_1_1_3_n60), .A2(
        npu_inst_pe_1_1_3_n2), .ZN(npu_inst_pe_1_1_3_n58) );
  NOR2_X1 npu_inst_pe_1_1_3_U20 ( .A1(npu_inst_pe_1_1_3_n56), .A2(
        npu_inst_pe_1_1_3_n2), .ZN(npu_inst_pe_1_1_3_n54) );
  NOR2_X1 npu_inst_pe_1_1_3_U19 ( .A1(npu_inst_pe_1_1_3_n52), .A2(
        npu_inst_pe_1_1_3_n2), .ZN(npu_inst_pe_1_1_3_n50) );
  NOR2_X1 npu_inst_pe_1_1_3_U18 ( .A1(npu_inst_pe_1_1_3_n48), .A2(
        npu_inst_pe_1_1_3_n2), .ZN(npu_inst_pe_1_1_3_n46) );
  NOR2_X1 npu_inst_pe_1_1_3_U17 ( .A1(npu_inst_pe_1_1_3_n40), .A2(
        npu_inst_pe_1_1_3_n2), .ZN(npu_inst_pe_1_1_3_n38) );
  NOR2_X1 npu_inst_pe_1_1_3_U16 ( .A1(npu_inst_pe_1_1_3_n44), .A2(
        npu_inst_pe_1_1_3_n2), .ZN(npu_inst_pe_1_1_3_n42) );
  BUF_X1 npu_inst_pe_1_1_3_U15 ( .A(npu_inst_n87), .Z(npu_inst_pe_1_1_3_n7) );
  INV_X1 npu_inst_pe_1_1_3_U14 ( .A(npu_inst_n108), .ZN(npu_inst_pe_1_1_3_n11)
         );
  INV_X1 npu_inst_pe_1_1_3_U13 ( .A(npu_inst_pe_1_1_3_n38), .ZN(
        npu_inst_pe_1_1_3_n113) );
  INV_X1 npu_inst_pe_1_1_3_U12 ( .A(npu_inst_pe_1_1_3_n58), .ZN(
        npu_inst_pe_1_1_3_n118) );
  INV_X1 npu_inst_pe_1_1_3_U11 ( .A(npu_inst_pe_1_1_3_n54), .ZN(
        npu_inst_pe_1_1_3_n117) );
  INV_X1 npu_inst_pe_1_1_3_U10 ( .A(npu_inst_pe_1_1_3_n50), .ZN(
        npu_inst_pe_1_1_3_n116) );
  INV_X1 npu_inst_pe_1_1_3_U9 ( .A(npu_inst_pe_1_1_3_n46), .ZN(
        npu_inst_pe_1_1_3_n115) );
  INV_X1 npu_inst_pe_1_1_3_U8 ( .A(npu_inst_pe_1_1_3_n42), .ZN(
        npu_inst_pe_1_1_3_n114) );
  BUF_X1 npu_inst_pe_1_1_3_U7 ( .A(npu_inst_pe_1_1_3_n11), .Z(
        npu_inst_pe_1_1_3_n10) );
  BUF_X1 npu_inst_pe_1_1_3_U6 ( .A(npu_inst_pe_1_1_3_n11), .Z(
        npu_inst_pe_1_1_3_n9) );
  BUF_X1 npu_inst_pe_1_1_3_U5 ( .A(npu_inst_pe_1_1_3_n11), .Z(
        npu_inst_pe_1_1_3_n8) );
  NOR2_X1 npu_inst_pe_1_1_3_U4 ( .A1(npu_inst_pe_1_1_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_3_n1), .ZN(npu_inst_pe_1_1_3_n76) );
  NOR2_X1 npu_inst_pe_1_1_3_U3 ( .A1(npu_inst_pe_1_1_3_n27), .A2(
        npu_inst_pe_1_1_3_n1), .ZN(npu_inst_pe_1_1_3_n77) );
  FA_X1 npu_inst_pe_1_1_3_sub_77_U2_1 ( .A(npu_inst_int_data_res_1__3__1_), 
        .B(npu_inst_pe_1_1_3_n13), .CI(npu_inst_pe_1_1_3_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_1_3_sub_77_carry_2_), .S(npu_inst_pe_1_1_3_N66) );
  FA_X1 npu_inst_pe_1_1_3_add_79_U1_1 ( .A(npu_inst_int_data_res_1__3__1_), 
        .B(npu_inst_pe_1_1_3_int_data_1_), .CI(
        npu_inst_pe_1_1_3_add_79_carry_1_), .CO(
        npu_inst_pe_1_1_3_add_79_carry_2_), .S(npu_inst_pe_1_1_3_N74) );
  NAND3_X1 npu_inst_pe_1_1_3_U101 ( .A1(npu_inst_pe_1_1_3_n4), .A2(
        npu_inst_pe_1_1_3_n6), .A3(npu_inst_pe_1_1_3_n7), .ZN(
        npu_inst_pe_1_1_3_n44) );
  NAND3_X1 npu_inst_pe_1_1_3_U100 ( .A1(npu_inst_pe_1_1_3_n3), .A2(
        npu_inst_pe_1_1_3_n6), .A3(npu_inst_pe_1_1_3_n7), .ZN(
        npu_inst_pe_1_1_3_n40) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_3_n33), .CK(
        npu_inst_pe_1_1_3_net4225), .RN(npu_inst_pe_1_1_3_n8), .Q(
        npu_inst_int_data_res_1__3__6_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_3_n34), .CK(
        npu_inst_pe_1_1_3_net4225), .RN(npu_inst_pe_1_1_3_n8), .Q(
        npu_inst_int_data_res_1__3__5_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_3_n35), .CK(
        npu_inst_pe_1_1_3_net4225), .RN(npu_inst_pe_1_1_3_n8), .Q(
        npu_inst_int_data_res_1__3__4_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_3_n36), .CK(
        npu_inst_pe_1_1_3_net4225), .RN(npu_inst_pe_1_1_3_n8), .Q(
        npu_inst_int_data_res_1__3__3_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_3_n98), .CK(
        npu_inst_pe_1_1_3_net4225), .RN(npu_inst_pe_1_1_3_n8), .Q(
        npu_inst_int_data_res_1__3__2_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_3_n99), .CK(
        npu_inst_pe_1_1_3_net4225), .RN(npu_inst_pe_1_1_3_n8), .Q(
        npu_inst_int_data_res_1__3__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_3_n32), .CK(
        npu_inst_pe_1_1_3_net4225), .RN(npu_inst_pe_1_1_3_n8), .Q(
        npu_inst_int_data_res_1__3__7_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_3_n100), 
        .CK(npu_inst_pe_1_1_3_net4225), .RN(npu_inst_pe_1_1_3_n8), .Q(
        npu_inst_int_data_res_1__3__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_weight_reg_0_ ( .D(npu_inst_n94), .CK(
        npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n8), .Q(
        npu_inst_pe_1_1_3_int_q_weight_0_), .QN(npu_inst_pe_1_1_3_n27) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_weight_reg_1_ ( .D(npu_inst_n100), .CK(
        npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n8), .Q(
        npu_inst_pe_1_1_3_int_q_weight_1_), .QN(npu_inst_pe_1_1_3_n26) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_3_n112), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n8), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_3_n106), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n8), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_3_n111), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_3_n105), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_3_n110), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_3_n104), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_3_n109), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_3_n103), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_3_n108), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_3_n102), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_3_n107), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_3_n101), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_3_n86), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_3_n87), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n9), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_3_n88), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_3_n89), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_3_n90), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_3_n91), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_3_n92), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_3_n93), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_3_n94), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_3_n95), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_3_n96), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_3_n97), 
        .CK(npu_inst_pe_1_1_3_net4231), .RN(npu_inst_pe_1_1_3_n10), .Q(
        npu_inst_pe_1_1_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_3_net4225) );
  CLKGATETST_X1 npu_inst_pe_1_1_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n47), .SE(1'b0), .GCK(npu_inst_pe_1_1_3_net4231) );
  MUX2_X1 npu_inst_pe_1_1_4_U153 ( .A(npu_inst_pe_1_1_4_n31), .B(
        npu_inst_pe_1_1_4_n28), .S(npu_inst_pe_1_1_4_n7), .Z(
        npu_inst_pe_1_1_4_N93) );
  MUX2_X1 npu_inst_pe_1_1_4_U152 ( .A(npu_inst_pe_1_1_4_n30), .B(
        npu_inst_pe_1_1_4_n29), .S(npu_inst_pe_1_1_4_n5), .Z(
        npu_inst_pe_1_1_4_n31) );
  MUX2_X1 npu_inst_pe_1_1_4_U151 ( .A(npu_inst_pe_1_1_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_4_n3), .Z(
        npu_inst_pe_1_1_4_n30) );
  MUX2_X1 npu_inst_pe_1_1_4_U150 ( .A(npu_inst_pe_1_1_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_4_n3), .Z(
        npu_inst_pe_1_1_4_n29) );
  MUX2_X1 npu_inst_pe_1_1_4_U149 ( .A(npu_inst_pe_1_1_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_4_n3), .Z(
        npu_inst_pe_1_1_4_n28) );
  MUX2_X1 npu_inst_pe_1_1_4_U148 ( .A(npu_inst_pe_1_1_4_n25), .B(
        npu_inst_pe_1_1_4_n22), .S(npu_inst_pe_1_1_4_n7), .Z(
        npu_inst_pe_1_1_4_N94) );
  MUX2_X1 npu_inst_pe_1_1_4_U147 ( .A(npu_inst_pe_1_1_4_n24), .B(
        npu_inst_pe_1_1_4_n23), .S(npu_inst_pe_1_1_4_n5), .Z(
        npu_inst_pe_1_1_4_n25) );
  MUX2_X1 npu_inst_pe_1_1_4_U146 ( .A(npu_inst_pe_1_1_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_4_n3), .Z(
        npu_inst_pe_1_1_4_n24) );
  MUX2_X1 npu_inst_pe_1_1_4_U145 ( .A(npu_inst_pe_1_1_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_4_n3), .Z(
        npu_inst_pe_1_1_4_n23) );
  MUX2_X1 npu_inst_pe_1_1_4_U144 ( .A(npu_inst_pe_1_1_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_4_n3), .Z(
        npu_inst_pe_1_1_4_n22) );
  MUX2_X1 npu_inst_pe_1_1_4_U143 ( .A(npu_inst_pe_1_1_4_n21), .B(
        npu_inst_pe_1_1_4_n18), .S(npu_inst_pe_1_1_4_n7), .Z(
        npu_inst_int_data_x_1__4__1_) );
  MUX2_X1 npu_inst_pe_1_1_4_U142 ( .A(npu_inst_pe_1_1_4_n20), .B(
        npu_inst_pe_1_1_4_n19), .S(npu_inst_pe_1_1_4_n5), .Z(
        npu_inst_pe_1_1_4_n21) );
  MUX2_X1 npu_inst_pe_1_1_4_U141 ( .A(npu_inst_pe_1_1_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_4_n3), .Z(
        npu_inst_pe_1_1_4_n20) );
  MUX2_X1 npu_inst_pe_1_1_4_U140 ( .A(npu_inst_pe_1_1_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_4_n3), .Z(
        npu_inst_pe_1_1_4_n19) );
  MUX2_X1 npu_inst_pe_1_1_4_U139 ( .A(npu_inst_pe_1_1_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_4_n3), .Z(
        npu_inst_pe_1_1_4_n18) );
  MUX2_X1 npu_inst_pe_1_1_4_U138 ( .A(npu_inst_pe_1_1_4_n17), .B(
        npu_inst_pe_1_1_4_n14), .S(npu_inst_pe_1_1_4_n7), .Z(
        npu_inst_int_data_x_1__4__0_) );
  MUX2_X1 npu_inst_pe_1_1_4_U137 ( .A(npu_inst_pe_1_1_4_n16), .B(
        npu_inst_pe_1_1_4_n15), .S(npu_inst_pe_1_1_4_n5), .Z(
        npu_inst_pe_1_1_4_n17) );
  MUX2_X1 npu_inst_pe_1_1_4_U136 ( .A(npu_inst_pe_1_1_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_4_n3), .Z(
        npu_inst_pe_1_1_4_n16) );
  MUX2_X1 npu_inst_pe_1_1_4_U135 ( .A(npu_inst_pe_1_1_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_4_n3), .Z(
        npu_inst_pe_1_1_4_n15) );
  MUX2_X1 npu_inst_pe_1_1_4_U134 ( .A(npu_inst_pe_1_1_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_4_n3), .Z(
        npu_inst_pe_1_1_4_n14) );
  XOR2_X1 npu_inst_pe_1_1_4_U133 ( .A(npu_inst_pe_1_1_4_int_data_0_), .B(
        npu_inst_int_data_res_1__4__0_), .Z(npu_inst_pe_1_1_4_N73) );
  AND2_X1 npu_inst_pe_1_1_4_U132 ( .A1(npu_inst_int_data_res_1__4__0_), .A2(
        npu_inst_pe_1_1_4_int_data_0_), .ZN(npu_inst_pe_1_1_4_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_4_U131 ( .A(npu_inst_int_data_res_1__4__0_), .B(
        npu_inst_pe_1_1_4_n12), .ZN(npu_inst_pe_1_1_4_N65) );
  OR2_X1 npu_inst_pe_1_1_4_U130 ( .A1(npu_inst_pe_1_1_4_n12), .A2(
        npu_inst_int_data_res_1__4__0_), .ZN(npu_inst_pe_1_1_4_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_4_U129 ( .A(npu_inst_int_data_res_1__4__2_), .B(
        npu_inst_pe_1_1_4_add_79_carry_2_), .Z(npu_inst_pe_1_1_4_N75) );
  AND2_X1 npu_inst_pe_1_1_4_U128 ( .A1(npu_inst_pe_1_1_4_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_1__4__2_), .ZN(
        npu_inst_pe_1_1_4_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_4_U127 ( .A(npu_inst_int_data_res_1__4__3_), .B(
        npu_inst_pe_1_1_4_add_79_carry_3_), .Z(npu_inst_pe_1_1_4_N76) );
  AND2_X1 npu_inst_pe_1_1_4_U126 ( .A1(npu_inst_pe_1_1_4_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_1__4__3_), .ZN(
        npu_inst_pe_1_1_4_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_4_U125 ( .A(npu_inst_int_data_res_1__4__4_), .B(
        npu_inst_pe_1_1_4_add_79_carry_4_), .Z(npu_inst_pe_1_1_4_N77) );
  AND2_X1 npu_inst_pe_1_1_4_U124 ( .A1(npu_inst_pe_1_1_4_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_1__4__4_), .ZN(
        npu_inst_pe_1_1_4_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_4_U123 ( .A(npu_inst_int_data_res_1__4__5_), .B(
        npu_inst_pe_1_1_4_add_79_carry_5_), .Z(npu_inst_pe_1_1_4_N78) );
  AND2_X1 npu_inst_pe_1_1_4_U122 ( .A1(npu_inst_pe_1_1_4_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_1__4__5_), .ZN(
        npu_inst_pe_1_1_4_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_4_U121 ( .A(npu_inst_int_data_res_1__4__6_), .B(
        npu_inst_pe_1_1_4_add_79_carry_6_), .Z(npu_inst_pe_1_1_4_N79) );
  AND2_X1 npu_inst_pe_1_1_4_U120 ( .A1(npu_inst_pe_1_1_4_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_1__4__6_), .ZN(
        npu_inst_pe_1_1_4_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_4_U119 ( .A(npu_inst_int_data_res_1__4__7_), .B(
        npu_inst_pe_1_1_4_add_79_carry_7_), .Z(npu_inst_pe_1_1_4_N80) );
  XNOR2_X1 npu_inst_pe_1_1_4_U118 ( .A(npu_inst_pe_1_1_4_sub_77_carry_2_), .B(
        npu_inst_int_data_res_1__4__2_), .ZN(npu_inst_pe_1_1_4_N67) );
  OR2_X1 npu_inst_pe_1_1_4_U117 ( .A1(npu_inst_int_data_res_1__4__2_), .A2(
        npu_inst_pe_1_1_4_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_1_4_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_4_U116 ( .A(npu_inst_pe_1_1_4_sub_77_carry_3_), .B(
        npu_inst_int_data_res_1__4__3_), .ZN(npu_inst_pe_1_1_4_N68) );
  OR2_X1 npu_inst_pe_1_1_4_U115 ( .A1(npu_inst_int_data_res_1__4__3_), .A2(
        npu_inst_pe_1_1_4_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_1_4_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_4_U114 ( .A(npu_inst_pe_1_1_4_sub_77_carry_4_), .B(
        npu_inst_int_data_res_1__4__4_), .ZN(npu_inst_pe_1_1_4_N69) );
  OR2_X1 npu_inst_pe_1_1_4_U113 ( .A1(npu_inst_int_data_res_1__4__4_), .A2(
        npu_inst_pe_1_1_4_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_1_4_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_4_U112 ( .A(npu_inst_pe_1_1_4_sub_77_carry_5_), .B(
        npu_inst_int_data_res_1__4__5_), .ZN(npu_inst_pe_1_1_4_N70) );
  OR2_X1 npu_inst_pe_1_1_4_U111 ( .A1(npu_inst_int_data_res_1__4__5_), .A2(
        npu_inst_pe_1_1_4_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_1_4_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_4_U110 ( .A(npu_inst_pe_1_1_4_sub_77_carry_6_), .B(
        npu_inst_int_data_res_1__4__6_), .ZN(npu_inst_pe_1_1_4_N71) );
  OR2_X1 npu_inst_pe_1_1_4_U109 ( .A1(npu_inst_int_data_res_1__4__6_), .A2(
        npu_inst_pe_1_1_4_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_1_4_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_4_U108 ( .A(npu_inst_int_data_res_1__4__7_), .B(
        npu_inst_pe_1_1_4_sub_77_carry_7_), .ZN(npu_inst_pe_1_1_4_N72) );
  INV_X1 npu_inst_pe_1_1_4_U107 ( .A(npu_inst_n61), .ZN(npu_inst_pe_1_1_4_n6)
         );
  INV_X1 npu_inst_pe_1_1_4_U106 ( .A(npu_inst_pe_1_1_4_n6), .ZN(
        npu_inst_pe_1_1_4_n5) );
  INV_X1 npu_inst_pe_1_1_4_U105 ( .A(npu_inst_n41), .ZN(npu_inst_pe_1_1_4_n2)
         );
  AOI22_X1 npu_inst_pe_1_1_4_U104 ( .A1(npu_inst_int_data_y_2__4__0_), .A2(
        npu_inst_pe_1_1_4_n58), .B1(npu_inst_pe_1_1_4_n118), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_4_n57) );
  INV_X1 npu_inst_pe_1_1_4_U103 ( .A(npu_inst_pe_1_1_4_n57), .ZN(
        npu_inst_pe_1_1_4_n107) );
  AOI22_X1 npu_inst_pe_1_1_4_U102 ( .A1(npu_inst_int_data_y_2__4__0_), .A2(
        npu_inst_pe_1_1_4_n54), .B1(npu_inst_pe_1_1_4_n117), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_4_n53) );
  INV_X1 npu_inst_pe_1_1_4_U99 ( .A(npu_inst_pe_1_1_4_n53), .ZN(
        npu_inst_pe_1_1_4_n108) );
  AOI22_X1 npu_inst_pe_1_1_4_U98 ( .A1(npu_inst_int_data_y_2__4__0_), .A2(
        npu_inst_pe_1_1_4_n50), .B1(npu_inst_pe_1_1_4_n116), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_4_n49) );
  INV_X1 npu_inst_pe_1_1_4_U97 ( .A(npu_inst_pe_1_1_4_n49), .ZN(
        npu_inst_pe_1_1_4_n109) );
  AOI22_X1 npu_inst_pe_1_1_4_U96 ( .A1(npu_inst_int_data_y_2__4__0_), .A2(
        npu_inst_pe_1_1_4_n46), .B1(npu_inst_pe_1_1_4_n115), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_4_n45) );
  INV_X1 npu_inst_pe_1_1_4_U95 ( .A(npu_inst_pe_1_1_4_n45), .ZN(
        npu_inst_pe_1_1_4_n110) );
  AOI22_X1 npu_inst_pe_1_1_4_U94 ( .A1(npu_inst_int_data_y_2__4__0_), .A2(
        npu_inst_pe_1_1_4_n42), .B1(npu_inst_pe_1_1_4_n114), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_4_n41) );
  INV_X1 npu_inst_pe_1_1_4_U93 ( .A(npu_inst_pe_1_1_4_n41), .ZN(
        npu_inst_pe_1_1_4_n111) );
  AOI22_X1 npu_inst_pe_1_1_4_U92 ( .A1(npu_inst_int_data_y_2__4__1_), .A2(
        npu_inst_pe_1_1_4_n58), .B1(npu_inst_pe_1_1_4_n118), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_4_n59) );
  INV_X1 npu_inst_pe_1_1_4_U91 ( .A(npu_inst_pe_1_1_4_n59), .ZN(
        npu_inst_pe_1_1_4_n101) );
  AOI22_X1 npu_inst_pe_1_1_4_U90 ( .A1(npu_inst_int_data_y_2__4__1_), .A2(
        npu_inst_pe_1_1_4_n54), .B1(npu_inst_pe_1_1_4_n117), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_4_n55) );
  INV_X1 npu_inst_pe_1_1_4_U89 ( .A(npu_inst_pe_1_1_4_n55), .ZN(
        npu_inst_pe_1_1_4_n102) );
  AOI22_X1 npu_inst_pe_1_1_4_U88 ( .A1(npu_inst_int_data_y_2__4__1_), .A2(
        npu_inst_pe_1_1_4_n50), .B1(npu_inst_pe_1_1_4_n116), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_4_n51) );
  INV_X1 npu_inst_pe_1_1_4_U87 ( .A(npu_inst_pe_1_1_4_n51), .ZN(
        npu_inst_pe_1_1_4_n103) );
  AOI22_X1 npu_inst_pe_1_1_4_U86 ( .A1(npu_inst_int_data_y_2__4__1_), .A2(
        npu_inst_pe_1_1_4_n46), .B1(npu_inst_pe_1_1_4_n115), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_4_n47) );
  INV_X1 npu_inst_pe_1_1_4_U85 ( .A(npu_inst_pe_1_1_4_n47), .ZN(
        npu_inst_pe_1_1_4_n104) );
  AOI22_X1 npu_inst_pe_1_1_4_U84 ( .A1(npu_inst_int_data_y_2__4__1_), .A2(
        npu_inst_pe_1_1_4_n42), .B1(npu_inst_pe_1_1_4_n114), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_4_n43) );
  INV_X1 npu_inst_pe_1_1_4_U83 ( .A(npu_inst_pe_1_1_4_n43), .ZN(
        npu_inst_pe_1_1_4_n105) );
  AOI22_X1 npu_inst_pe_1_1_4_U82 ( .A1(npu_inst_pe_1_1_4_n38), .A2(
        npu_inst_int_data_y_2__4__1_), .B1(npu_inst_pe_1_1_4_n113), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_4_n39) );
  INV_X1 npu_inst_pe_1_1_4_U81 ( .A(npu_inst_pe_1_1_4_n39), .ZN(
        npu_inst_pe_1_1_4_n106) );
  AND2_X1 npu_inst_pe_1_1_4_U80 ( .A1(npu_inst_pe_1_1_4_N93), .A2(npu_inst_n41), .ZN(npu_inst_int_data_y_1__4__0_) );
  NAND2_X1 npu_inst_pe_1_1_4_U79 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_4_n60), .ZN(npu_inst_pe_1_1_4_n74) );
  OAI21_X1 npu_inst_pe_1_1_4_U78 ( .B1(npu_inst_pe_1_1_4_n63), .B2(
        npu_inst_pe_1_1_4_n60), .A(npu_inst_pe_1_1_4_n74), .ZN(
        npu_inst_pe_1_1_4_n97) );
  NAND2_X1 npu_inst_pe_1_1_4_U77 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_4_n60), .ZN(npu_inst_pe_1_1_4_n73) );
  OAI21_X1 npu_inst_pe_1_1_4_U76 ( .B1(npu_inst_pe_1_1_4_n61), .B2(
        npu_inst_pe_1_1_4_n60), .A(npu_inst_pe_1_1_4_n73), .ZN(
        npu_inst_pe_1_1_4_n96) );
  NAND2_X1 npu_inst_pe_1_1_4_U75 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_4_n56), .ZN(npu_inst_pe_1_1_4_n72) );
  OAI21_X1 npu_inst_pe_1_1_4_U74 ( .B1(npu_inst_pe_1_1_4_n63), .B2(
        npu_inst_pe_1_1_4_n56), .A(npu_inst_pe_1_1_4_n72), .ZN(
        npu_inst_pe_1_1_4_n95) );
  NAND2_X1 npu_inst_pe_1_1_4_U73 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_4_n56), .ZN(npu_inst_pe_1_1_4_n71) );
  OAI21_X1 npu_inst_pe_1_1_4_U72 ( .B1(npu_inst_pe_1_1_4_n61), .B2(
        npu_inst_pe_1_1_4_n56), .A(npu_inst_pe_1_1_4_n71), .ZN(
        npu_inst_pe_1_1_4_n94) );
  NAND2_X1 npu_inst_pe_1_1_4_U71 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_4_n52), .ZN(npu_inst_pe_1_1_4_n70) );
  OAI21_X1 npu_inst_pe_1_1_4_U70 ( .B1(npu_inst_pe_1_1_4_n63), .B2(
        npu_inst_pe_1_1_4_n52), .A(npu_inst_pe_1_1_4_n70), .ZN(
        npu_inst_pe_1_1_4_n93) );
  NAND2_X1 npu_inst_pe_1_1_4_U69 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_4_n52), .ZN(npu_inst_pe_1_1_4_n69) );
  OAI21_X1 npu_inst_pe_1_1_4_U68 ( .B1(npu_inst_pe_1_1_4_n61), .B2(
        npu_inst_pe_1_1_4_n52), .A(npu_inst_pe_1_1_4_n69), .ZN(
        npu_inst_pe_1_1_4_n92) );
  NAND2_X1 npu_inst_pe_1_1_4_U67 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_4_n48), .ZN(npu_inst_pe_1_1_4_n68) );
  OAI21_X1 npu_inst_pe_1_1_4_U66 ( .B1(npu_inst_pe_1_1_4_n63), .B2(
        npu_inst_pe_1_1_4_n48), .A(npu_inst_pe_1_1_4_n68), .ZN(
        npu_inst_pe_1_1_4_n91) );
  NAND2_X1 npu_inst_pe_1_1_4_U65 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_4_n48), .ZN(npu_inst_pe_1_1_4_n67) );
  OAI21_X1 npu_inst_pe_1_1_4_U64 ( .B1(npu_inst_pe_1_1_4_n61), .B2(
        npu_inst_pe_1_1_4_n48), .A(npu_inst_pe_1_1_4_n67), .ZN(
        npu_inst_pe_1_1_4_n90) );
  NAND2_X1 npu_inst_pe_1_1_4_U63 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_4_n44), .ZN(npu_inst_pe_1_1_4_n66) );
  OAI21_X1 npu_inst_pe_1_1_4_U62 ( .B1(npu_inst_pe_1_1_4_n63), .B2(
        npu_inst_pe_1_1_4_n44), .A(npu_inst_pe_1_1_4_n66), .ZN(
        npu_inst_pe_1_1_4_n89) );
  NAND2_X1 npu_inst_pe_1_1_4_U61 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_4_n44), .ZN(npu_inst_pe_1_1_4_n65) );
  OAI21_X1 npu_inst_pe_1_1_4_U60 ( .B1(npu_inst_pe_1_1_4_n61), .B2(
        npu_inst_pe_1_1_4_n44), .A(npu_inst_pe_1_1_4_n65), .ZN(
        npu_inst_pe_1_1_4_n88) );
  NAND2_X1 npu_inst_pe_1_1_4_U59 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_4_n40), .ZN(npu_inst_pe_1_1_4_n64) );
  OAI21_X1 npu_inst_pe_1_1_4_U58 ( .B1(npu_inst_pe_1_1_4_n63), .B2(
        npu_inst_pe_1_1_4_n40), .A(npu_inst_pe_1_1_4_n64), .ZN(
        npu_inst_pe_1_1_4_n87) );
  NAND2_X1 npu_inst_pe_1_1_4_U57 ( .A1(npu_inst_pe_1_1_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_4_n40), .ZN(npu_inst_pe_1_1_4_n62) );
  OAI21_X1 npu_inst_pe_1_1_4_U56 ( .B1(npu_inst_pe_1_1_4_n61), .B2(
        npu_inst_pe_1_1_4_n40), .A(npu_inst_pe_1_1_4_n62), .ZN(
        npu_inst_pe_1_1_4_n86) );
  AOI22_X1 npu_inst_pe_1_1_4_U55 ( .A1(npu_inst_pe_1_1_4_n38), .A2(
        npu_inst_int_data_y_2__4__0_), .B1(npu_inst_pe_1_1_4_n113), .B2(
        npu_inst_pe_1_1_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_4_n37) );
  INV_X1 npu_inst_pe_1_1_4_U54 ( .A(npu_inst_pe_1_1_4_n37), .ZN(
        npu_inst_pe_1_1_4_n112) );
  AND2_X1 npu_inst_pe_1_1_4_U53 ( .A1(npu_inst_n41), .A2(npu_inst_pe_1_1_4_N94), .ZN(npu_inst_int_data_y_1__4__1_) );
  AOI222_X1 npu_inst_pe_1_1_4_U52 ( .A1(npu_inst_int_data_res_2__4__0_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N73), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N65), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n84) );
  INV_X1 npu_inst_pe_1_1_4_U51 ( .A(npu_inst_pe_1_1_4_n84), .ZN(
        npu_inst_pe_1_1_4_n100) );
  AOI222_X1 npu_inst_pe_1_1_4_U50 ( .A1(npu_inst_pe_1_1_4_n1), .A2(
        npu_inst_int_data_res_2__4__7_), .B1(npu_inst_pe_1_1_4_N80), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N72), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n75) );
  INV_X1 npu_inst_pe_1_1_4_U49 ( .A(npu_inst_pe_1_1_4_n75), .ZN(
        npu_inst_pe_1_1_4_n32) );
  AOI222_X1 npu_inst_pe_1_1_4_U48 ( .A1(npu_inst_int_data_res_2__4__1_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N74), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N66), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n83) );
  INV_X1 npu_inst_pe_1_1_4_U47 ( .A(npu_inst_pe_1_1_4_n83), .ZN(
        npu_inst_pe_1_1_4_n99) );
  AOI222_X1 npu_inst_pe_1_1_4_U46 ( .A1(npu_inst_int_data_res_2__4__3_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N76), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N68), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n81) );
  INV_X1 npu_inst_pe_1_1_4_U45 ( .A(npu_inst_pe_1_1_4_n81), .ZN(
        npu_inst_pe_1_1_4_n36) );
  AOI222_X1 npu_inst_pe_1_1_4_U44 ( .A1(npu_inst_int_data_res_2__4__4_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N77), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N69), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n80) );
  INV_X1 npu_inst_pe_1_1_4_U43 ( .A(npu_inst_pe_1_1_4_n80), .ZN(
        npu_inst_pe_1_1_4_n35) );
  AOI222_X1 npu_inst_pe_1_1_4_U42 ( .A1(npu_inst_int_data_res_2__4__5_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N78), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N70), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n79) );
  INV_X1 npu_inst_pe_1_1_4_U41 ( .A(npu_inst_pe_1_1_4_n79), .ZN(
        npu_inst_pe_1_1_4_n34) );
  AOI222_X1 npu_inst_pe_1_1_4_U40 ( .A1(npu_inst_int_data_res_2__4__6_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N79), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N71), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n78) );
  INV_X1 npu_inst_pe_1_1_4_U39 ( .A(npu_inst_pe_1_1_4_n78), .ZN(
        npu_inst_pe_1_1_4_n33) );
  AND2_X1 npu_inst_pe_1_1_4_U38 ( .A1(npu_inst_int_data_x_1__4__1_), .A2(
        npu_inst_pe_1_1_4_int_q_weight_1_), .ZN(npu_inst_pe_1_1_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_4_U37 ( .A1(npu_inst_int_data_x_1__4__0_), .A2(
        npu_inst_pe_1_1_4_int_q_weight_1_), .ZN(npu_inst_pe_1_1_4_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_1_4_U36 ( .A(npu_inst_pe_1_1_4_int_data_1_), .ZN(
        npu_inst_pe_1_1_4_n13) );
  NOR3_X1 npu_inst_pe_1_1_4_U35 ( .A1(npu_inst_pe_1_1_4_n26), .A2(npu_inst_n41), .A3(npu_inst_int_ckg[51]), .ZN(npu_inst_pe_1_1_4_n85) );
  OR2_X1 npu_inst_pe_1_1_4_U34 ( .A1(npu_inst_pe_1_1_4_n85), .A2(
        npu_inst_pe_1_1_4_n1), .ZN(npu_inst_pe_1_1_4_N84) );
  AOI222_X1 npu_inst_pe_1_1_4_U33 ( .A1(npu_inst_int_data_res_2__4__2_), .A2(
        npu_inst_pe_1_1_4_n1), .B1(npu_inst_pe_1_1_4_N75), .B2(
        npu_inst_pe_1_1_4_n76), .C1(npu_inst_pe_1_1_4_N67), .C2(
        npu_inst_pe_1_1_4_n77), .ZN(npu_inst_pe_1_1_4_n82) );
  INV_X1 npu_inst_pe_1_1_4_U32 ( .A(npu_inst_pe_1_1_4_n82), .ZN(
        npu_inst_pe_1_1_4_n98) );
  AOI22_X1 npu_inst_pe_1_1_4_U31 ( .A1(npu_inst_n41), .A2(
        npu_inst_int_data_y_2__4__1_), .B1(npu_inst_pe_1_1_4_n2), .B2(
        npu_inst_int_data_x_1__5__1_), .ZN(npu_inst_pe_1_1_4_n63) );
  AOI22_X1 npu_inst_pe_1_1_4_U30 ( .A1(npu_inst_n41), .A2(
        npu_inst_int_data_y_2__4__0_), .B1(npu_inst_pe_1_1_4_n2), .B2(
        npu_inst_int_data_x_1__5__0_), .ZN(npu_inst_pe_1_1_4_n61) );
  INV_X1 npu_inst_pe_1_1_4_U29 ( .A(npu_inst_pe_1_1_4_int_data_0_), .ZN(
        npu_inst_pe_1_1_4_n12) );
  INV_X1 npu_inst_pe_1_1_4_U28 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_1_4_n4)
         );
  OR3_X1 npu_inst_pe_1_1_4_U27 ( .A1(npu_inst_pe_1_1_4_n5), .A2(
        npu_inst_pe_1_1_4_n7), .A3(npu_inst_pe_1_1_4_n4), .ZN(
        npu_inst_pe_1_1_4_n56) );
  OR3_X1 npu_inst_pe_1_1_4_U26 ( .A1(npu_inst_pe_1_1_4_n4), .A2(
        npu_inst_pe_1_1_4_n7), .A3(npu_inst_pe_1_1_4_n6), .ZN(
        npu_inst_pe_1_1_4_n48) );
  INV_X1 npu_inst_pe_1_1_4_U25 ( .A(npu_inst_pe_1_1_4_n4), .ZN(
        npu_inst_pe_1_1_4_n3) );
  OR3_X1 npu_inst_pe_1_1_4_U24 ( .A1(npu_inst_pe_1_1_4_n3), .A2(
        npu_inst_pe_1_1_4_n7), .A3(npu_inst_pe_1_1_4_n6), .ZN(
        npu_inst_pe_1_1_4_n52) );
  OR3_X1 npu_inst_pe_1_1_4_U23 ( .A1(npu_inst_pe_1_1_4_n5), .A2(
        npu_inst_pe_1_1_4_n7), .A3(npu_inst_pe_1_1_4_n3), .ZN(
        npu_inst_pe_1_1_4_n60) );
  BUF_X1 npu_inst_pe_1_1_4_U22 ( .A(npu_inst_n28), .Z(npu_inst_pe_1_1_4_n1) );
  NOR2_X1 npu_inst_pe_1_1_4_U21 ( .A1(npu_inst_pe_1_1_4_n60), .A2(
        npu_inst_pe_1_1_4_n2), .ZN(npu_inst_pe_1_1_4_n58) );
  NOR2_X1 npu_inst_pe_1_1_4_U20 ( .A1(npu_inst_pe_1_1_4_n56), .A2(
        npu_inst_pe_1_1_4_n2), .ZN(npu_inst_pe_1_1_4_n54) );
  NOR2_X1 npu_inst_pe_1_1_4_U19 ( .A1(npu_inst_pe_1_1_4_n52), .A2(
        npu_inst_pe_1_1_4_n2), .ZN(npu_inst_pe_1_1_4_n50) );
  NOR2_X1 npu_inst_pe_1_1_4_U18 ( .A1(npu_inst_pe_1_1_4_n48), .A2(
        npu_inst_pe_1_1_4_n2), .ZN(npu_inst_pe_1_1_4_n46) );
  NOR2_X1 npu_inst_pe_1_1_4_U17 ( .A1(npu_inst_pe_1_1_4_n40), .A2(
        npu_inst_pe_1_1_4_n2), .ZN(npu_inst_pe_1_1_4_n38) );
  NOR2_X1 npu_inst_pe_1_1_4_U16 ( .A1(npu_inst_pe_1_1_4_n44), .A2(
        npu_inst_pe_1_1_4_n2), .ZN(npu_inst_pe_1_1_4_n42) );
  BUF_X1 npu_inst_pe_1_1_4_U15 ( .A(npu_inst_n86), .Z(npu_inst_pe_1_1_4_n7) );
  INV_X1 npu_inst_pe_1_1_4_U14 ( .A(npu_inst_n108), .ZN(npu_inst_pe_1_1_4_n11)
         );
  INV_X1 npu_inst_pe_1_1_4_U13 ( .A(npu_inst_pe_1_1_4_n38), .ZN(
        npu_inst_pe_1_1_4_n113) );
  INV_X1 npu_inst_pe_1_1_4_U12 ( .A(npu_inst_pe_1_1_4_n58), .ZN(
        npu_inst_pe_1_1_4_n118) );
  INV_X1 npu_inst_pe_1_1_4_U11 ( .A(npu_inst_pe_1_1_4_n54), .ZN(
        npu_inst_pe_1_1_4_n117) );
  INV_X1 npu_inst_pe_1_1_4_U10 ( .A(npu_inst_pe_1_1_4_n50), .ZN(
        npu_inst_pe_1_1_4_n116) );
  INV_X1 npu_inst_pe_1_1_4_U9 ( .A(npu_inst_pe_1_1_4_n46), .ZN(
        npu_inst_pe_1_1_4_n115) );
  INV_X1 npu_inst_pe_1_1_4_U8 ( .A(npu_inst_pe_1_1_4_n42), .ZN(
        npu_inst_pe_1_1_4_n114) );
  BUF_X1 npu_inst_pe_1_1_4_U7 ( .A(npu_inst_pe_1_1_4_n11), .Z(
        npu_inst_pe_1_1_4_n10) );
  BUF_X1 npu_inst_pe_1_1_4_U6 ( .A(npu_inst_pe_1_1_4_n11), .Z(
        npu_inst_pe_1_1_4_n9) );
  BUF_X1 npu_inst_pe_1_1_4_U5 ( .A(npu_inst_pe_1_1_4_n11), .Z(
        npu_inst_pe_1_1_4_n8) );
  NOR2_X1 npu_inst_pe_1_1_4_U4 ( .A1(npu_inst_pe_1_1_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_4_n1), .ZN(npu_inst_pe_1_1_4_n76) );
  NOR2_X1 npu_inst_pe_1_1_4_U3 ( .A1(npu_inst_pe_1_1_4_n27), .A2(
        npu_inst_pe_1_1_4_n1), .ZN(npu_inst_pe_1_1_4_n77) );
  FA_X1 npu_inst_pe_1_1_4_sub_77_U2_1 ( .A(npu_inst_int_data_res_1__4__1_), 
        .B(npu_inst_pe_1_1_4_n13), .CI(npu_inst_pe_1_1_4_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_1_4_sub_77_carry_2_), .S(npu_inst_pe_1_1_4_N66) );
  FA_X1 npu_inst_pe_1_1_4_add_79_U1_1 ( .A(npu_inst_int_data_res_1__4__1_), 
        .B(npu_inst_pe_1_1_4_int_data_1_), .CI(
        npu_inst_pe_1_1_4_add_79_carry_1_), .CO(
        npu_inst_pe_1_1_4_add_79_carry_2_), .S(npu_inst_pe_1_1_4_N74) );
  NAND3_X1 npu_inst_pe_1_1_4_U101 ( .A1(npu_inst_pe_1_1_4_n4), .A2(
        npu_inst_pe_1_1_4_n6), .A3(npu_inst_pe_1_1_4_n7), .ZN(
        npu_inst_pe_1_1_4_n44) );
  NAND3_X1 npu_inst_pe_1_1_4_U100 ( .A1(npu_inst_pe_1_1_4_n3), .A2(
        npu_inst_pe_1_1_4_n6), .A3(npu_inst_pe_1_1_4_n7), .ZN(
        npu_inst_pe_1_1_4_n40) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_4_n33), .CK(
        npu_inst_pe_1_1_4_net4202), .RN(npu_inst_pe_1_1_4_n8), .Q(
        npu_inst_int_data_res_1__4__6_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_4_n34), .CK(
        npu_inst_pe_1_1_4_net4202), .RN(npu_inst_pe_1_1_4_n8), .Q(
        npu_inst_int_data_res_1__4__5_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_4_n35), .CK(
        npu_inst_pe_1_1_4_net4202), .RN(npu_inst_pe_1_1_4_n8), .Q(
        npu_inst_int_data_res_1__4__4_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_4_n36), .CK(
        npu_inst_pe_1_1_4_net4202), .RN(npu_inst_pe_1_1_4_n8), .Q(
        npu_inst_int_data_res_1__4__3_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_4_n98), .CK(
        npu_inst_pe_1_1_4_net4202), .RN(npu_inst_pe_1_1_4_n8), .Q(
        npu_inst_int_data_res_1__4__2_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_4_n99), .CK(
        npu_inst_pe_1_1_4_net4202), .RN(npu_inst_pe_1_1_4_n8), .Q(
        npu_inst_int_data_res_1__4__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_4_n32), .CK(
        npu_inst_pe_1_1_4_net4202), .RN(npu_inst_pe_1_1_4_n8), .Q(
        npu_inst_int_data_res_1__4__7_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_4_n100), 
        .CK(npu_inst_pe_1_1_4_net4202), .RN(npu_inst_pe_1_1_4_n8), .Q(
        npu_inst_int_data_res_1__4__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_weight_reg_0_ ( .D(npu_inst_n94), .CK(
        npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n8), .Q(
        npu_inst_pe_1_1_4_int_q_weight_0_), .QN(npu_inst_pe_1_1_4_n27) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_weight_reg_1_ ( .D(npu_inst_n100), .CK(
        npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n8), .Q(
        npu_inst_pe_1_1_4_int_q_weight_1_), .QN(npu_inst_pe_1_1_4_n26) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_4_n112), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n8), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_4_n106), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n8), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_4_n111), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_4_n105), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_4_n110), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_4_n104), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_4_n109), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_4_n103), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_4_n108), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_4_n102), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_4_n107), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_4_n101), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_4_n86), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_4_n87), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n9), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_4_n88), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_4_n89), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_4_n90), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_4_n91), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_4_n92), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_4_n93), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_4_n94), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_4_n95), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_4_n96), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_4_n97), 
        .CK(npu_inst_pe_1_1_4_net4208), .RN(npu_inst_pe_1_1_4_n10), .Q(
        npu_inst_pe_1_1_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_4_net4202) );
  CLKGATETST_X1 npu_inst_pe_1_1_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n47), .SE(1'b0), .GCK(npu_inst_pe_1_1_4_net4208) );
  MUX2_X1 npu_inst_pe_1_1_5_U153 ( .A(npu_inst_pe_1_1_5_n31), .B(
        npu_inst_pe_1_1_5_n28), .S(npu_inst_pe_1_1_5_n7), .Z(
        npu_inst_pe_1_1_5_N93) );
  MUX2_X1 npu_inst_pe_1_1_5_U152 ( .A(npu_inst_pe_1_1_5_n30), .B(
        npu_inst_pe_1_1_5_n29), .S(npu_inst_pe_1_1_5_n5), .Z(
        npu_inst_pe_1_1_5_n31) );
  MUX2_X1 npu_inst_pe_1_1_5_U151 ( .A(npu_inst_pe_1_1_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_5_n3), .Z(
        npu_inst_pe_1_1_5_n30) );
  MUX2_X1 npu_inst_pe_1_1_5_U150 ( .A(npu_inst_pe_1_1_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_5_n3), .Z(
        npu_inst_pe_1_1_5_n29) );
  MUX2_X1 npu_inst_pe_1_1_5_U149 ( .A(npu_inst_pe_1_1_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_5_n3), .Z(
        npu_inst_pe_1_1_5_n28) );
  MUX2_X1 npu_inst_pe_1_1_5_U148 ( .A(npu_inst_pe_1_1_5_n25), .B(
        npu_inst_pe_1_1_5_n22), .S(npu_inst_pe_1_1_5_n7), .Z(
        npu_inst_pe_1_1_5_N94) );
  MUX2_X1 npu_inst_pe_1_1_5_U147 ( .A(npu_inst_pe_1_1_5_n24), .B(
        npu_inst_pe_1_1_5_n23), .S(npu_inst_pe_1_1_5_n5), .Z(
        npu_inst_pe_1_1_5_n25) );
  MUX2_X1 npu_inst_pe_1_1_5_U146 ( .A(npu_inst_pe_1_1_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_5_n3), .Z(
        npu_inst_pe_1_1_5_n24) );
  MUX2_X1 npu_inst_pe_1_1_5_U145 ( .A(npu_inst_pe_1_1_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_5_n3), .Z(
        npu_inst_pe_1_1_5_n23) );
  MUX2_X1 npu_inst_pe_1_1_5_U144 ( .A(npu_inst_pe_1_1_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_5_n3), .Z(
        npu_inst_pe_1_1_5_n22) );
  MUX2_X1 npu_inst_pe_1_1_5_U143 ( .A(npu_inst_pe_1_1_5_n21), .B(
        npu_inst_pe_1_1_5_n18), .S(npu_inst_pe_1_1_5_n7), .Z(
        npu_inst_int_data_x_1__5__1_) );
  MUX2_X1 npu_inst_pe_1_1_5_U142 ( .A(npu_inst_pe_1_1_5_n20), .B(
        npu_inst_pe_1_1_5_n19), .S(npu_inst_pe_1_1_5_n5), .Z(
        npu_inst_pe_1_1_5_n21) );
  MUX2_X1 npu_inst_pe_1_1_5_U141 ( .A(npu_inst_pe_1_1_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_5_n3), .Z(
        npu_inst_pe_1_1_5_n20) );
  MUX2_X1 npu_inst_pe_1_1_5_U140 ( .A(npu_inst_pe_1_1_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_5_n3), .Z(
        npu_inst_pe_1_1_5_n19) );
  MUX2_X1 npu_inst_pe_1_1_5_U139 ( .A(npu_inst_pe_1_1_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_5_n3), .Z(
        npu_inst_pe_1_1_5_n18) );
  MUX2_X1 npu_inst_pe_1_1_5_U138 ( .A(npu_inst_pe_1_1_5_n17), .B(
        npu_inst_pe_1_1_5_n14), .S(npu_inst_pe_1_1_5_n7), .Z(
        npu_inst_int_data_x_1__5__0_) );
  MUX2_X1 npu_inst_pe_1_1_5_U137 ( .A(npu_inst_pe_1_1_5_n16), .B(
        npu_inst_pe_1_1_5_n15), .S(npu_inst_pe_1_1_5_n5), .Z(
        npu_inst_pe_1_1_5_n17) );
  MUX2_X1 npu_inst_pe_1_1_5_U136 ( .A(npu_inst_pe_1_1_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_5_n3), .Z(
        npu_inst_pe_1_1_5_n16) );
  MUX2_X1 npu_inst_pe_1_1_5_U135 ( .A(npu_inst_pe_1_1_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_5_n3), .Z(
        npu_inst_pe_1_1_5_n15) );
  MUX2_X1 npu_inst_pe_1_1_5_U134 ( .A(npu_inst_pe_1_1_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_5_n3), .Z(
        npu_inst_pe_1_1_5_n14) );
  XOR2_X1 npu_inst_pe_1_1_5_U133 ( .A(npu_inst_pe_1_1_5_int_data_0_), .B(
        npu_inst_int_data_res_1__5__0_), .Z(npu_inst_pe_1_1_5_N73) );
  AND2_X1 npu_inst_pe_1_1_5_U132 ( .A1(npu_inst_int_data_res_1__5__0_), .A2(
        npu_inst_pe_1_1_5_int_data_0_), .ZN(npu_inst_pe_1_1_5_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_5_U131 ( .A(npu_inst_int_data_res_1__5__0_), .B(
        npu_inst_pe_1_1_5_n12), .ZN(npu_inst_pe_1_1_5_N65) );
  OR2_X1 npu_inst_pe_1_1_5_U130 ( .A1(npu_inst_pe_1_1_5_n12), .A2(
        npu_inst_int_data_res_1__5__0_), .ZN(npu_inst_pe_1_1_5_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_5_U129 ( .A(npu_inst_int_data_res_1__5__2_), .B(
        npu_inst_pe_1_1_5_add_79_carry_2_), .Z(npu_inst_pe_1_1_5_N75) );
  AND2_X1 npu_inst_pe_1_1_5_U128 ( .A1(npu_inst_pe_1_1_5_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_1__5__2_), .ZN(
        npu_inst_pe_1_1_5_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_5_U127 ( .A(npu_inst_int_data_res_1__5__3_), .B(
        npu_inst_pe_1_1_5_add_79_carry_3_), .Z(npu_inst_pe_1_1_5_N76) );
  AND2_X1 npu_inst_pe_1_1_5_U126 ( .A1(npu_inst_pe_1_1_5_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_1__5__3_), .ZN(
        npu_inst_pe_1_1_5_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_5_U125 ( .A(npu_inst_int_data_res_1__5__4_), .B(
        npu_inst_pe_1_1_5_add_79_carry_4_), .Z(npu_inst_pe_1_1_5_N77) );
  AND2_X1 npu_inst_pe_1_1_5_U124 ( .A1(npu_inst_pe_1_1_5_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_1__5__4_), .ZN(
        npu_inst_pe_1_1_5_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_5_U123 ( .A(npu_inst_int_data_res_1__5__5_), .B(
        npu_inst_pe_1_1_5_add_79_carry_5_), .Z(npu_inst_pe_1_1_5_N78) );
  AND2_X1 npu_inst_pe_1_1_5_U122 ( .A1(npu_inst_pe_1_1_5_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_1__5__5_), .ZN(
        npu_inst_pe_1_1_5_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_5_U121 ( .A(npu_inst_int_data_res_1__5__6_), .B(
        npu_inst_pe_1_1_5_add_79_carry_6_), .Z(npu_inst_pe_1_1_5_N79) );
  AND2_X1 npu_inst_pe_1_1_5_U120 ( .A1(npu_inst_pe_1_1_5_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_1__5__6_), .ZN(
        npu_inst_pe_1_1_5_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_5_U119 ( .A(npu_inst_int_data_res_1__5__7_), .B(
        npu_inst_pe_1_1_5_add_79_carry_7_), .Z(npu_inst_pe_1_1_5_N80) );
  XNOR2_X1 npu_inst_pe_1_1_5_U118 ( .A(npu_inst_pe_1_1_5_sub_77_carry_2_), .B(
        npu_inst_int_data_res_1__5__2_), .ZN(npu_inst_pe_1_1_5_N67) );
  OR2_X1 npu_inst_pe_1_1_5_U117 ( .A1(npu_inst_int_data_res_1__5__2_), .A2(
        npu_inst_pe_1_1_5_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_1_5_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_5_U116 ( .A(npu_inst_pe_1_1_5_sub_77_carry_3_), .B(
        npu_inst_int_data_res_1__5__3_), .ZN(npu_inst_pe_1_1_5_N68) );
  OR2_X1 npu_inst_pe_1_1_5_U115 ( .A1(npu_inst_int_data_res_1__5__3_), .A2(
        npu_inst_pe_1_1_5_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_1_5_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_5_U114 ( .A(npu_inst_pe_1_1_5_sub_77_carry_4_), .B(
        npu_inst_int_data_res_1__5__4_), .ZN(npu_inst_pe_1_1_5_N69) );
  OR2_X1 npu_inst_pe_1_1_5_U113 ( .A1(npu_inst_int_data_res_1__5__4_), .A2(
        npu_inst_pe_1_1_5_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_1_5_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_5_U112 ( .A(npu_inst_pe_1_1_5_sub_77_carry_5_), .B(
        npu_inst_int_data_res_1__5__5_), .ZN(npu_inst_pe_1_1_5_N70) );
  OR2_X1 npu_inst_pe_1_1_5_U111 ( .A1(npu_inst_int_data_res_1__5__5_), .A2(
        npu_inst_pe_1_1_5_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_1_5_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_5_U110 ( .A(npu_inst_pe_1_1_5_sub_77_carry_6_), .B(
        npu_inst_int_data_res_1__5__6_), .ZN(npu_inst_pe_1_1_5_N71) );
  OR2_X1 npu_inst_pe_1_1_5_U109 ( .A1(npu_inst_int_data_res_1__5__6_), .A2(
        npu_inst_pe_1_1_5_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_1_5_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_5_U108 ( .A(npu_inst_int_data_res_1__5__7_), .B(
        npu_inst_pe_1_1_5_sub_77_carry_7_), .ZN(npu_inst_pe_1_1_5_N72) );
  INV_X1 npu_inst_pe_1_1_5_U107 ( .A(npu_inst_n61), .ZN(npu_inst_pe_1_1_5_n6)
         );
  INV_X1 npu_inst_pe_1_1_5_U106 ( .A(npu_inst_pe_1_1_5_n6), .ZN(
        npu_inst_pe_1_1_5_n5) );
  INV_X1 npu_inst_pe_1_1_5_U105 ( .A(npu_inst_n41), .ZN(npu_inst_pe_1_1_5_n2)
         );
  AOI22_X1 npu_inst_pe_1_1_5_U104 ( .A1(npu_inst_int_data_y_2__5__0_), .A2(
        npu_inst_pe_1_1_5_n58), .B1(npu_inst_pe_1_1_5_n118), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_5_n57) );
  INV_X1 npu_inst_pe_1_1_5_U103 ( .A(npu_inst_pe_1_1_5_n57), .ZN(
        npu_inst_pe_1_1_5_n107) );
  AOI22_X1 npu_inst_pe_1_1_5_U102 ( .A1(npu_inst_int_data_y_2__5__0_), .A2(
        npu_inst_pe_1_1_5_n54), .B1(npu_inst_pe_1_1_5_n117), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_5_n53) );
  INV_X1 npu_inst_pe_1_1_5_U99 ( .A(npu_inst_pe_1_1_5_n53), .ZN(
        npu_inst_pe_1_1_5_n108) );
  AOI22_X1 npu_inst_pe_1_1_5_U98 ( .A1(npu_inst_int_data_y_2__5__0_), .A2(
        npu_inst_pe_1_1_5_n50), .B1(npu_inst_pe_1_1_5_n116), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_5_n49) );
  INV_X1 npu_inst_pe_1_1_5_U97 ( .A(npu_inst_pe_1_1_5_n49), .ZN(
        npu_inst_pe_1_1_5_n109) );
  AOI22_X1 npu_inst_pe_1_1_5_U96 ( .A1(npu_inst_int_data_y_2__5__0_), .A2(
        npu_inst_pe_1_1_5_n46), .B1(npu_inst_pe_1_1_5_n115), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_5_n45) );
  INV_X1 npu_inst_pe_1_1_5_U95 ( .A(npu_inst_pe_1_1_5_n45), .ZN(
        npu_inst_pe_1_1_5_n110) );
  AOI22_X1 npu_inst_pe_1_1_5_U94 ( .A1(npu_inst_int_data_y_2__5__0_), .A2(
        npu_inst_pe_1_1_5_n42), .B1(npu_inst_pe_1_1_5_n114), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_5_n41) );
  INV_X1 npu_inst_pe_1_1_5_U93 ( .A(npu_inst_pe_1_1_5_n41), .ZN(
        npu_inst_pe_1_1_5_n111) );
  AOI22_X1 npu_inst_pe_1_1_5_U92 ( .A1(npu_inst_int_data_y_2__5__1_), .A2(
        npu_inst_pe_1_1_5_n58), .B1(npu_inst_pe_1_1_5_n118), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_5_n59) );
  INV_X1 npu_inst_pe_1_1_5_U91 ( .A(npu_inst_pe_1_1_5_n59), .ZN(
        npu_inst_pe_1_1_5_n101) );
  AOI22_X1 npu_inst_pe_1_1_5_U90 ( .A1(npu_inst_int_data_y_2__5__1_), .A2(
        npu_inst_pe_1_1_5_n54), .B1(npu_inst_pe_1_1_5_n117), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_5_n55) );
  INV_X1 npu_inst_pe_1_1_5_U89 ( .A(npu_inst_pe_1_1_5_n55), .ZN(
        npu_inst_pe_1_1_5_n102) );
  AOI22_X1 npu_inst_pe_1_1_5_U88 ( .A1(npu_inst_int_data_y_2__5__1_), .A2(
        npu_inst_pe_1_1_5_n50), .B1(npu_inst_pe_1_1_5_n116), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_5_n51) );
  INV_X1 npu_inst_pe_1_1_5_U87 ( .A(npu_inst_pe_1_1_5_n51), .ZN(
        npu_inst_pe_1_1_5_n103) );
  AOI22_X1 npu_inst_pe_1_1_5_U86 ( .A1(npu_inst_int_data_y_2__5__1_), .A2(
        npu_inst_pe_1_1_5_n46), .B1(npu_inst_pe_1_1_5_n115), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_5_n47) );
  INV_X1 npu_inst_pe_1_1_5_U85 ( .A(npu_inst_pe_1_1_5_n47), .ZN(
        npu_inst_pe_1_1_5_n104) );
  AOI22_X1 npu_inst_pe_1_1_5_U84 ( .A1(npu_inst_int_data_y_2__5__1_), .A2(
        npu_inst_pe_1_1_5_n42), .B1(npu_inst_pe_1_1_5_n114), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_5_n43) );
  INV_X1 npu_inst_pe_1_1_5_U83 ( .A(npu_inst_pe_1_1_5_n43), .ZN(
        npu_inst_pe_1_1_5_n105) );
  AOI22_X1 npu_inst_pe_1_1_5_U82 ( .A1(npu_inst_pe_1_1_5_n38), .A2(
        npu_inst_int_data_y_2__5__1_), .B1(npu_inst_pe_1_1_5_n113), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_5_n39) );
  INV_X1 npu_inst_pe_1_1_5_U81 ( .A(npu_inst_pe_1_1_5_n39), .ZN(
        npu_inst_pe_1_1_5_n106) );
  AND2_X1 npu_inst_pe_1_1_5_U80 ( .A1(npu_inst_pe_1_1_5_N93), .A2(npu_inst_n41), .ZN(npu_inst_int_data_y_1__5__0_) );
  NAND2_X1 npu_inst_pe_1_1_5_U79 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_5_n60), .ZN(npu_inst_pe_1_1_5_n74) );
  OAI21_X1 npu_inst_pe_1_1_5_U78 ( .B1(npu_inst_pe_1_1_5_n63), .B2(
        npu_inst_pe_1_1_5_n60), .A(npu_inst_pe_1_1_5_n74), .ZN(
        npu_inst_pe_1_1_5_n97) );
  NAND2_X1 npu_inst_pe_1_1_5_U77 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_5_n60), .ZN(npu_inst_pe_1_1_5_n73) );
  OAI21_X1 npu_inst_pe_1_1_5_U76 ( .B1(npu_inst_pe_1_1_5_n61), .B2(
        npu_inst_pe_1_1_5_n60), .A(npu_inst_pe_1_1_5_n73), .ZN(
        npu_inst_pe_1_1_5_n96) );
  NAND2_X1 npu_inst_pe_1_1_5_U75 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_5_n56), .ZN(npu_inst_pe_1_1_5_n72) );
  OAI21_X1 npu_inst_pe_1_1_5_U74 ( .B1(npu_inst_pe_1_1_5_n63), .B2(
        npu_inst_pe_1_1_5_n56), .A(npu_inst_pe_1_1_5_n72), .ZN(
        npu_inst_pe_1_1_5_n95) );
  NAND2_X1 npu_inst_pe_1_1_5_U73 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_5_n56), .ZN(npu_inst_pe_1_1_5_n71) );
  OAI21_X1 npu_inst_pe_1_1_5_U72 ( .B1(npu_inst_pe_1_1_5_n61), .B2(
        npu_inst_pe_1_1_5_n56), .A(npu_inst_pe_1_1_5_n71), .ZN(
        npu_inst_pe_1_1_5_n94) );
  NAND2_X1 npu_inst_pe_1_1_5_U71 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_5_n52), .ZN(npu_inst_pe_1_1_5_n70) );
  OAI21_X1 npu_inst_pe_1_1_5_U70 ( .B1(npu_inst_pe_1_1_5_n63), .B2(
        npu_inst_pe_1_1_5_n52), .A(npu_inst_pe_1_1_5_n70), .ZN(
        npu_inst_pe_1_1_5_n93) );
  NAND2_X1 npu_inst_pe_1_1_5_U69 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_5_n52), .ZN(npu_inst_pe_1_1_5_n69) );
  OAI21_X1 npu_inst_pe_1_1_5_U68 ( .B1(npu_inst_pe_1_1_5_n61), .B2(
        npu_inst_pe_1_1_5_n52), .A(npu_inst_pe_1_1_5_n69), .ZN(
        npu_inst_pe_1_1_5_n92) );
  NAND2_X1 npu_inst_pe_1_1_5_U67 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_5_n48), .ZN(npu_inst_pe_1_1_5_n68) );
  OAI21_X1 npu_inst_pe_1_1_5_U66 ( .B1(npu_inst_pe_1_1_5_n63), .B2(
        npu_inst_pe_1_1_5_n48), .A(npu_inst_pe_1_1_5_n68), .ZN(
        npu_inst_pe_1_1_5_n91) );
  NAND2_X1 npu_inst_pe_1_1_5_U65 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_5_n48), .ZN(npu_inst_pe_1_1_5_n67) );
  OAI21_X1 npu_inst_pe_1_1_5_U64 ( .B1(npu_inst_pe_1_1_5_n61), .B2(
        npu_inst_pe_1_1_5_n48), .A(npu_inst_pe_1_1_5_n67), .ZN(
        npu_inst_pe_1_1_5_n90) );
  NAND2_X1 npu_inst_pe_1_1_5_U63 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_5_n44), .ZN(npu_inst_pe_1_1_5_n66) );
  OAI21_X1 npu_inst_pe_1_1_5_U62 ( .B1(npu_inst_pe_1_1_5_n63), .B2(
        npu_inst_pe_1_1_5_n44), .A(npu_inst_pe_1_1_5_n66), .ZN(
        npu_inst_pe_1_1_5_n89) );
  NAND2_X1 npu_inst_pe_1_1_5_U61 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_5_n44), .ZN(npu_inst_pe_1_1_5_n65) );
  OAI21_X1 npu_inst_pe_1_1_5_U60 ( .B1(npu_inst_pe_1_1_5_n61), .B2(
        npu_inst_pe_1_1_5_n44), .A(npu_inst_pe_1_1_5_n65), .ZN(
        npu_inst_pe_1_1_5_n88) );
  NAND2_X1 npu_inst_pe_1_1_5_U59 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_5_n40), .ZN(npu_inst_pe_1_1_5_n64) );
  OAI21_X1 npu_inst_pe_1_1_5_U58 ( .B1(npu_inst_pe_1_1_5_n63), .B2(
        npu_inst_pe_1_1_5_n40), .A(npu_inst_pe_1_1_5_n64), .ZN(
        npu_inst_pe_1_1_5_n87) );
  NAND2_X1 npu_inst_pe_1_1_5_U57 ( .A1(npu_inst_pe_1_1_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_5_n40), .ZN(npu_inst_pe_1_1_5_n62) );
  OAI21_X1 npu_inst_pe_1_1_5_U56 ( .B1(npu_inst_pe_1_1_5_n61), .B2(
        npu_inst_pe_1_1_5_n40), .A(npu_inst_pe_1_1_5_n62), .ZN(
        npu_inst_pe_1_1_5_n86) );
  AOI22_X1 npu_inst_pe_1_1_5_U55 ( .A1(npu_inst_pe_1_1_5_n38), .A2(
        npu_inst_int_data_y_2__5__0_), .B1(npu_inst_pe_1_1_5_n113), .B2(
        npu_inst_pe_1_1_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_5_n37) );
  INV_X1 npu_inst_pe_1_1_5_U54 ( .A(npu_inst_pe_1_1_5_n37), .ZN(
        npu_inst_pe_1_1_5_n112) );
  AND2_X1 npu_inst_pe_1_1_5_U53 ( .A1(npu_inst_n41), .A2(npu_inst_pe_1_1_5_N94), .ZN(npu_inst_int_data_y_1__5__1_) );
  AOI222_X1 npu_inst_pe_1_1_5_U52 ( .A1(npu_inst_int_data_res_2__5__0_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N73), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N65), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n84) );
  INV_X1 npu_inst_pe_1_1_5_U51 ( .A(npu_inst_pe_1_1_5_n84), .ZN(
        npu_inst_pe_1_1_5_n100) );
  AOI222_X1 npu_inst_pe_1_1_5_U50 ( .A1(npu_inst_pe_1_1_5_n1), .A2(
        npu_inst_int_data_res_2__5__7_), .B1(npu_inst_pe_1_1_5_N80), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N72), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n75) );
  INV_X1 npu_inst_pe_1_1_5_U49 ( .A(npu_inst_pe_1_1_5_n75), .ZN(
        npu_inst_pe_1_1_5_n32) );
  AOI222_X1 npu_inst_pe_1_1_5_U48 ( .A1(npu_inst_int_data_res_2__5__1_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N74), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N66), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n83) );
  INV_X1 npu_inst_pe_1_1_5_U47 ( .A(npu_inst_pe_1_1_5_n83), .ZN(
        npu_inst_pe_1_1_5_n99) );
  AOI222_X1 npu_inst_pe_1_1_5_U46 ( .A1(npu_inst_int_data_res_2__5__3_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N76), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N68), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n81) );
  INV_X1 npu_inst_pe_1_1_5_U45 ( .A(npu_inst_pe_1_1_5_n81), .ZN(
        npu_inst_pe_1_1_5_n36) );
  AOI222_X1 npu_inst_pe_1_1_5_U44 ( .A1(npu_inst_int_data_res_2__5__4_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N77), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N69), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n80) );
  INV_X1 npu_inst_pe_1_1_5_U43 ( .A(npu_inst_pe_1_1_5_n80), .ZN(
        npu_inst_pe_1_1_5_n35) );
  AOI222_X1 npu_inst_pe_1_1_5_U42 ( .A1(npu_inst_int_data_res_2__5__5_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N78), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N70), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n79) );
  INV_X1 npu_inst_pe_1_1_5_U41 ( .A(npu_inst_pe_1_1_5_n79), .ZN(
        npu_inst_pe_1_1_5_n34) );
  AOI222_X1 npu_inst_pe_1_1_5_U40 ( .A1(npu_inst_int_data_res_2__5__6_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N79), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N71), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n78) );
  INV_X1 npu_inst_pe_1_1_5_U39 ( .A(npu_inst_pe_1_1_5_n78), .ZN(
        npu_inst_pe_1_1_5_n33) );
  AND2_X1 npu_inst_pe_1_1_5_U38 ( .A1(npu_inst_int_data_x_1__5__1_), .A2(
        npu_inst_pe_1_1_5_int_q_weight_1_), .ZN(npu_inst_pe_1_1_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_5_U37 ( .A1(npu_inst_int_data_x_1__5__0_), .A2(
        npu_inst_pe_1_1_5_int_q_weight_1_), .ZN(npu_inst_pe_1_1_5_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_1_5_U36 ( .A(npu_inst_pe_1_1_5_int_data_1_), .ZN(
        npu_inst_pe_1_1_5_n13) );
  NOR3_X1 npu_inst_pe_1_1_5_U35 ( .A1(npu_inst_pe_1_1_5_n26), .A2(npu_inst_n41), .A3(npu_inst_int_ckg[50]), .ZN(npu_inst_pe_1_1_5_n85) );
  OR2_X1 npu_inst_pe_1_1_5_U34 ( .A1(npu_inst_pe_1_1_5_n85), .A2(
        npu_inst_pe_1_1_5_n1), .ZN(npu_inst_pe_1_1_5_N84) );
  AOI222_X1 npu_inst_pe_1_1_5_U33 ( .A1(npu_inst_int_data_res_2__5__2_), .A2(
        npu_inst_pe_1_1_5_n1), .B1(npu_inst_pe_1_1_5_N75), .B2(
        npu_inst_pe_1_1_5_n76), .C1(npu_inst_pe_1_1_5_N67), .C2(
        npu_inst_pe_1_1_5_n77), .ZN(npu_inst_pe_1_1_5_n82) );
  INV_X1 npu_inst_pe_1_1_5_U32 ( .A(npu_inst_pe_1_1_5_n82), .ZN(
        npu_inst_pe_1_1_5_n98) );
  AOI22_X1 npu_inst_pe_1_1_5_U31 ( .A1(npu_inst_n41), .A2(
        npu_inst_int_data_y_2__5__1_), .B1(npu_inst_pe_1_1_5_n2), .B2(
        npu_inst_int_data_x_1__6__1_), .ZN(npu_inst_pe_1_1_5_n63) );
  AOI22_X1 npu_inst_pe_1_1_5_U30 ( .A1(npu_inst_n41), .A2(
        npu_inst_int_data_y_2__5__0_), .B1(npu_inst_pe_1_1_5_n2), .B2(
        npu_inst_int_data_x_1__6__0_), .ZN(npu_inst_pe_1_1_5_n61) );
  INV_X1 npu_inst_pe_1_1_5_U29 ( .A(npu_inst_pe_1_1_5_int_data_0_), .ZN(
        npu_inst_pe_1_1_5_n12) );
  INV_X1 npu_inst_pe_1_1_5_U28 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_1_5_n4)
         );
  OR3_X1 npu_inst_pe_1_1_5_U27 ( .A1(npu_inst_pe_1_1_5_n5), .A2(
        npu_inst_pe_1_1_5_n7), .A3(npu_inst_pe_1_1_5_n4), .ZN(
        npu_inst_pe_1_1_5_n56) );
  OR3_X1 npu_inst_pe_1_1_5_U26 ( .A1(npu_inst_pe_1_1_5_n4), .A2(
        npu_inst_pe_1_1_5_n7), .A3(npu_inst_pe_1_1_5_n6), .ZN(
        npu_inst_pe_1_1_5_n48) );
  INV_X1 npu_inst_pe_1_1_5_U25 ( .A(npu_inst_pe_1_1_5_n4), .ZN(
        npu_inst_pe_1_1_5_n3) );
  OR3_X1 npu_inst_pe_1_1_5_U24 ( .A1(npu_inst_pe_1_1_5_n3), .A2(
        npu_inst_pe_1_1_5_n7), .A3(npu_inst_pe_1_1_5_n6), .ZN(
        npu_inst_pe_1_1_5_n52) );
  OR3_X1 npu_inst_pe_1_1_5_U23 ( .A1(npu_inst_pe_1_1_5_n5), .A2(
        npu_inst_pe_1_1_5_n7), .A3(npu_inst_pe_1_1_5_n3), .ZN(
        npu_inst_pe_1_1_5_n60) );
  BUF_X1 npu_inst_pe_1_1_5_U22 ( .A(npu_inst_n27), .Z(npu_inst_pe_1_1_5_n1) );
  NOR2_X1 npu_inst_pe_1_1_5_U21 ( .A1(npu_inst_pe_1_1_5_n60), .A2(
        npu_inst_pe_1_1_5_n2), .ZN(npu_inst_pe_1_1_5_n58) );
  NOR2_X1 npu_inst_pe_1_1_5_U20 ( .A1(npu_inst_pe_1_1_5_n56), .A2(
        npu_inst_pe_1_1_5_n2), .ZN(npu_inst_pe_1_1_5_n54) );
  NOR2_X1 npu_inst_pe_1_1_5_U19 ( .A1(npu_inst_pe_1_1_5_n52), .A2(
        npu_inst_pe_1_1_5_n2), .ZN(npu_inst_pe_1_1_5_n50) );
  NOR2_X1 npu_inst_pe_1_1_5_U18 ( .A1(npu_inst_pe_1_1_5_n48), .A2(
        npu_inst_pe_1_1_5_n2), .ZN(npu_inst_pe_1_1_5_n46) );
  NOR2_X1 npu_inst_pe_1_1_5_U17 ( .A1(npu_inst_pe_1_1_5_n40), .A2(
        npu_inst_pe_1_1_5_n2), .ZN(npu_inst_pe_1_1_5_n38) );
  NOR2_X1 npu_inst_pe_1_1_5_U16 ( .A1(npu_inst_pe_1_1_5_n44), .A2(
        npu_inst_pe_1_1_5_n2), .ZN(npu_inst_pe_1_1_5_n42) );
  BUF_X1 npu_inst_pe_1_1_5_U15 ( .A(npu_inst_n86), .Z(npu_inst_pe_1_1_5_n7) );
  INV_X1 npu_inst_pe_1_1_5_U14 ( .A(npu_inst_n108), .ZN(npu_inst_pe_1_1_5_n11)
         );
  INV_X1 npu_inst_pe_1_1_5_U13 ( .A(npu_inst_pe_1_1_5_n38), .ZN(
        npu_inst_pe_1_1_5_n113) );
  INV_X1 npu_inst_pe_1_1_5_U12 ( .A(npu_inst_pe_1_1_5_n58), .ZN(
        npu_inst_pe_1_1_5_n118) );
  INV_X1 npu_inst_pe_1_1_5_U11 ( .A(npu_inst_pe_1_1_5_n54), .ZN(
        npu_inst_pe_1_1_5_n117) );
  INV_X1 npu_inst_pe_1_1_5_U10 ( .A(npu_inst_pe_1_1_5_n50), .ZN(
        npu_inst_pe_1_1_5_n116) );
  INV_X1 npu_inst_pe_1_1_5_U9 ( .A(npu_inst_pe_1_1_5_n46), .ZN(
        npu_inst_pe_1_1_5_n115) );
  INV_X1 npu_inst_pe_1_1_5_U8 ( .A(npu_inst_pe_1_1_5_n42), .ZN(
        npu_inst_pe_1_1_5_n114) );
  BUF_X1 npu_inst_pe_1_1_5_U7 ( .A(npu_inst_pe_1_1_5_n11), .Z(
        npu_inst_pe_1_1_5_n10) );
  BUF_X1 npu_inst_pe_1_1_5_U6 ( .A(npu_inst_pe_1_1_5_n11), .Z(
        npu_inst_pe_1_1_5_n9) );
  BUF_X1 npu_inst_pe_1_1_5_U5 ( .A(npu_inst_pe_1_1_5_n11), .Z(
        npu_inst_pe_1_1_5_n8) );
  NOR2_X1 npu_inst_pe_1_1_5_U4 ( .A1(npu_inst_pe_1_1_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_5_n1), .ZN(npu_inst_pe_1_1_5_n76) );
  NOR2_X1 npu_inst_pe_1_1_5_U3 ( .A1(npu_inst_pe_1_1_5_n27), .A2(
        npu_inst_pe_1_1_5_n1), .ZN(npu_inst_pe_1_1_5_n77) );
  FA_X1 npu_inst_pe_1_1_5_sub_77_U2_1 ( .A(npu_inst_int_data_res_1__5__1_), 
        .B(npu_inst_pe_1_1_5_n13), .CI(npu_inst_pe_1_1_5_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_1_5_sub_77_carry_2_), .S(npu_inst_pe_1_1_5_N66) );
  FA_X1 npu_inst_pe_1_1_5_add_79_U1_1 ( .A(npu_inst_int_data_res_1__5__1_), 
        .B(npu_inst_pe_1_1_5_int_data_1_), .CI(
        npu_inst_pe_1_1_5_add_79_carry_1_), .CO(
        npu_inst_pe_1_1_5_add_79_carry_2_), .S(npu_inst_pe_1_1_5_N74) );
  NAND3_X1 npu_inst_pe_1_1_5_U101 ( .A1(npu_inst_pe_1_1_5_n4), .A2(
        npu_inst_pe_1_1_5_n6), .A3(npu_inst_pe_1_1_5_n7), .ZN(
        npu_inst_pe_1_1_5_n44) );
  NAND3_X1 npu_inst_pe_1_1_5_U100 ( .A1(npu_inst_pe_1_1_5_n3), .A2(
        npu_inst_pe_1_1_5_n6), .A3(npu_inst_pe_1_1_5_n7), .ZN(
        npu_inst_pe_1_1_5_n40) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_5_n33), .CK(
        npu_inst_pe_1_1_5_net4179), .RN(npu_inst_pe_1_1_5_n8), .Q(
        npu_inst_int_data_res_1__5__6_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_5_n34), .CK(
        npu_inst_pe_1_1_5_net4179), .RN(npu_inst_pe_1_1_5_n8), .Q(
        npu_inst_int_data_res_1__5__5_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_5_n35), .CK(
        npu_inst_pe_1_1_5_net4179), .RN(npu_inst_pe_1_1_5_n8), .Q(
        npu_inst_int_data_res_1__5__4_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_5_n36), .CK(
        npu_inst_pe_1_1_5_net4179), .RN(npu_inst_pe_1_1_5_n8), .Q(
        npu_inst_int_data_res_1__5__3_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_5_n98), .CK(
        npu_inst_pe_1_1_5_net4179), .RN(npu_inst_pe_1_1_5_n8), .Q(
        npu_inst_int_data_res_1__5__2_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_5_n99), .CK(
        npu_inst_pe_1_1_5_net4179), .RN(npu_inst_pe_1_1_5_n8), .Q(
        npu_inst_int_data_res_1__5__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_5_n32), .CK(
        npu_inst_pe_1_1_5_net4179), .RN(npu_inst_pe_1_1_5_n8), .Q(
        npu_inst_int_data_res_1__5__7_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_5_n100), 
        .CK(npu_inst_pe_1_1_5_net4179), .RN(npu_inst_pe_1_1_5_n8), .Q(
        npu_inst_int_data_res_1__5__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_weight_reg_0_ ( .D(npu_inst_n94), .CK(
        npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n8), .Q(
        npu_inst_pe_1_1_5_int_q_weight_0_), .QN(npu_inst_pe_1_1_5_n27) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_weight_reg_1_ ( .D(npu_inst_n100), .CK(
        npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n8), .Q(
        npu_inst_pe_1_1_5_int_q_weight_1_), .QN(npu_inst_pe_1_1_5_n26) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_5_n112), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n8), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_5_n106), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n8), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_5_n111), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_5_n105), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_5_n110), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_5_n104), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_5_n109), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_5_n103), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_5_n108), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_5_n102), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_5_n107), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_5_n101), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_5_n86), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_5_n87), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n9), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_5_n88), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_5_n89), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_5_n90), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_5_n91), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_5_n92), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_5_n93), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_5_n94), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_5_n95), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_5_n96), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_5_n97), 
        .CK(npu_inst_pe_1_1_5_net4185), .RN(npu_inst_pe_1_1_5_n10), .Q(
        npu_inst_pe_1_1_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_5_net4179) );
  CLKGATETST_X1 npu_inst_pe_1_1_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n47), .SE(1'b0), .GCK(npu_inst_pe_1_1_5_net4185) );
  MUX2_X1 npu_inst_pe_1_1_6_U153 ( .A(npu_inst_pe_1_1_6_n31), .B(
        npu_inst_pe_1_1_6_n28), .S(npu_inst_pe_1_1_6_n7), .Z(
        npu_inst_pe_1_1_6_N93) );
  MUX2_X1 npu_inst_pe_1_1_6_U152 ( .A(npu_inst_pe_1_1_6_n30), .B(
        npu_inst_pe_1_1_6_n29), .S(npu_inst_pe_1_1_6_n5), .Z(
        npu_inst_pe_1_1_6_n31) );
  MUX2_X1 npu_inst_pe_1_1_6_U151 ( .A(npu_inst_pe_1_1_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_6_n3), .Z(
        npu_inst_pe_1_1_6_n30) );
  MUX2_X1 npu_inst_pe_1_1_6_U150 ( .A(npu_inst_pe_1_1_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_6_n3), .Z(
        npu_inst_pe_1_1_6_n29) );
  MUX2_X1 npu_inst_pe_1_1_6_U149 ( .A(npu_inst_pe_1_1_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_6_n3), .Z(
        npu_inst_pe_1_1_6_n28) );
  MUX2_X1 npu_inst_pe_1_1_6_U148 ( .A(npu_inst_pe_1_1_6_n25), .B(
        npu_inst_pe_1_1_6_n22), .S(npu_inst_pe_1_1_6_n7), .Z(
        npu_inst_pe_1_1_6_N94) );
  MUX2_X1 npu_inst_pe_1_1_6_U147 ( .A(npu_inst_pe_1_1_6_n24), .B(
        npu_inst_pe_1_1_6_n23), .S(npu_inst_pe_1_1_6_n5), .Z(
        npu_inst_pe_1_1_6_n25) );
  MUX2_X1 npu_inst_pe_1_1_6_U146 ( .A(npu_inst_pe_1_1_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_6_n3), .Z(
        npu_inst_pe_1_1_6_n24) );
  MUX2_X1 npu_inst_pe_1_1_6_U145 ( .A(npu_inst_pe_1_1_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_6_n3), .Z(
        npu_inst_pe_1_1_6_n23) );
  MUX2_X1 npu_inst_pe_1_1_6_U144 ( .A(npu_inst_pe_1_1_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_6_n3), .Z(
        npu_inst_pe_1_1_6_n22) );
  MUX2_X1 npu_inst_pe_1_1_6_U143 ( .A(npu_inst_pe_1_1_6_n21), .B(
        npu_inst_pe_1_1_6_n18), .S(npu_inst_pe_1_1_6_n7), .Z(
        npu_inst_int_data_x_1__6__1_) );
  MUX2_X1 npu_inst_pe_1_1_6_U142 ( .A(npu_inst_pe_1_1_6_n20), .B(
        npu_inst_pe_1_1_6_n19), .S(npu_inst_pe_1_1_6_n5), .Z(
        npu_inst_pe_1_1_6_n21) );
  MUX2_X1 npu_inst_pe_1_1_6_U141 ( .A(npu_inst_pe_1_1_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_6_n3), .Z(
        npu_inst_pe_1_1_6_n20) );
  MUX2_X1 npu_inst_pe_1_1_6_U140 ( .A(npu_inst_pe_1_1_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_6_n3), .Z(
        npu_inst_pe_1_1_6_n19) );
  MUX2_X1 npu_inst_pe_1_1_6_U139 ( .A(npu_inst_pe_1_1_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_6_n3), .Z(
        npu_inst_pe_1_1_6_n18) );
  MUX2_X1 npu_inst_pe_1_1_6_U138 ( .A(npu_inst_pe_1_1_6_n17), .B(
        npu_inst_pe_1_1_6_n14), .S(npu_inst_pe_1_1_6_n7), .Z(
        npu_inst_int_data_x_1__6__0_) );
  MUX2_X1 npu_inst_pe_1_1_6_U137 ( .A(npu_inst_pe_1_1_6_n16), .B(
        npu_inst_pe_1_1_6_n15), .S(npu_inst_pe_1_1_6_n5), .Z(
        npu_inst_pe_1_1_6_n17) );
  MUX2_X1 npu_inst_pe_1_1_6_U136 ( .A(npu_inst_pe_1_1_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_6_n3), .Z(
        npu_inst_pe_1_1_6_n16) );
  MUX2_X1 npu_inst_pe_1_1_6_U135 ( .A(npu_inst_pe_1_1_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_6_n3), .Z(
        npu_inst_pe_1_1_6_n15) );
  MUX2_X1 npu_inst_pe_1_1_6_U134 ( .A(npu_inst_pe_1_1_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_6_n3), .Z(
        npu_inst_pe_1_1_6_n14) );
  XOR2_X1 npu_inst_pe_1_1_6_U133 ( .A(npu_inst_pe_1_1_6_int_data_0_), .B(
        npu_inst_int_data_res_1__6__0_), .Z(npu_inst_pe_1_1_6_N73) );
  AND2_X1 npu_inst_pe_1_1_6_U132 ( .A1(npu_inst_int_data_res_1__6__0_), .A2(
        npu_inst_pe_1_1_6_int_data_0_), .ZN(npu_inst_pe_1_1_6_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_6_U131 ( .A(npu_inst_int_data_res_1__6__0_), .B(
        npu_inst_pe_1_1_6_n12), .ZN(npu_inst_pe_1_1_6_N65) );
  OR2_X1 npu_inst_pe_1_1_6_U130 ( .A1(npu_inst_pe_1_1_6_n12), .A2(
        npu_inst_int_data_res_1__6__0_), .ZN(npu_inst_pe_1_1_6_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_6_U129 ( .A(npu_inst_int_data_res_1__6__2_), .B(
        npu_inst_pe_1_1_6_add_79_carry_2_), .Z(npu_inst_pe_1_1_6_N75) );
  AND2_X1 npu_inst_pe_1_1_6_U128 ( .A1(npu_inst_pe_1_1_6_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_1__6__2_), .ZN(
        npu_inst_pe_1_1_6_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_6_U127 ( .A(npu_inst_int_data_res_1__6__3_), .B(
        npu_inst_pe_1_1_6_add_79_carry_3_), .Z(npu_inst_pe_1_1_6_N76) );
  AND2_X1 npu_inst_pe_1_1_6_U126 ( .A1(npu_inst_pe_1_1_6_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_1__6__3_), .ZN(
        npu_inst_pe_1_1_6_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_6_U125 ( .A(npu_inst_int_data_res_1__6__4_), .B(
        npu_inst_pe_1_1_6_add_79_carry_4_), .Z(npu_inst_pe_1_1_6_N77) );
  AND2_X1 npu_inst_pe_1_1_6_U124 ( .A1(npu_inst_pe_1_1_6_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_1__6__4_), .ZN(
        npu_inst_pe_1_1_6_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_6_U123 ( .A(npu_inst_int_data_res_1__6__5_), .B(
        npu_inst_pe_1_1_6_add_79_carry_5_), .Z(npu_inst_pe_1_1_6_N78) );
  AND2_X1 npu_inst_pe_1_1_6_U122 ( .A1(npu_inst_pe_1_1_6_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_1__6__5_), .ZN(
        npu_inst_pe_1_1_6_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_6_U121 ( .A(npu_inst_int_data_res_1__6__6_), .B(
        npu_inst_pe_1_1_6_add_79_carry_6_), .Z(npu_inst_pe_1_1_6_N79) );
  AND2_X1 npu_inst_pe_1_1_6_U120 ( .A1(npu_inst_pe_1_1_6_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_1__6__6_), .ZN(
        npu_inst_pe_1_1_6_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_6_U119 ( .A(npu_inst_int_data_res_1__6__7_), .B(
        npu_inst_pe_1_1_6_add_79_carry_7_), .Z(npu_inst_pe_1_1_6_N80) );
  XNOR2_X1 npu_inst_pe_1_1_6_U118 ( .A(npu_inst_pe_1_1_6_sub_77_carry_2_), .B(
        npu_inst_int_data_res_1__6__2_), .ZN(npu_inst_pe_1_1_6_N67) );
  OR2_X1 npu_inst_pe_1_1_6_U117 ( .A1(npu_inst_int_data_res_1__6__2_), .A2(
        npu_inst_pe_1_1_6_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_1_6_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_6_U116 ( .A(npu_inst_pe_1_1_6_sub_77_carry_3_), .B(
        npu_inst_int_data_res_1__6__3_), .ZN(npu_inst_pe_1_1_6_N68) );
  OR2_X1 npu_inst_pe_1_1_6_U115 ( .A1(npu_inst_int_data_res_1__6__3_), .A2(
        npu_inst_pe_1_1_6_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_1_6_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_6_U114 ( .A(npu_inst_pe_1_1_6_sub_77_carry_4_), .B(
        npu_inst_int_data_res_1__6__4_), .ZN(npu_inst_pe_1_1_6_N69) );
  OR2_X1 npu_inst_pe_1_1_6_U113 ( .A1(npu_inst_int_data_res_1__6__4_), .A2(
        npu_inst_pe_1_1_6_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_1_6_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_6_U112 ( .A(npu_inst_pe_1_1_6_sub_77_carry_5_), .B(
        npu_inst_int_data_res_1__6__5_), .ZN(npu_inst_pe_1_1_6_N70) );
  OR2_X1 npu_inst_pe_1_1_6_U111 ( .A1(npu_inst_int_data_res_1__6__5_), .A2(
        npu_inst_pe_1_1_6_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_1_6_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_6_U110 ( .A(npu_inst_pe_1_1_6_sub_77_carry_6_), .B(
        npu_inst_int_data_res_1__6__6_), .ZN(npu_inst_pe_1_1_6_N71) );
  OR2_X1 npu_inst_pe_1_1_6_U109 ( .A1(npu_inst_int_data_res_1__6__6_), .A2(
        npu_inst_pe_1_1_6_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_1_6_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_6_U108 ( .A(npu_inst_int_data_res_1__6__7_), .B(
        npu_inst_pe_1_1_6_sub_77_carry_7_), .ZN(npu_inst_pe_1_1_6_N72) );
  INV_X1 npu_inst_pe_1_1_6_U107 ( .A(npu_inst_n61), .ZN(npu_inst_pe_1_1_6_n6)
         );
  INV_X1 npu_inst_pe_1_1_6_U106 ( .A(npu_inst_pe_1_1_6_n6), .ZN(
        npu_inst_pe_1_1_6_n5) );
  INV_X1 npu_inst_pe_1_1_6_U105 ( .A(npu_inst_n41), .ZN(npu_inst_pe_1_1_6_n2)
         );
  AOI22_X1 npu_inst_pe_1_1_6_U104 ( .A1(npu_inst_int_data_y_2__6__0_), .A2(
        npu_inst_pe_1_1_6_n58), .B1(npu_inst_pe_1_1_6_n118), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_6_n57) );
  INV_X1 npu_inst_pe_1_1_6_U103 ( .A(npu_inst_pe_1_1_6_n57), .ZN(
        npu_inst_pe_1_1_6_n107) );
  AOI22_X1 npu_inst_pe_1_1_6_U102 ( .A1(npu_inst_int_data_y_2__6__0_), .A2(
        npu_inst_pe_1_1_6_n54), .B1(npu_inst_pe_1_1_6_n117), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_6_n53) );
  INV_X1 npu_inst_pe_1_1_6_U99 ( .A(npu_inst_pe_1_1_6_n53), .ZN(
        npu_inst_pe_1_1_6_n108) );
  AOI22_X1 npu_inst_pe_1_1_6_U98 ( .A1(npu_inst_int_data_y_2__6__0_), .A2(
        npu_inst_pe_1_1_6_n50), .B1(npu_inst_pe_1_1_6_n116), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_6_n49) );
  INV_X1 npu_inst_pe_1_1_6_U97 ( .A(npu_inst_pe_1_1_6_n49), .ZN(
        npu_inst_pe_1_1_6_n109) );
  AOI22_X1 npu_inst_pe_1_1_6_U96 ( .A1(npu_inst_int_data_y_2__6__0_), .A2(
        npu_inst_pe_1_1_6_n46), .B1(npu_inst_pe_1_1_6_n115), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_6_n45) );
  INV_X1 npu_inst_pe_1_1_6_U95 ( .A(npu_inst_pe_1_1_6_n45), .ZN(
        npu_inst_pe_1_1_6_n110) );
  AOI22_X1 npu_inst_pe_1_1_6_U94 ( .A1(npu_inst_int_data_y_2__6__0_), .A2(
        npu_inst_pe_1_1_6_n42), .B1(npu_inst_pe_1_1_6_n114), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_6_n41) );
  INV_X1 npu_inst_pe_1_1_6_U93 ( .A(npu_inst_pe_1_1_6_n41), .ZN(
        npu_inst_pe_1_1_6_n111) );
  AOI22_X1 npu_inst_pe_1_1_6_U92 ( .A1(npu_inst_int_data_y_2__6__1_), .A2(
        npu_inst_pe_1_1_6_n58), .B1(npu_inst_pe_1_1_6_n118), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_6_n59) );
  INV_X1 npu_inst_pe_1_1_6_U91 ( .A(npu_inst_pe_1_1_6_n59), .ZN(
        npu_inst_pe_1_1_6_n101) );
  AOI22_X1 npu_inst_pe_1_1_6_U90 ( .A1(npu_inst_int_data_y_2__6__1_), .A2(
        npu_inst_pe_1_1_6_n54), .B1(npu_inst_pe_1_1_6_n117), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_6_n55) );
  INV_X1 npu_inst_pe_1_1_6_U89 ( .A(npu_inst_pe_1_1_6_n55), .ZN(
        npu_inst_pe_1_1_6_n102) );
  AOI22_X1 npu_inst_pe_1_1_6_U88 ( .A1(npu_inst_int_data_y_2__6__1_), .A2(
        npu_inst_pe_1_1_6_n50), .B1(npu_inst_pe_1_1_6_n116), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_6_n51) );
  INV_X1 npu_inst_pe_1_1_6_U87 ( .A(npu_inst_pe_1_1_6_n51), .ZN(
        npu_inst_pe_1_1_6_n103) );
  AOI22_X1 npu_inst_pe_1_1_6_U86 ( .A1(npu_inst_int_data_y_2__6__1_), .A2(
        npu_inst_pe_1_1_6_n46), .B1(npu_inst_pe_1_1_6_n115), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_6_n47) );
  INV_X1 npu_inst_pe_1_1_6_U85 ( .A(npu_inst_pe_1_1_6_n47), .ZN(
        npu_inst_pe_1_1_6_n104) );
  AOI22_X1 npu_inst_pe_1_1_6_U84 ( .A1(npu_inst_int_data_y_2__6__1_), .A2(
        npu_inst_pe_1_1_6_n42), .B1(npu_inst_pe_1_1_6_n114), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_6_n43) );
  INV_X1 npu_inst_pe_1_1_6_U83 ( .A(npu_inst_pe_1_1_6_n43), .ZN(
        npu_inst_pe_1_1_6_n105) );
  AOI22_X1 npu_inst_pe_1_1_6_U82 ( .A1(npu_inst_pe_1_1_6_n38), .A2(
        npu_inst_int_data_y_2__6__1_), .B1(npu_inst_pe_1_1_6_n113), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_6_n39) );
  INV_X1 npu_inst_pe_1_1_6_U81 ( .A(npu_inst_pe_1_1_6_n39), .ZN(
        npu_inst_pe_1_1_6_n106) );
  AND2_X1 npu_inst_pe_1_1_6_U80 ( .A1(npu_inst_pe_1_1_6_N93), .A2(npu_inst_n41), .ZN(npu_inst_int_data_y_1__6__0_) );
  NAND2_X1 npu_inst_pe_1_1_6_U79 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_6_n60), .ZN(npu_inst_pe_1_1_6_n74) );
  OAI21_X1 npu_inst_pe_1_1_6_U78 ( .B1(npu_inst_pe_1_1_6_n63), .B2(
        npu_inst_pe_1_1_6_n60), .A(npu_inst_pe_1_1_6_n74), .ZN(
        npu_inst_pe_1_1_6_n97) );
  NAND2_X1 npu_inst_pe_1_1_6_U77 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_6_n60), .ZN(npu_inst_pe_1_1_6_n73) );
  OAI21_X1 npu_inst_pe_1_1_6_U76 ( .B1(npu_inst_pe_1_1_6_n61), .B2(
        npu_inst_pe_1_1_6_n60), .A(npu_inst_pe_1_1_6_n73), .ZN(
        npu_inst_pe_1_1_6_n96) );
  NAND2_X1 npu_inst_pe_1_1_6_U75 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_6_n56), .ZN(npu_inst_pe_1_1_6_n72) );
  OAI21_X1 npu_inst_pe_1_1_6_U74 ( .B1(npu_inst_pe_1_1_6_n63), .B2(
        npu_inst_pe_1_1_6_n56), .A(npu_inst_pe_1_1_6_n72), .ZN(
        npu_inst_pe_1_1_6_n95) );
  NAND2_X1 npu_inst_pe_1_1_6_U73 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_6_n56), .ZN(npu_inst_pe_1_1_6_n71) );
  OAI21_X1 npu_inst_pe_1_1_6_U72 ( .B1(npu_inst_pe_1_1_6_n61), .B2(
        npu_inst_pe_1_1_6_n56), .A(npu_inst_pe_1_1_6_n71), .ZN(
        npu_inst_pe_1_1_6_n94) );
  NAND2_X1 npu_inst_pe_1_1_6_U71 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_6_n52), .ZN(npu_inst_pe_1_1_6_n70) );
  OAI21_X1 npu_inst_pe_1_1_6_U70 ( .B1(npu_inst_pe_1_1_6_n63), .B2(
        npu_inst_pe_1_1_6_n52), .A(npu_inst_pe_1_1_6_n70), .ZN(
        npu_inst_pe_1_1_6_n93) );
  NAND2_X1 npu_inst_pe_1_1_6_U69 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_6_n52), .ZN(npu_inst_pe_1_1_6_n69) );
  OAI21_X1 npu_inst_pe_1_1_6_U68 ( .B1(npu_inst_pe_1_1_6_n61), .B2(
        npu_inst_pe_1_1_6_n52), .A(npu_inst_pe_1_1_6_n69), .ZN(
        npu_inst_pe_1_1_6_n92) );
  NAND2_X1 npu_inst_pe_1_1_6_U67 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_6_n48), .ZN(npu_inst_pe_1_1_6_n68) );
  OAI21_X1 npu_inst_pe_1_1_6_U66 ( .B1(npu_inst_pe_1_1_6_n63), .B2(
        npu_inst_pe_1_1_6_n48), .A(npu_inst_pe_1_1_6_n68), .ZN(
        npu_inst_pe_1_1_6_n91) );
  NAND2_X1 npu_inst_pe_1_1_6_U65 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_6_n48), .ZN(npu_inst_pe_1_1_6_n67) );
  OAI21_X1 npu_inst_pe_1_1_6_U64 ( .B1(npu_inst_pe_1_1_6_n61), .B2(
        npu_inst_pe_1_1_6_n48), .A(npu_inst_pe_1_1_6_n67), .ZN(
        npu_inst_pe_1_1_6_n90) );
  NAND2_X1 npu_inst_pe_1_1_6_U63 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_6_n44), .ZN(npu_inst_pe_1_1_6_n66) );
  OAI21_X1 npu_inst_pe_1_1_6_U62 ( .B1(npu_inst_pe_1_1_6_n63), .B2(
        npu_inst_pe_1_1_6_n44), .A(npu_inst_pe_1_1_6_n66), .ZN(
        npu_inst_pe_1_1_6_n89) );
  NAND2_X1 npu_inst_pe_1_1_6_U61 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_6_n44), .ZN(npu_inst_pe_1_1_6_n65) );
  OAI21_X1 npu_inst_pe_1_1_6_U60 ( .B1(npu_inst_pe_1_1_6_n61), .B2(
        npu_inst_pe_1_1_6_n44), .A(npu_inst_pe_1_1_6_n65), .ZN(
        npu_inst_pe_1_1_6_n88) );
  NAND2_X1 npu_inst_pe_1_1_6_U59 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_6_n40), .ZN(npu_inst_pe_1_1_6_n64) );
  OAI21_X1 npu_inst_pe_1_1_6_U58 ( .B1(npu_inst_pe_1_1_6_n63), .B2(
        npu_inst_pe_1_1_6_n40), .A(npu_inst_pe_1_1_6_n64), .ZN(
        npu_inst_pe_1_1_6_n87) );
  NAND2_X1 npu_inst_pe_1_1_6_U57 ( .A1(npu_inst_pe_1_1_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_6_n40), .ZN(npu_inst_pe_1_1_6_n62) );
  OAI21_X1 npu_inst_pe_1_1_6_U56 ( .B1(npu_inst_pe_1_1_6_n61), .B2(
        npu_inst_pe_1_1_6_n40), .A(npu_inst_pe_1_1_6_n62), .ZN(
        npu_inst_pe_1_1_6_n86) );
  AOI22_X1 npu_inst_pe_1_1_6_U55 ( .A1(npu_inst_pe_1_1_6_n38), .A2(
        npu_inst_int_data_y_2__6__0_), .B1(npu_inst_pe_1_1_6_n113), .B2(
        npu_inst_pe_1_1_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_6_n37) );
  INV_X1 npu_inst_pe_1_1_6_U54 ( .A(npu_inst_pe_1_1_6_n37), .ZN(
        npu_inst_pe_1_1_6_n112) );
  AND2_X1 npu_inst_pe_1_1_6_U53 ( .A1(npu_inst_n41), .A2(npu_inst_pe_1_1_6_N94), .ZN(npu_inst_int_data_y_1__6__1_) );
  AOI222_X1 npu_inst_pe_1_1_6_U52 ( .A1(npu_inst_int_data_res_2__6__0_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N73), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N65), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n84) );
  INV_X1 npu_inst_pe_1_1_6_U51 ( .A(npu_inst_pe_1_1_6_n84), .ZN(
        npu_inst_pe_1_1_6_n100) );
  AOI222_X1 npu_inst_pe_1_1_6_U50 ( .A1(npu_inst_pe_1_1_6_n1), .A2(
        npu_inst_int_data_res_2__6__7_), .B1(npu_inst_pe_1_1_6_N80), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N72), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n75) );
  INV_X1 npu_inst_pe_1_1_6_U49 ( .A(npu_inst_pe_1_1_6_n75), .ZN(
        npu_inst_pe_1_1_6_n32) );
  AOI222_X1 npu_inst_pe_1_1_6_U48 ( .A1(npu_inst_int_data_res_2__6__1_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N74), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N66), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n83) );
  INV_X1 npu_inst_pe_1_1_6_U47 ( .A(npu_inst_pe_1_1_6_n83), .ZN(
        npu_inst_pe_1_1_6_n99) );
  AOI222_X1 npu_inst_pe_1_1_6_U46 ( .A1(npu_inst_int_data_res_2__6__3_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N76), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N68), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n81) );
  INV_X1 npu_inst_pe_1_1_6_U45 ( .A(npu_inst_pe_1_1_6_n81), .ZN(
        npu_inst_pe_1_1_6_n36) );
  AOI222_X1 npu_inst_pe_1_1_6_U44 ( .A1(npu_inst_int_data_res_2__6__4_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N77), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N69), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n80) );
  INV_X1 npu_inst_pe_1_1_6_U43 ( .A(npu_inst_pe_1_1_6_n80), .ZN(
        npu_inst_pe_1_1_6_n35) );
  AOI222_X1 npu_inst_pe_1_1_6_U42 ( .A1(npu_inst_int_data_res_2__6__5_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N78), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N70), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n79) );
  INV_X1 npu_inst_pe_1_1_6_U41 ( .A(npu_inst_pe_1_1_6_n79), .ZN(
        npu_inst_pe_1_1_6_n34) );
  AOI222_X1 npu_inst_pe_1_1_6_U40 ( .A1(npu_inst_int_data_res_2__6__6_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N79), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N71), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n78) );
  INV_X1 npu_inst_pe_1_1_6_U39 ( .A(npu_inst_pe_1_1_6_n78), .ZN(
        npu_inst_pe_1_1_6_n33) );
  AND2_X1 npu_inst_pe_1_1_6_U38 ( .A1(npu_inst_int_data_x_1__6__1_), .A2(
        npu_inst_pe_1_1_6_int_q_weight_1_), .ZN(npu_inst_pe_1_1_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_6_U37 ( .A1(npu_inst_int_data_x_1__6__0_), .A2(
        npu_inst_pe_1_1_6_int_q_weight_1_), .ZN(npu_inst_pe_1_1_6_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_1_6_U36 ( .A(npu_inst_pe_1_1_6_int_data_1_), .ZN(
        npu_inst_pe_1_1_6_n13) );
  NOR3_X1 npu_inst_pe_1_1_6_U35 ( .A1(npu_inst_pe_1_1_6_n26), .A2(npu_inst_n41), .A3(npu_inst_int_ckg[49]), .ZN(npu_inst_pe_1_1_6_n85) );
  OR2_X1 npu_inst_pe_1_1_6_U34 ( .A1(npu_inst_pe_1_1_6_n85), .A2(
        npu_inst_pe_1_1_6_n1), .ZN(npu_inst_pe_1_1_6_N84) );
  AOI222_X1 npu_inst_pe_1_1_6_U33 ( .A1(npu_inst_int_data_res_2__6__2_), .A2(
        npu_inst_pe_1_1_6_n1), .B1(npu_inst_pe_1_1_6_N75), .B2(
        npu_inst_pe_1_1_6_n76), .C1(npu_inst_pe_1_1_6_N67), .C2(
        npu_inst_pe_1_1_6_n77), .ZN(npu_inst_pe_1_1_6_n82) );
  INV_X1 npu_inst_pe_1_1_6_U32 ( .A(npu_inst_pe_1_1_6_n82), .ZN(
        npu_inst_pe_1_1_6_n98) );
  AOI22_X1 npu_inst_pe_1_1_6_U31 ( .A1(npu_inst_n41), .A2(
        npu_inst_int_data_y_2__6__1_), .B1(npu_inst_pe_1_1_6_n2), .B2(
        npu_inst_int_data_x_1__7__1_), .ZN(npu_inst_pe_1_1_6_n63) );
  AOI22_X1 npu_inst_pe_1_1_6_U30 ( .A1(npu_inst_n41), .A2(
        npu_inst_int_data_y_2__6__0_), .B1(npu_inst_pe_1_1_6_n2), .B2(
        npu_inst_int_data_x_1__7__0_), .ZN(npu_inst_pe_1_1_6_n61) );
  INV_X1 npu_inst_pe_1_1_6_U29 ( .A(npu_inst_pe_1_1_6_int_data_0_), .ZN(
        npu_inst_pe_1_1_6_n12) );
  INV_X1 npu_inst_pe_1_1_6_U28 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_1_6_n4)
         );
  OR3_X1 npu_inst_pe_1_1_6_U27 ( .A1(npu_inst_pe_1_1_6_n5), .A2(
        npu_inst_pe_1_1_6_n7), .A3(npu_inst_pe_1_1_6_n4), .ZN(
        npu_inst_pe_1_1_6_n56) );
  OR3_X1 npu_inst_pe_1_1_6_U26 ( .A1(npu_inst_pe_1_1_6_n4), .A2(
        npu_inst_pe_1_1_6_n7), .A3(npu_inst_pe_1_1_6_n6), .ZN(
        npu_inst_pe_1_1_6_n48) );
  INV_X1 npu_inst_pe_1_1_6_U25 ( .A(npu_inst_pe_1_1_6_n4), .ZN(
        npu_inst_pe_1_1_6_n3) );
  OR3_X1 npu_inst_pe_1_1_6_U24 ( .A1(npu_inst_pe_1_1_6_n3), .A2(
        npu_inst_pe_1_1_6_n7), .A3(npu_inst_pe_1_1_6_n6), .ZN(
        npu_inst_pe_1_1_6_n52) );
  OR3_X1 npu_inst_pe_1_1_6_U23 ( .A1(npu_inst_pe_1_1_6_n5), .A2(
        npu_inst_pe_1_1_6_n7), .A3(npu_inst_pe_1_1_6_n3), .ZN(
        npu_inst_pe_1_1_6_n60) );
  BUF_X1 npu_inst_pe_1_1_6_U22 ( .A(npu_inst_n27), .Z(npu_inst_pe_1_1_6_n1) );
  NOR2_X1 npu_inst_pe_1_1_6_U21 ( .A1(npu_inst_pe_1_1_6_n60), .A2(
        npu_inst_pe_1_1_6_n2), .ZN(npu_inst_pe_1_1_6_n58) );
  NOR2_X1 npu_inst_pe_1_1_6_U20 ( .A1(npu_inst_pe_1_1_6_n56), .A2(
        npu_inst_pe_1_1_6_n2), .ZN(npu_inst_pe_1_1_6_n54) );
  NOR2_X1 npu_inst_pe_1_1_6_U19 ( .A1(npu_inst_pe_1_1_6_n52), .A2(
        npu_inst_pe_1_1_6_n2), .ZN(npu_inst_pe_1_1_6_n50) );
  NOR2_X1 npu_inst_pe_1_1_6_U18 ( .A1(npu_inst_pe_1_1_6_n48), .A2(
        npu_inst_pe_1_1_6_n2), .ZN(npu_inst_pe_1_1_6_n46) );
  NOR2_X1 npu_inst_pe_1_1_6_U17 ( .A1(npu_inst_pe_1_1_6_n40), .A2(
        npu_inst_pe_1_1_6_n2), .ZN(npu_inst_pe_1_1_6_n38) );
  NOR2_X1 npu_inst_pe_1_1_6_U16 ( .A1(npu_inst_pe_1_1_6_n44), .A2(
        npu_inst_pe_1_1_6_n2), .ZN(npu_inst_pe_1_1_6_n42) );
  BUF_X1 npu_inst_pe_1_1_6_U15 ( .A(npu_inst_n86), .Z(npu_inst_pe_1_1_6_n7) );
  INV_X1 npu_inst_pe_1_1_6_U14 ( .A(npu_inst_n108), .ZN(npu_inst_pe_1_1_6_n11)
         );
  INV_X1 npu_inst_pe_1_1_6_U13 ( .A(npu_inst_pe_1_1_6_n38), .ZN(
        npu_inst_pe_1_1_6_n113) );
  INV_X1 npu_inst_pe_1_1_6_U12 ( .A(npu_inst_pe_1_1_6_n58), .ZN(
        npu_inst_pe_1_1_6_n118) );
  INV_X1 npu_inst_pe_1_1_6_U11 ( .A(npu_inst_pe_1_1_6_n54), .ZN(
        npu_inst_pe_1_1_6_n117) );
  INV_X1 npu_inst_pe_1_1_6_U10 ( .A(npu_inst_pe_1_1_6_n50), .ZN(
        npu_inst_pe_1_1_6_n116) );
  INV_X1 npu_inst_pe_1_1_6_U9 ( .A(npu_inst_pe_1_1_6_n46), .ZN(
        npu_inst_pe_1_1_6_n115) );
  INV_X1 npu_inst_pe_1_1_6_U8 ( .A(npu_inst_pe_1_1_6_n42), .ZN(
        npu_inst_pe_1_1_6_n114) );
  BUF_X1 npu_inst_pe_1_1_6_U7 ( .A(npu_inst_pe_1_1_6_n11), .Z(
        npu_inst_pe_1_1_6_n10) );
  BUF_X1 npu_inst_pe_1_1_6_U6 ( .A(npu_inst_pe_1_1_6_n11), .Z(
        npu_inst_pe_1_1_6_n9) );
  BUF_X1 npu_inst_pe_1_1_6_U5 ( .A(npu_inst_pe_1_1_6_n11), .Z(
        npu_inst_pe_1_1_6_n8) );
  NOR2_X1 npu_inst_pe_1_1_6_U4 ( .A1(npu_inst_pe_1_1_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_6_n1), .ZN(npu_inst_pe_1_1_6_n76) );
  NOR2_X1 npu_inst_pe_1_1_6_U3 ( .A1(npu_inst_pe_1_1_6_n27), .A2(
        npu_inst_pe_1_1_6_n1), .ZN(npu_inst_pe_1_1_6_n77) );
  FA_X1 npu_inst_pe_1_1_6_sub_77_U2_1 ( .A(npu_inst_int_data_res_1__6__1_), 
        .B(npu_inst_pe_1_1_6_n13), .CI(npu_inst_pe_1_1_6_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_1_6_sub_77_carry_2_), .S(npu_inst_pe_1_1_6_N66) );
  FA_X1 npu_inst_pe_1_1_6_add_79_U1_1 ( .A(npu_inst_int_data_res_1__6__1_), 
        .B(npu_inst_pe_1_1_6_int_data_1_), .CI(
        npu_inst_pe_1_1_6_add_79_carry_1_), .CO(
        npu_inst_pe_1_1_6_add_79_carry_2_), .S(npu_inst_pe_1_1_6_N74) );
  NAND3_X1 npu_inst_pe_1_1_6_U101 ( .A1(npu_inst_pe_1_1_6_n4), .A2(
        npu_inst_pe_1_1_6_n6), .A3(npu_inst_pe_1_1_6_n7), .ZN(
        npu_inst_pe_1_1_6_n44) );
  NAND3_X1 npu_inst_pe_1_1_6_U100 ( .A1(npu_inst_pe_1_1_6_n3), .A2(
        npu_inst_pe_1_1_6_n6), .A3(npu_inst_pe_1_1_6_n7), .ZN(
        npu_inst_pe_1_1_6_n40) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_6_n33), .CK(
        npu_inst_pe_1_1_6_net4156), .RN(npu_inst_pe_1_1_6_n8), .Q(
        npu_inst_int_data_res_1__6__6_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_6_n34), .CK(
        npu_inst_pe_1_1_6_net4156), .RN(npu_inst_pe_1_1_6_n8), .Q(
        npu_inst_int_data_res_1__6__5_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_6_n35), .CK(
        npu_inst_pe_1_1_6_net4156), .RN(npu_inst_pe_1_1_6_n8), .Q(
        npu_inst_int_data_res_1__6__4_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_6_n36), .CK(
        npu_inst_pe_1_1_6_net4156), .RN(npu_inst_pe_1_1_6_n8), .Q(
        npu_inst_int_data_res_1__6__3_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_6_n98), .CK(
        npu_inst_pe_1_1_6_net4156), .RN(npu_inst_pe_1_1_6_n8), .Q(
        npu_inst_int_data_res_1__6__2_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_6_n99), .CK(
        npu_inst_pe_1_1_6_net4156), .RN(npu_inst_pe_1_1_6_n8), .Q(
        npu_inst_int_data_res_1__6__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_6_n32), .CK(
        npu_inst_pe_1_1_6_net4156), .RN(npu_inst_pe_1_1_6_n8), .Q(
        npu_inst_int_data_res_1__6__7_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_6_n100), 
        .CK(npu_inst_pe_1_1_6_net4156), .RN(npu_inst_pe_1_1_6_n8), .Q(
        npu_inst_int_data_res_1__6__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_weight_reg_0_ ( .D(npu_inst_n94), .CK(
        npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n8), .Q(
        npu_inst_pe_1_1_6_int_q_weight_0_), .QN(npu_inst_pe_1_1_6_n27) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_weight_reg_1_ ( .D(npu_inst_n100), .CK(
        npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n8), .Q(
        npu_inst_pe_1_1_6_int_q_weight_1_), .QN(npu_inst_pe_1_1_6_n26) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_6_n112), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n8), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_6_n106), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n8), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_6_n111), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_6_n105), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_6_n110), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_6_n104), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_6_n109), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_6_n103), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_6_n108), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_6_n102), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_6_n107), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_6_n101), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_6_n86), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_6_n87), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n9), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_6_n88), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_6_n89), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_6_n90), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_6_n91), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_6_n92), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_6_n93), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_6_n94), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_6_n95), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_6_n96), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_6_n97), 
        .CK(npu_inst_pe_1_1_6_net4162), .RN(npu_inst_pe_1_1_6_n10), .Q(
        npu_inst_pe_1_1_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_6_net4156) );
  CLKGATETST_X1 npu_inst_pe_1_1_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n47), .SE(1'b0), .GCK(npu_inst_pe_1_1_6_net4162) );
  MUX2_X1 npu_inst_pe_1_1_7_U153 ( .A(npu_inst_pe_1_1_7_n31), .B(
        npu_inst_pe_1_1_7_n28), .S(npu_inst_pe_1_1_7_n7), .Z(
        npu_inst_pe_1_1_7_N93) );
  MUX2_X1 npu_inst_pe_1_1_7_U152 ( .A(npu_inst_pe_1_1_7_n30), .B(
        npu_inst_pe_1_1_7_n29), .S(npu_inst_pe_1_1_7_n5), .Z(
        npu_inst_pe_1_1_7_n31) );
  MUX2_X1 npu_inst_pe_1_1_7_U151 ( .A(npu_inst_pe_1_1_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_1_7_n3), .Z(
        npu_inst_pe_1_1_7_n30) );
  MUX2_X1 npu_inst_pe_1_1_7_U150 ( .A(npu_inst_pe_1_1_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_1_7_n3), .Z(
        npu_inst_pe_1_1_7_n29) );
  MUX2_X1 npu_inst_pe_1_1_7_U149 ( .A(npu_inst_pe_1_1_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_1_7_n3), .Z(
        npu_inst_pe_1_1_7_n28) );
  MUX2_X1 npu_inst_pe_1_1_7_U148 ( .A(npu_inst_pe_1_1_7_n25), .B(
        npu_inst_pe_1_1_7_n22), .S(npu_inst_pe_1_1_7_n7), .Z(
        npu_inst_pe_1_1_7_N94) );
  MUX2_X1 npu_inst_pe_1_1_7_U147 ( .A(npu_inst_pe_1_1_7_n24), .B(
        npu_inst_pe_1_1_7_n23), .S(npu_inst_pe_1_1_7_n5), .Z(
        npu_inst_pe_1_1_7_n25) );
  MUX2_X1 npu_inst_pe_1_1_7_U146 ( .A(npu_inst_pe_1_1_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_1_7_n3), .Z(
        npu_inst_pe_1_1_7_n24) );
  MUX2_X1 npu_inst_pe_1_1_7_U145 ( .A(npu_inst_pe_1_1_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_1_7_n3), .Z(
        npu_inst_pe_1_1_7_n23) );
  MUX2_X1 npu_inst_pe_1_1_7_U144 ( .A(npu_inst_pe_1_1_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_1_7_n3), .Z(
        npu_inst_pe_1_1_7_n22) );
  MUX2_X1 npu_inst_pe_1_1_7_U143 ( .A(npu_inst_pe_1_1_7_n21), .B(
        npu_inst_pe_1_1_7_n18), .S(npu_inst_pe_1_1_7_n7), .Z(
        npu_inst_int_data_x_1__7__1_) );
  MUX2_X1 npu_inst_pe_1_1_7_U142 ( .A(npu_inst_pe_1_1_7_n20), .B(
        npu_inst_pe_1_1_7_n19), .S(npu_inst_pe_1_1_7_n5), .Z(
        npu_inst_pe_1_1_7_n21) );
  MUX2_X1 npu_inst_pe_1_1_7_U141 ( .A(npu_inst_pe_1_1_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_1_7_n3), .Z(
        npu_inst_pe_1_1_7_n20) );
  MUX2_X1 npu_inst_pe_1_1_7_U140 ( .A(npu_inst_pe_1_1_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_1_7_n3), .Z(
        npu_inst_pe_1_1_7_n19) );
  MUX2_X1 npu_inst_pe_1_1_7_U139 ( .A(npu_inst_pe_1_1_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_1_7_n3), .Z(
        npu_inst_pe_1_1_7_n18) );
  MUX2_X1 npu_inst_pe_1_1_7_U138 ( .A(npu_inst_pe_1_1_7_n17), .B(
        npu_inst_pe_1_1_7_n14), .S(npu_inst_pe_1_1_7_n7), .Z(
        npu_inst_int_data_x_1__7__0_) );
  MUX2_X1 npu_inst_pe_1_1_7_U137 ( .A(npu_inst_pe_1_1_7_n16), .B(
        npu_inst_pe_1_1_7_n15), .S(npu_inst_pe_1_1_7_n5), .Z(
        npu_inst_pe_1_1_7_n17) );
  MUX2_X1 npu_inst_pe_1_1_7_U136 ( .A(npu_inst_pe_1_1_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_1_7_n3), .Z(
        npu_inst_pe_1_1_7_n16) );
  MUX2_X1 npu_inst_pe_1_1_7_U135 ( .A(npu_inst_pe_1_1_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_1_7_n3), .Z(
        npu_inst_pe_1_1_7_n15) );
  MUX2_X1 npu_inst_pe_1_1_7_U134 ( .A(npu_inst_pe_1_1_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_1_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_1_7_n3), .Z(
        npu_inst_pe_1_1_7_n14) );
  XOR2_X1 npu_inst_pe_1_1_7_U133 ( .A(npu_inst_pe_1_1_7_int_data_0_), .B(
        npu_inst_int_data_res_1__7__0_), .Z(npu_inst_pe_1_1_7_N73) );
  AND2_X1 npu_inst_pe_1_1_7_U132 ( .A1(npu_inst_int_data_res_1__7__0_), .A2(
        npu_inst_pe_1_1_7_int_data_0_), .ZN(npu_inst_pe_1_1_7_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_1_7_U131 ( .A(npu_inst_int_data_res_1__7__0_), .B(
        npu_inst_pe_1_1_7_n12), .ZN(npu_inst_pe_1_1_7_N65) );
  OR2_X1 npu_inst_pe_1_1_7_U130 ( .A1(npu_inst_pe_1_1_7_n12), .A2(
        npu_inst_int_data_res_1__7__0_), .ZN(npu_inst_pe_1_1_7_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_1_7_U129 ( .A(npu_inst_int_data_res_1__7__2_), .B(
        npu_inst_pe_1_1_7_add_79_carry_2_), .Z(npu_inst_pe_1_1_7_N75) );
  AND2_X1 npu_inst_pe_1_1_7_U128 ( .A1(npu_inst_pe_1_1_7_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_1__7__2_), .ZN(
        npu_inst_pe_1_1_7_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_1_7_U127 ( .A(npu_inst_int_data_res_1__7__3_), .B(
        npu_inst_pe_1_1_7_add_79_carry_3_), .Z(npu_inst_pe_1_1_7_N76) );
  AND2_X1 npu_inst_pe_1_1_7_U126 ( .A1(npu_inst_pe_1_1_7_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_1__7__3_), .ZN(
        npu_inst_pe_1_1_7_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_1_7_U125 ( .A(npu_inst_int_data_res_1__7__4_), .B(
        npu_inst_pe_1_1_7_add_79_carry_4_), .Z(npu_inst_pe_1_1_7_N77) );
  AND2_X1 npu_inst_pe_1_1_7_U124 ( .A1(npu_inst_pe_1_1_7_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_1__7__4_), .ZN(
        npu_inst_pe_1_1_7_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_1_7_U123 ( .A(npu_inst_int_data_res_1__7__5_), .B(
        npu_inst_pe_1_1_7_add_79_carry_5_), .Z(npu_inst_pe_1_1_7_N78) );
  AND2_X1 npu_inst_pe_1_1_7_U122 ( .A1(npu_inst_pe_1_1_7_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_1__7__5_), .ZN(
        npu_inst_pe_1_1_7_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_1_7_U121 ( .A(npu_inst_int_data_res_1__7__6_), .B(
        npu_inst_pe_1_1_7_add_79_carry_6_), .Z(npu_inst_pe_1_1_7_N79) );
  AND2_X1 npu_inst_pe_1_1_7_U120 ( .A1(npu_inst_pe_1_1_7_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_1__7__6_), .ZN(
        npu_inst_pe_1_1_7_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_1_7_U119 ( .A(npu_inst_int_data_res_1__7__7_), .B(
        npu_inst_pe_1_1_7_add_79_carry_7_), .Z(npu_inst_pe_1_1_7_N80) );
  XNOR2_X1 npu_inst_pe_1_1_7_U118 ( .A(npu_inst_pe_1_1_7_sub_77_carry_2_), .B(
        npu_inst_int_data_res_1__7__2_), .ZN(npu_inst_pe_1_1_7_N67) );
  OR2_X1 npu_inst_pe_1_1_7_U117 ( .A1(npu_inst_int_data_res_1__7__2_), .A2(
        npu_inst_pe_1_1_7_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_1_7_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_1_7_U116 ( .A(npu_inst_pe_1_1_7_sub_77_carry_3_), .B(
        npu_inst_int_data_res_1__7__3_), .ZN(npu_inst_pe_1_1_7_N68) );
  OR2_X1 npu_inst_pe_1_1_7_U115 ( .A1(npu_inst_int_data_res_1__7__3_), .A2(
        npu_inst_pe_1_1_7_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_1_7_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_1_7_U114 ( .A(npu_inst_pe_1_1_7_sub_77_carry_4_), .B(
        npu_inst_int_data_res_1__7__4_), .ZN(npu_inst_pe_1_1_7_N69) );
  OR2_X1 npu_inst_pe_1_1_7_U113 ( .A1(npu_inst_int_data_res_1__7__4_), .A2(
        npu_inst_pe_1_1_7_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_1_7_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_1_7_U112 ( .A(npu_inst_pe_1_1_7_sub_77_carry_5_), .B(
        npu_inst_int_data_res_1__7__5_), .ZN(npu_inst_pe_1_1_7_N70) );
  OR2_X1 npu_inst_pe_1_1_7_U111 ( .A1(npu_inst_int_data_res_1__7__5_), .A2(
        npu_inst_pe_1_1_7_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_1_7_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_1_7_U110 ( .A(npu_inst_pe_1_1_7_sub_77_carry_6_), .B(
        npu_inst_int_data_res_1__7__6_), .ZN(npu_inst_pe_1_1_7_N71) );
  OR2_X1 npu_inst_pe_1_1_7_U109 ( .A1(npu_inst_int_data_res_1__7__6_), .A2(
        npu_inst_pe_1_1_7_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_1_7_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_1_7_U108 ( .A(npu_inst_int_data_res_1__7__7_), .B(
        npu_inst_pe_1_1_7_sub_77_carry_7_), .ZN(npu_inst_pe_1_1_7_N72) );
  INV_X1 npu_inst_pe_1_1_7_U107 ( .A(npu_inst_n61), .ZN(npu_inst_pe_1_1_7_n6)
         );
  INV_X1 npu_inst_pe_1_1_7_U106 ( .A(npu_inst_pe_1_1_7_n6), .ZN(
        npu_inst_pe_1_1_7_n5) );
  INV_X1 npu_inst_pe_1_1_7_U105 ( .A(npu_inst_n40), .ZN(npu_inst_pe_1_1_7_n2)
         );
  AOI22_X1 npu_inst_pe_1_1_7_U104 ( .A1(npu_inst_int_data_y_2__7__0_), .A2(
        npu_inst_pe_1_1_7_n58), .B1(npu_inst_pe_1_1_7_n118), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_1_7_n57) );
  INV_X1 npu_inst_pe_1_1_7_U103 ( .A(npu_inst_pe_1_1_7_n57), .ZN(
        npu_inst_pe_1_1_7_n107) );
  AOI22_X1 npu_inst_pe_1_1_7_U102 ( .A1(npu_inst_int_data_y_2__7__0_), .A2(
        npu_inst_pe_1_1_7_n54), .B1(npu_inst_pe_1_1_7_n117), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_1_7_n53) );
  INV_X1 npu_inst_pe_1_1_7_U99 ( .A(npu_inst_pe_1_1_7_n53), .ZN(
        npu_inst_pe_1_1_7_n108) );
  AOI22_X1 npu_inst_pe_1_1_7_U98 ( .A1(npu_inst_int_data_y_2__7__0_), .A2(
        npu_inst_pe_1_1_7_n50), .B1(npu_inst_pe_1_1_7_n116), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_1_7_n49) );
  INV_X1 npu_inst_pe_1_1_7_U97 ( .A(npu_inst_pe_1_1_7_n49), .ZN(
        npu_inst_pe_1_1_7_n109) );
  AOI22_X1 npu_inst_pe_1_1_7_U96 ( .A1(npu_inst_int_data_y_2__7__0_), .A2(
        npu_inst_pe_1_1_7_n46), .B1(npu_inst_pe_1_1_7_n115), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_1_7_n45) );
  INV_X1 npu_inst_pe_1_1_7_U95 ( .A(npu_inst_pe_1_1_7_n45), .ZN(
        npu_inst_pe_1_1_7_n110) );
  AOI22_X1 npu_inst_pe_1_1_7_U94 ( .A1(npu_inst_int_data_y_2__7__0_), .A2(
        npu_inst_pe_1_1_7_n42), .B1(npu_inst_pe_1_1_7_n114), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_1_7_n41) );
  INV_X1 npu_inst_pe_1_1_7_U93 ( .A(npu_inst_pe_1_1_7_n41), .ZN(
        npu_inst_pe_1_1_7_n111) );
  AOI22_X1 npu_inst_pe_1_1_7_U92 ( .A1(npu_inst_int_data_y_2__7__1_), .A2(
        npu_inst_pe_1_1_7_n58), .B1(npu_inst_pe_1_1_7_n118), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_1_7_n59) );
  INV_X1 npu_inst_pe_1_1_7_U91 ( .A(npu_inst_pe_1_1_7_n59), .ZN(
        npu_inst_pe_1_1_7_n101) );
  AOI22_X1 npu_inst_pe_1_1_7_U90 ( .A1(npu_inst_int_data_y_2__7__1_), .A2(
        npu_inst_pe_1_1_7_n54), .B1(npu_inst_pe_1_1_7_n117), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_1_7_n55) );
  INV_X1 npu_inst_pe_1_1_7_U89 ( .A(npu_inst_pe_1_1_7_n55), .ZN(
        npu_inst_pe_1_1_7_n102) );
  AOI22_X1 npu_inst_pe_1_1_7_U88 ( .A1(npu_inst_int_data_y_2__7__1_), .A2(
        npu_inst_pe_1_1_7_n50), .B1(npu_inst_pe_1_1_7_n116), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_1_7_n51) );
  INV_X1 npu_inst_pe_1_1_7_U87 ( .A(npu_inst_pe_1_1_7_n51), .ZN(
        npu_inst_pe_1_1_7_n103) );
  AOI22_X1 npu_inst_pe_1_1_7_U86 ( .A1(npu_inst_int_data_y_2__7__1_), .A2(
        npu_inst_pe_1_1_7_n46), .B1(npu_inst_pe_1_1_7_n115), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_1_7_n47) );
  INV_X1 npu_inst_pe_1_1_7_U85 ( .A(npu_inst_pe_1_1_7_n47), .ZN(
        npu_inst_pe_1_1_7_n104) );
  AOI22_X1 npu_inst_pe_1_1_7_U84 ( .A1(npu_inst_int_data_y_2__7__1_), .A2(
        npu_inst_pe_1_1_7_n42), .B1(npu_inst_pe_1_1_7_n114), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_1_7_n43) );
  INV_X1 npu_inst_pe_1_1_7_U83 ( .A(npu_inst_pe_1_1_7_n43), .ZN(
        npu_inst_pe_1_1_7_n105) );
  AOI22_X1 npu_inst_pe_1_1_7_U82 ( .A1(npu_inst_pe_1_1_7_n38), .A2(
        npu_inst_int_data_y_2__7__1_), .B1(npu_inst_pe_1_1_7_n113), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_1_7_n39) );
  INV_X1 npu_inst_pe_1_1_7_U81 ( .A(npu_inst_pe_1_1_7_n39), .ZN(
        npu_inst_pe_1_1_7_n106) );
  AND2_X1 npu_inst_pe_1_1_7_U80 ( .A1(npu_inst_pe_1_1_7_N93), .A2(npu_inst_n40), .ZN(npu_inst_int_data_y_1__7__0_) );
  AOI22_X1 npu_inst_pe_1_1_7_U79 ( .A1(npu_inst_pe_1_1_7_n38), .A2(
        npu_inst_int_data_y_2__7__0_), .B1(npu_inst_pe_1_1_7_n113), .B2(
        npu_inst_pe_1_1_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_1_7_n37) );
  INV_X1 npu_inst_pe_1_1_7_U78 ( .A(npu_inst_pe_1_1_7_n37), .ZN(
        npu_inst_pe_1_1_7_n112) );
  AND2_X1 npu_inst_pe_1_1_7_U77 ( .A1(npu_inst_n40), .A2(npu_inst_pe_1_1_7_N94), .ZN(npu_inst_int_data_y_1__7__1_) );
  AOI222_X1 npu_inst_pe_1_1_7_U76 ( .A1(npu_inst_int_data_res_2__7__0_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N73), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N65), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n84) );
  INV_X1 npu_inst_pe_1_1_7_U75 ( .A(npu_inst_pe_1_1_7_n84), .ZN(
        npu_inst_pe_1_1_7_n100) );
  AOI222_X1 npu_inst_pe_1_1_7_U74 ( .A1(npu_inst_pe_1_1_7_n1), .A2(
        npu_inst_int_data_res_2__7__7_), .B1(npu_inst_pe_1_1_7_N80), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N72), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n75) );
  INV_X1 npu_inst_pe_1_1_7_U73 ( .A(npu_inst_pe_1_1_7_n75), .ZN(
        npu_inst_pe_1_1_7_n32) );
  AOI222_X1 npu_inst_pe_1_1_7_U72 ( .A1(npu_inst_int_data_res_2__7__1_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N74), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N66), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n83) );
  INV_X1 npu_inst_pe_1_1_7_U71 ( .A(npu_inst_pe_1_1_7_n83), .ZN(
        npu_inst_pe_1_1_7_n99) );
  AOI222_X1 npu_inst_pe_1_1_7_U70 ( .A1(npu_inst_int_data_res_2__7__3_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N76), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N68), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n81) );
  INV_X1 npu_inst_pe_1_1_7_U69 ( .A(npu_inst_pe_1_1_7_n81), .ZN(
        npu_inst_pe_1_1_7_n36) );
  AOI222_X1 npu_inst_pe_1_1_7_U68 ( .A1(npu_inst_int_data_res_2__7__4_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N77), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N69), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n80) );
  INV_X1 npu_inst_pe_1_1_7_U67 ( .A(npu_inst_pe_1_1_7_n80), .ZN(
        npu_inst_pe_1_1_7_n35) );
  AOI222_X1 npu_inst_pe_1_1_7_U66 ( .A1(npu_inst_int_data_res_2__7__5_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N78), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N70), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n79) );
  INV_X1 npu_inst_pe_1_1_7_U65 ( .A(npu_inst_pe_1_1_7_n79), .ZN(
        npu_inst_pe_1_1_7_n34) );
  AOI222_X1 npu_inst_pe_1_1_7_U64 ( .A1(npu_inst_int_data_res_2__7__6_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N79), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N71), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n78) );
  INV_X1 npu_inst_pe_1_1_7_U63 ( .A(npu_inst_pe_1_1_7_n78), .ZN(
        npu_inst_pe_1_1_7_n33) );
  AND2_X1 npu_inst_pe_1_1_7_U62 ( .A1(npu_inst_int_data_x_1__7__1_), .A2(
        npu_inst_pe_1_1_7_int_q_weight_1_), .ZN(npu_inst_pe_1_1_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_1_7_U61 ( .A1(npu_inst_int_data_x_1__7__0_), .A2(
        npu_inst_pe_1_1_7_int_q_weight_1_), .ZN(npu_inst_pe_1_1_7_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_1_7_U60 ( .A(npu_inst_pe_1_1_7_int_data_1_), .ZN(
        npu_inst_pe_1_1_7_n13) );
  NAND2_X1 npu_inst_pe_1_1_7_U59 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_1_7_n60), .ZN(npu_inst_pe_1_1_7_n74) );
  OAI21_X1 npu_inst_pe_1_1_7_U58 ( .B1(npu_inst_pe_1_1_7_n63), .B2(
        npu_inst_pe_1_1_7_n60), .A(npu_inst_pe_1_1_7_n74), .ZN(
        npu_inst_pe_1_1_7_n97) );
  NAND2_X1 npu_inst_pe_1_1_7_U57 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_1_7_n60), .ZN(npu_inst_pe_1_1_7_n73) );
  OAI21_X1 npu_inst_pe_1_1_7_U56 ( .B1(npu_inst_pe_1_1_7_n61), .B2(
        npu_inst_pe_1_1_7_n60), .A(npu_inst_pe_1_1_7_n73), .ZN(
        npu_inst_pe_1_1_7_n96) );
  NAND2_X1 npu_inst_pe_1_1_7_U55 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_1_7_n56), .ZN(npu_inst_pe_1_1_7_n72) );
  OAI21_X1 npu_inst_pe_1_1_7_U54 ( .B1(npu_inst_pe_1_1_7_n63), .B2(
        npu_inst_pe_1_1_7_n56), .A(npu_inst_pe_1_1_7_n72), .ZN(
        npu_inst_pe_1_1_7_n95) );
  NAND2_X1 npu_inst_pe_1_1_7_U53 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_1_7_n56), .ZN(npu_inst_pe_1_1_7_n71) );
  OAI21_X1 npu_inst_pe_1_1_7_U52 ( .B1(npu_inst_pe_1_1_7_n61), .B2(
        npu_inst_pe_1_1_7_n56), .A(npu_inst_pe_1_1_7_n71), .ZN(
        npu_inst_pe_1_1_7_n94) );
  NAND2_X1 npu_inst_pe_1_1_7_U51 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_1_7_n52), .ZN(npu_inst_pe_1_1_7_n70) );
  OAI21_X1 npu_inst_pe_1_1_7_U50 ( .B1(npu_inst_pe_1_1_7_n63), .B2(
        npu_inst_pe_1_1_7_n52), .A(npu_inst_pe_1_1_7_n70), .ZN(
        npu_inst_pe_1_1_7_n93) );
  NAND2_X1 npu_inst_pe_1_1_7_U49 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_1_7_n52), .ZN(npu_inst_pe_1_1_7_n69) );
  OAI21_X1 npu_inst_pe_1_1_7_U48 ( .B1(npu_inst_pe_1_1_7_n61), .B2(
        npu_inst_pe_1_1_7_n52), .A(npu_inst_pe_1_1_7_n69), .ZN(
        npu_inst_pe_1_1_7_n92) );
  NAND2_X1 npu_inst_pe_1_1_7_U47 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_1_7_n48), .ZN(npu_inst_pe_1_1_7_n68) );
  OAI21_X1 npu_inst_pe_1_1_7_U46 ( .B1(npu_inst_pe_1_1_7_n63), .B2(
        npu_inst_pe_1_1_7_n48), .A(npu_inst_pe_1_1_7_n68), .ZN(
        npu_inst_pe_1_1_7_n91) );
  NAND2_X1 npu_inst_pe_1_1_7_U45 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_1_7_n48), .ZN(npu_inst_pe_1_1_7_n67) );
  OAI21_X1 npu_inst_pe_1_1_7_U44 ( .B1(npu_inst_pe_1_1_7_n61), .B2(
        npu_inst_pe_1_1_7_n48), .A(npu_inst_pe_1_1_7_n67), .ZN(
        npu_inst_pe_1_1_7_n90) );
  NAND2_X1 npu_inst_pe_1_1_7_U43 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_1_7_n44), .ZN(npu_inst_pe_1_1_7_n66) );
  OAI21_X1 npu_inst_pe_1_1_7_U42 ( .B1(npu_inst_pe_1_1_7_n63), .B2(
        npu_inst_pe_1_1_7_n44), .A(npu_inst_pe_1_1_7_n66), .ZN(
        npu_inst_pe_1_1_7_n89) );
  NAND2_X1 npu_inst_pe_1_1_7_U41 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_1_7_n44), .ZN(npu_inst_pe_1_1_7_n65) );
  OAI21_X1 npu_inst_pe_1_1_7_U40 ( .B1(npu_inst_pe_1_1_7_n61), .B2(
        npu_inst_pe_1_1_7_n44), .A(npu_inst_pe_1_1_7_n65), .ZN(
        npu_inst_pe_1_1_7_n88) );
  NAND2_X1 npu_inst_pe_1_1_7_U39 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_1_7_n40), .ZN(npu_inst_pe_1_1_7_n64) );
  OAI21_X1 npu_inst_pe_1_1_7_U38 ( .B1(npu_inst_pe_1_1_7_n63), .B2(
        npu_inst_pe_1_1_7_n40), .A(npu_inst_pe_1_1_7_n64), .ZN(
        npu_inst_pe_1_1_7_n87) );
  NAND2_X1 npu_inst_pe_1_1_7_U37 ( .A1(npu_inst_pe_1_1_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_1_7_n40), .ZN(npu_inst_pe_1_1_7_n62) );
  OAI21_X1 npu_inst_pe_1_1_7_U36 ( .B1(npu_inst_pe_1_1_7_n61), .B2(
        npu_inst_pe_1_1_7_n40), .A(npu_inst_pe_1_1_7_n62), .ZN(
        npu_inst_pe_1_1_7_n86) );
  NOR3_X1 npu_inst_pe_1_1_7_U35 ( .A1(npu_inst_pe_1_1_7_n26), .A2(npu_inst_n40), .A3(npu_inst_int_ckg[48]), .ZN(npu_inst_pe_1_1_7_n85) );
  OR2_X1 npu_inst_pe_1_1_7_U34 ( .A1(npu_inst_pe_1_1_7_n85), .A2(
        npu_inst_pe_1_1_7_n1), .ZN(npu_inst_pe_1_1_7_N84) );
  AOI222_X1 npu_inst_pe_1_1_7_U33 ( .A1(npu_inst_int_data_res_2__7__2_), .A2(
        npu_inst_pe_1_1_7_n1), .B1(npu_inst_pe_1_1_7_N75), .B2(
        npu_inst_pe_1_1_7_n76), .C1(npu_inst_pe_1_1_7_N67), .C2(
        npu_inst_pe_1_1_7_n77), .ZN(npu_inst_pe_1_1_7_n82) );
  INV_X1 npu_inst_pe_1_1_7_U32 ( .A(npu_inst_pe_1_1_7_n82), .ZN(
        npu_inst_pe_1_1_7_n98) );
  INV_X1 npu_inst_pe_1_1_7_U31 ( .A(npu_inst_pe_1_1_7_int_data_0_), .ZN(
        npu_inst_pe_1_1_7_n12) );
  INV_X1 npu_inst_pe_1_1_7_U30 ( .A(npu_inst_n53), .ZN(npu_inst_pe_1_1_7_n4)
         );
  AOI22_X1 npu_inst_pe_1_1_7_U29 ( .A1(npu_inst_n40), .A2(
        npu_inst_int_data_y_2__7__1_), .B1(npu_inst_pe_1_1_7_n2), .B2(
        int_i_data_h_npu[13]), .ZN(npu_inst_pe_1_1_7_n63) );
  AOI22_X1 npu_inst_pe_1_1_7_U28 ( .A1(npu_inst_n40), .A2(
        npu_inst_int_data_y_2__7__0_), .B1(npu_inst_pe_1_1_7_n2), .B2(
        int_i_data_h_npu[12]), .ZN(npu_inst_pe_1_1_7_n61) );
  OR3_X1 npu_inst_pe_1_1_7_U27 ( .A1(npu_inst_pe_1_1_7_n5), .A2(
        npu_inst_pe_1_1_7_n7), .A3(npu_inst_pe_1_1_7_n4), .ZN(
        npu_inst_pe_1_1_7_n56) );
  OR3_X1 npu_inst_pe_1_1_7_U26 ( .A1(npu_inst_pe_1_1_7_n4), .A2(
        npu_inst_pe_1_1_7_n7), .A3(npu_inst_pe_1_1_7_n6), .ZN(
        npu_inst_pe_1_1_7_n48) );
  INV_X1 npu_inst_pe_1_1_7_U25 ( .A(npu_inst_pe_1_1_7_n4), .ZN(
        npu_inst_pe_1_1_7_n3) );
  OR3_X1 npu_inst_pe_1_1_7_U24 ( .A1(npu_inst_pe_1_1_7_n3), .A2(
        npu_inst_pe_1_1_7_n7), .A3(npu_inst_pe_1_1_7_n6), .ZN(
        npu_inst_pe_1_1_7_n52) );
  OR3_X1 npu_inst_pe_1_1_7_U23 ( .A1(npu_inst_pe_1_1_7_n5), .A2(
        npu_inst_pe_1_1_7_n7), .A3(npu_inst_pe_1_1_7_n3), .ZN(
        npu_inst_pe_1_1_7_n60) );
  BUF_X1 npu_inst_pe_1_1_7_U22 ( .A(npu_inst_n27), .Z(npu_inst_pe_1_1_7_n1) );
  NOR2_X1 npu_inst_pe_1_1_7_U21 ( .A1(npu_inst_pe_1_1_7_n60), .A2(
        npu_inst_pe_1_1_7_n2), .ZN(npu_inst_pe_1_1_7_n58) );
  NOR2_X1 npu_inst_pe_1_1_7_U20 ( .A1(npu_inst_pe_1_1_7_n56), .A2(
        npu_inst_pe_1_1_7_n2), .ZN(npu_inst_pe_1_1_7_n54) );
  NOR2_X1 npu_inst_pe_1_1_7_U19 ( .A1(npu_inst_pe_1_1_7_n52), .A2(
        npu_inst_pe_1_1_7_n2), .ZN(npu_inst_pe_1_1_7_n50) );
  NOR2_X1 npu_inst_pe_1_1_7_U18 ( .A1(npu_inst_pe_1_1_7_n48), .A2(
        npu_inst_pe_1_1_7_n2), .ZN(npu_inst_pe_1_1_7_n46) );
  NOR2_X1 npu_inst_pe_1_1_7_U17 ( .A1(npu_inst_pe_1_1_7_n40), .A2(
        npu_inst_pe_1_1_7_n2), .ZN(npu_inst_pe_1_1_7_n38) );
  NOR2_X1 npu_inst_pe_1_1_7_U16 ( .A1(npu_inst_pe_1_1_7_n44), .A2(
        npu_inst_pe_1_1_7_n2), .ZN(npu_inst_pe_1_1_7_n42) );
  BUF_X1 npu_inst_pe_1_1_7_U15 ( .A(npu_inst_n86), .Z(npu_inst_pe_1_1_7_n7) );
  INV_X1 npu_inst_pe_1_1_7_U14 ( .A(npu_inst_n108), .ZN(npu_inst_pe_1_1_7_n11)
         );
  INV_X1 npu_inst_pe_1_1_7_U13 ( .A(npu_inst_pe_1_1_7_n38), .ZN(
        npu_inst_pe_1_1_7_n113) );
  INV_X1 npu_inst_pe_1_1_7_U12 ( .A(npu_inst_pe_1_1_7_n58), .ZN(
        npu_inst_pe_1_1_7_n118) );
  INV_X1 npu_inst_pe_1_1_7_U11 ( .A(npu_inst_pe_1_1_7_n54), .ZN(
        npu_inst_pe_1_1_7_n117) );
  INV_X1 npu_inst_pe_1_1_7_U10 ( .A(npu_inst_pe_1_1_7_n50), .ZN(
        npu_inst_pe_1_1_7_n116) );
  INV_X1 npu_inst_pe_1_1_7_U9 ( .A(npu_inst_pe_1_1_7_n46), .ZN(
        npu_inst_pe_1_1_7_n115) );
  INV_X1 npu_inst_pe_1_1_7_U8 ( .A(npu_inst_pe_1_1_7_n42), .ZN(
        npu_inst_pe_1_1_7_n114) );
  BUF_X1 npu_inst_pe_1_1_7_U7 ( .A(npu_inst_pe_1_1_7_n11), .Z(
        npu_inst_pe_1_1_7_n10) );
  BUF_X1 npu_inst_pe_1_1_7_U6 ( .A(npu_inst_pe_1_1_7_n11), .Z(
        npu_inst_pe_1_1_7_n9) );
  BUF_X1 npu_inst_pe_1_1_7_U5 ( .A(npu_inst_pe_1_1_7_n11), .Z(
        npu_inst_pe_1_1_7_n8) );
  NOR2_X1 npu_inst_pe_1_1_7_U4 ( .A1(npu_inst_pe_1_1_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_1_7_n1), .ZN(npu_inst_pe_1_1_7_n76) );
  NOR2_X1 npu_inst_pe_1_1_7_U3 ( .A1(npu_inst_pe_1_1_7_n27), .A2(
        npu_inst_pe_1_1_7_n1), .ZN(npu_inst_pe_1_1_7_n77) );
  FA_X1 npu_inst_pe_1_1_7_sub_77_U2_1 ( .A(npu_inst_int_data_res_1__7__1_), 
        .B(npu_inst_pe_1_1_7_n13), .CI(npu_inst_pe_1_1_7_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_1_7_sub_77_carry_2_), .S(npu_inst_pe_1_1_7_N66) );
  FA_X1 npu_inst_pe_1_1_7_add_79_U1_1 ( .A(npu_inst_int_data_res_1__7__1_), 
        .B(npu_inst_pe_1_1_7_int_data_1_), .CI(
        npu_inst_pe_1_1_7_add_79_carry_1_), .CO(
        npu_inst_pe_1_1_7_add_79_carry_2_), .S(npu_inst_pe_1_1_7_N74) );
  NAND3_X1 npu_inst_pe_1_1_7_U101 ( .A1(npu_inst_pe_1_1_7_n4), .A2(
        npu_inst_pe_1_1_7_n6), .A3(npu_inst_pe_1_1_7_n7), .ZN(
        npu_inst_pe_1_1_7_n44) );
  NAND3_X1 npu_inst_pe_1_1_7_U100 ( .A1(npu_inst_pe_1_1_7_n3), .A2(
        npu_inst_pe_1_1_7_n6), .A3(npu_inst_pe_1_1_7_n7), .ZN(
        npu_inst_pe_1_1_7_n40) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_1_7_n33), .CK(
        npu_inst_pe_1_1_7_net4133), .RN(npu_inst_pe_1_1_7_n8), .Q(
        npu_inst_int_data_res_1__7__6_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_1_7_n34), .CK(
        npu_inst_pe_1_1_7_net4133), .RN(npu_inst_pe_1_1_7_n8), .Q(
        npu_inst_int_data_res_1__7__5_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_1_7_n35), .CK(
        npu_inst_pe_1_1_7_net4133), .RN(npu_inst_pe_1_1_7_n8), .Q(
        npu_inst_int_data_res_1__7__4_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_1_7_n36), .CK(
        npu_inst_pe_1_1_7_net4133), .RN(npu_inst_pe_1_1_7_n8), .Q(
        npu_inst_int_data_res_1__7__3_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_1_7_n98), .CK(
        npu_inst_pe_1_1_7_net4133), .RN(npu_inst_pe_1_1_7_n8), .Q(
        npu_inst_int_data_res_1__7__2_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_1_7_n99), .CK(
        npu_inst_pe_1_1_7_net4133), .RN(npu_inst_pe_1_1_7_n8), .Q(
        npu_inst_int_data_res_1__7__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_1_7_n32), .CK(
        npu_inst_pe_1_1_7_net4133), .RN(npu_inst_pe_1_1_7_n8), .Q(
        npu_inst_int_data_res_1__7__7_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_1_7_n100), 
        .CK(npu_inst_pe_1_1_7_net4133), .RN(npu_inst_pe_1_1_7_n8), .Q(
        npu_inst_int_data_res_1__7__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_weight_reg_0_ ( .D(npu_inst_n94), .CK(
        npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n8), .Q(
        npu_inst_pe_1_1_7_int_q_weight_0_), .QN(npu_inst_pe_1_1_7_n27) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_weight_reg_1_ ( .D(npu_inst_n100), .CK(
        npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n8), .Q(
        npu_inst_pe_1_1_7_int_q_weight_1_), .QN(npu_inst_pe_1_1_7_n26) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_1_7_n112), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n8), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_1_7_n106), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n8), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_1_7_n111), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_1_7_n105), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_1_7_n110), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_1_7_n104), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_1_7_n109), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_1_7_n103), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_1_7_n108), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_1_7_n102), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_1_7_n107), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_1_7_n101), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_1_7_n86), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_1_7_n87), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n9), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_1_7_n88), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_1_7_n89), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_1_7_n90), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_1_7_n91), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_1_7_n92), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_1_7_n93), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_1_7_n94), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_1_7_n95), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_1_7_n96), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_1_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_1_7_n97), 
        .CK(npu_inst_pe_1_1_7_net4139), .RN(npu_inst_pe_1_1_7_n10), .Q(
        npu_inst_pe_1_1_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_1_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_1_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_1_7_net4133) );
  CLKGATETST_X1 npu_inst_pe_1_1_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n47), .SE(1'b0), .GCK(npu_inst_pe_1_1_7_net4139) );
  MUX2_X1 npu_inst_pe_1_2_0_U152 ( .A(npu_inst_pe_1_2_0_n30), .B(
        npu_inst_pe_1_2_0_n25), .S(npu_inst_pe_1_2_0_n6), .Z(
        npu_inst_pe_1_2_0_N93) );
  MUX2_X1 npu_inst_pe_1_2_0_U151 ( .A(npu_inst_pe_1_2_0_n29), .B(
        npu_inst_pe_1_2_0_n28), .S(npu_inst_n60), .Z(npu_inst_pe_1_2_0_n30) );
  MUX2_X1 npu_inst_pe_1_2_0_U150 ( .A(npu_inst_pe_1_2_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_0_n3), .Z(
        npu_inst_pe_1_2_0_n29) );
  MUX2_X1 npu_inst_pe_1_2_0_U149 ( .A(npu_inst_pe_1_2_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_0_n3), .Z(
        npu_inst_pe_1_2_0_n28) );
  MUX2_X1 npu_inst_pe_1_2_0_U148 ( .A(npu_inst_pe_1_2_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_0_n3), .Z(
        npu_inst_pe_1_2_0_n25) );
  MUX2_X1 npu_inst_pe_1_2_0_U147 ( .A(npu_inst_pe_1_2_0_n24), .B(
        npu_inst_pe_1_2_0_n21), .S(npu_inst_pe_1_2_0_n6), .Z(
        npu_inst_pe_1_2_0_N94) );
  MUX2_X1 npu_inst_pe_1_2_0_U146 ( .A(npu_inst_pe_1_2_0_n23), .B(
        npu_inst_pe_1_2_0_n22), .S(npu_inst_n60), .Z(npu_inst_pe_1_2_0_n24) );
  MUX2_X1 npu_inst_pe_1_2_0_U145 ( .A(npu_inst_pe_1_2_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_0_n3), .Z(
        npu_inst_pe_1_2_0_n23) );
  MUX2_X1 npu_inst_pe_1_2_0_U144 ( .A(npu_inst_pe_1_2_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_0_n3), .Z(
        npu_inst_pe_1_2_0_n22) );
  MUX2_X1 npu_inst_pe_1_2_0_U143 ( .A(npu_inst_pe_1_2_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_0_n3), .Z(
        npu_inst_pe_1_2_0_n21) );
  MUX2_X1 npu_inst_pe_1_2_0_U142 ( .A(npu_inst_pe_1_2_0_n20), .B(
        npu_inst_pe_1_2_0_n17), .S(npu_inst_pe_1_2_0_n6), .Z(
        npu_inst_pe_1_2_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_2_0_U141 ( .A(npu_inst_pe_1_2_0_n19), .B(
        npu_inst_pe_1_2_0_n18), .S(npu_inst_n60), .Z(npu_inst_pe_1_2_0_n20) );
  MUX2_X1 npu_inst_pe_1_2_0_U140 ( .A(npu_inst_pe_1_2_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_0_n3), .Z(
        npu_inst_pe_1_2_0_n19) );
  MUX2_X1 npu_inst_pe_1_2_0_U139 ( .A(npu_inst_pe_1_2_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_0_n3), .Z(
        npu_inst_pe_1_2_0_n18) );
  MUX2_X1 npu_inst_pe_1_2_0_U138 ( .A(npu_inst_pe_1_2_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_0_n3), .Z(
        npu_inst_pe_1_2_0_n17) );
  MUX2_X1 npu_inst_pe_1_2_0_U137 ( .A(npu_inst_pe_1_2_0_n16), .B(
        npu_inst_pe_1_2_0_n13), .S(npu_inst_pe_1_2_0_n6), .Z(
        npu_inst_pe_1_2_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_2_0_U136 ( .A(npu_inst_pe_1_2_0_n15), .B(
        npu_inst_pe_1_2_0_n14), .S(npu_inst_n60), .Z(npu_inst_pe_1_2_0_n16) );
  MUX2_X1 npu_inst_pe_1_2_0_U135 ( .A(npu_inst_pe_1_2_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_0_n3), .Z(
        npu_inst_pe_1_2_0_n15) );
  MUX2_X1 npu_inst_pe_1_2_0_U134 ( .A(npu_inst_pe_1_2_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_0_n3), .Z(
        npu_inst_pe_1_2_0_n14) );
  MUX2_X1 npu_inst_pe_1_2_0_U133 ( .A(npu_inst_pe_1_2_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_0_n3), .Z(
        npu_inst_pe_1_2_0_n13) );
  XOR2_X1 npu_inst_pe_1_2_0_U132 ( .A(npu_inst_pe_1_2_0_int_data_0_), .B(
        npu_inst_int_data_res_2__0__0_), .Z(npu_inst_pe_1_2_0_N73) );
  AND2_X1 npu_inst_pe_1_2_0_U131 ( .A1(npu_inst_int_data_res_2__0__0_), .A2(
        npu_inst_pe_1_2_0_int_data_0_), .ZN(npu_inst_pe_1_2_0_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_0_U130 ( .A(npu_inst_int_data_res_2__0__0_), .B(
        npu_inst_pe_1_2_0_n11), .ZN(npu_inst_pe_1_2_0_N65) );
  OR2_X1 npu_inst_pe_1_2_0_U129 ( .A1(npu_inst_pe_1_2_0_n11), .A2(
        npu_inst_int_data_res_2__0__0_), .ZN(npu_inst_pe_1_2_0_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_0_U128 ( .A(npu_inst_int_data_res_2__0__2_), .B(
        npu_inst_pe_1_2_0_add_79_carry_2_), .Z(npu_inst_pe_1_2_0_N75) );
  AND2_X1 npu_inst_pe_1_2_0_U127 ( .A1(npu_inst_pe_1_2_0_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_2__0__2_), .ZN(
        npu_inst_pe_1_2_0_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_0_U126 ( .A(npu_inst_int_data_res_2__0__3_), .B(
        npu_inst_pe_1_2_0_add_79_carry_3_), .Z(npu_inst_pe_1_2_0_N76) );
  AND2_X1 npu_inst_pe_1_2_0_U125 ( .A1(npu_inst_pe_1_2_0_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_2__0__3_), .ZN(
        npu_inst_pe_1_2_0_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_0_U124 ( .A(npu_inst_int_data_res_2__0__4_), .B(
        npu_inst_pe_1_2_0_add_79_carry_4_), .Z(npu_inst_pe_1_2_0_N77) );
  AND2_X1 npu_inst_pe_1_2_0_U123 ( .A1(npu_inst_pe_1_2_0_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_2__0__4_), .ZN(
        npu_inst_pe_1_2_0_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_0_U122 ( .A(npu_inst_int_data_res_2__0__5_), .B(
        npu_inst_pe_1_2_0_add_79_carry_5_), .Z(npu_inst_pe_1_2_0_N78) );
  AND2_X1 npu_inst_pe_1_2_0_U121 ( .A1(npu_inst_pe_1_2_0_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_2__0__5_), .ZN(
        npu_inst_pe_1_2_0_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_0_U120 ( .A(npu_inst_int_data_res_2__0__6_), .B(
        npu_inst_pe_1_2_0_add_79_carry_6_), .Z(npu_inst_pe_1_2_0_N79) );
  AND2_X1 npu_inst_pe_1_2_0_U119 ( .A1(npu_inst_pe_1_2_0_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_2__0__6_), .ZN(
        npu_inst_pe_1_2_0_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_0_U118 ( .A(npu_inst_int_data_res_2__0__7_), .B(
        npu_inst_pe_1_2_0_add_79_carry_7_), .Z(npu_inst_pe_1_2_0_N80) );
  XNOR2_X1 npu_inst_pe_1_2_0_U117 ( .A(npu_inst_pe_1_2_0_sub_77_carry_2_), .B(
        npu_inst_int_data_res_2__0__2_), .ZN(npu_inst_pe_1_2_0_N67) );
  OR2_X1 npu_inst_pe_1_2_0_U116 ( .A1(npu_inst_int_data_res_2__0__2_), .A2(
        npu_inst_pe_1_2_0_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_2_0_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_0_U115 ( .A(npu_inst_pe_1_2_0_sub_77_carry_3_), .B(
        npu_inst_int_data_res_2__0__3_), .ZN(npu_inst_pe_1_2_0_N68) );
  OR2_X1 npu_inst_pe_1_2_0_U114 ( .A1(npu_inst_int_data_res_2__0__3_), .A2(
        npu_inst_pe_1_2_0_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_2_0_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_0_U113 ( .A(npu_inst_pe_1_2_0_sub_77_carry_4_), .B(
        npu_inst_int_data_res_2__0__4_), .ZN(npu_inst_pe_1_2_0_N69) );
  OR2_X1 npu_inst_pe_1_2_0_U112 ( .A1(npu_inst_int_data_res_2__0__4_), .A2(
        npu_inst_pe_1_2_0_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_2_0_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_0_U111 ( .A(npu_inst_pe_1_2_0_sub_77_carry_5_), .B(
        npu_inst_int_data_res_2__0__5_), .ZN(npu_inst_pe_1_2_0_N70) );
  OR2_X1 npu_inst_pe_1_2_0_U110 ( .A1(npu_inst_int_data_res_2__0__5_), .A2(
        npu_inst_pe_1_2_0_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_2_0_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_0_U109 ( .A(npu_inst_pe_1_2_0_sub_77_carry_6_), .B(
        npu_inst_int_data_res_2__0__6_), .ZN(npu_inst_pe_1_2_0_N71) );
  OR2_X1 npu_inst_pe_1_2_0_U108 ( .A1(npu_inst_int_data_res_2__0__6_), .A2(
        npu_inst_pe_1_2_0_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_2_0_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_0_U107 ( .A(npu_inst_int_data_res_2__0__7_), .B(
        npu_inst_pe_1_2_0_sub_77_carry_7_), .ZN(npu_inst_pe_1_2_0_N72) );
  INV_X1 npu_inst_pe_1_2_0_U106 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_2_0_n5)
         );
  INV_X1 npu_inst_pe_1_2_0_U105 ( .A(npu_inst_n40), .ZN(npu_inst_pe_1_2_0_n2)
         );
  AOI22_X1 npu_inst_pe_1_2_0_U104 ( .A1(npu_inst_int_data_y_3__0__0_), .A2(
        npu_inst_pe_1_2_0_n58), .B1(npu_inst_pe_1_2_0_n117), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_0_n57) );
  INV_X1 npu_inst_pe_1_2_0_U103 ( .A(npu_inst_pe_1_2_0_n57), .ZN(
        npu_inst_pe_1_2_0_n106) );
  AOI22_X1 npu_inst_pe_1_2_0_U102 ( .A1(npu_inst_int_data_y_3__0__0_), .A2(
        npu_inst_pe_1_2_0_n54), .B1(npu_inst_pe_1_2_0_n116), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_0_n53) );
  INV_X1 npu_inst_pe_1_2_0_U99 ( .A(npu_inst_pe_1_2_0_n53), .ZN(
        npu_inst_pe_1_2_0_n107) );
  AOI22_X1 npu_inst_pe_1_2_0_U98 ( .A1(npu_inst_int_data_y_3__0__0_), .A2(
        npu_inst_pe_1_2_0_n50), .B1(npu_inst_pe_1_2_0_n115), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_0_n49) );
  INV_X1 npu_inst_pe_1_2_0_U97 ( .A(npu_inst_pe_1_2_0_n49), .ZN(
        npu_inst_pe_1_2_0_n108) );
  AOI22_X1 npu_inst_pe_1_2_0_U96 ( .A1(npu_inst_int_data_y_3__0__0_), .A2(
        npu_inst_pe_1_2_0_n46), .B1(npu_inst_pe_1_2_0_n114), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_0_n45) );
  INV_X1 npu_inst_pe_1_2_0_U95 ( .A(npu_inst_pe_1_2_0_n45), .ZN(
        npu_inst_pe_1_2_0_n109) );
  AOI22_X1 npu_inst_pe_1_2_0_U94 ( .A1(npu_inst_int_data_y_3__0__0_), .A2(
        npu_inst_pe_1_2_0_n42), .B1(npu_inst_pe_1_2_0_n113), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_0_n41) );
  INV_X1 npu_inst_pe_1_2_0_U93 ( .A(npu_inst_pe_1_2_0_n41), .ZN(
        npu_inst_pe_1_2_0_n110) );
  AOI22_X1 npu_inst_pe_1_2_0_U92 ( .A1(npu_inst_int_data_y_3__0__1_), .A2(
        npu_inst_pe_1_2_0_n58), .B1(npu_inst_pe_1_2_0_n117), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_0_n59) );
  INV_X1 npu_inst_pe_1_2_0_U91 ( .A(npu_inst_pe_1_2_0_n59), .ZN(
        npu_inst_pe_1_2_0_n100) );
  AOI22_X1 npu_inst_pe_1_2_0_U90 ( .A1(npu_inst_int_data_y_3__0__1_), .A2(
        npu_inst_pe_1_2_0_n54), .B1(npu_inst_pe_1_2_0_n116), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_0_n55) );
  INV_X1 npu_inst_pe_1_2_0_U89 ( .A(npu_inst_pe_1_2_0_n55), .ZN(
        npu_inst_pe_1_2_0_n101) );
  AOI22_X1 npu_inst_pe_1_2_0_U88 ( .A1(npu_inst_int_data_y_3__0__1_), .A2(
        npu_inst_pe_1_2_0_n50), .B1(npu_inst_pe_1_2_0_n115), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_0_n51) );
  INV_X1 npu_inst_pe_1_2_0_U87 ( .A(npu_inst_pe_1_2_0_n51), .ZN(
        npu_inst_pe_1_2_0_n102) );
  AOI22_X1 npu_inst_pe_1_2_0_U86 ( .A1(npu_inst_int_data_y_3__0__1_), .A2(
        npu_inst_pe_1_2_0_n46), .B1(npu_inst_pe_1_2_0_n114), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_0_n47) );
  INV_X1 npu_inst_pe_1_2_0_U85 ( .A(npu_inst_pe_1_2_0_n47), .ZN(
        npu_inst_pe_1_2_0_n103) );
  AOI22_X1 npu_inst_pe_1_2_0_U84 ( .A1(npu_inst_int_data_y_3__0__1_), .A2(
        npu_inst_pe_1_2_0_n42), .B1(npu_inst_pe_1_2_0_n113), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_0_n43) );
  INV_X1 npu_inst_pe_1_2_0_U83 ( .A(npu_inst_pe_1_2_0_n43), .ZN(
        npu_inst_pe_1_2_0_n104) );
  AOI22_X1 npu_inst_pe_1_2_0_U82 ( .A1(npu_inst_pe_1_2_0_n38), .A2(
        npu_inst_int_data_y_3__0__1_), .B1(npu_inst_pe_1_2_0_n112), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_0_n39) );
  INV_X1 npu_inst_pe_1_2_0_U81 ( .A(npu_inst_pe_1_2_0_n39), .ZN(
        npu_inst_pe_1_2_0_n105) );
  AND2_X1 npu_inst_pe_1_2_0_U80 ( .A1(npu_inst_pe_1_2_0_N93), .A2(npu_inst_n40), .ZN(npu_inst_int_data_y_2__0__0_) );
  NAND2_X1 npu_inst_pe_1_2_0_U79 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_0_n60), .ZN(npu_inst_pe_1_2_0_n74) );
  OAI21_X1 npu_inst_pe_1_2_0_U78 ( .B1(npu_inst_pe_1_2_0_n63), .B2(
        npu_inst_pe_1_2_0_n60), .A(npu_inst_pe_1_2_0_n74), .ZN(
        npu_inst_pe_1_2_0_n97) );
  NAND2_X1 npu_inst_pe_1_2_0_U77 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_0_n60), .ZN(npu_inst_pe_1_2_0_n73) );
  OAI21_X1 npu_inst_pe_1_2_0_U76 ( .B1(npu_inst_pe_1_2_0_n61), .B2(
        npu_inst_pe_1_2_0_n60), .A(npu_inst_pe_1_2_0_n73), .ZN(
        npu_inst_pe_1_2_0_n96) );
  NAND2_X1 npu_inst_pe_1_2_0_U75 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_0_n56), .ZN(npu_inst_pe_1_2_0_n72) );
  OAI21_X1 npu_inst_pe_1_2_0_U74 ( .B1(npu_inst_pe_1_2_0_n63), .B2(
        npu_inst_pe_1_2_0_n56), .A(npu_inst_pe_1_2_0_n72), .ZN(
        npu_inst_pe_1_2_0_n95) );
  NAND2_X1 npu_inst_pe_1_2_0_U73 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_0_n56), .ZN(npu_inst_pe_1_2_0_n71) );
  OAI21_X1 npu_inst_pe_1_2_0_U72 ( .B1(npu_inst_pe_1_2_0_n61), .B2(
        npu_inst_pe_1_2_0_n56), .A(npu_inst_pe_1_2_0_n71), .ZN(
        npu_inst_pe_1_2_0_n94) );
  NAND2_X1 npu_inst_pe_1_2_0_U71 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_0_n52), .ZN(npu_inst_pe_1_2_0_n70) );
  OAI21_X1 npu_inst_pe_1_2_0_U70 ( .B1(npu_inst_pe_1_2_0_n63), .B2(
        npu_inst_pe_1_2_0_n52), .A(npu_inst_pe_1_2_0_n70), .ZN(
        npu_inst_pe_1_2_0_n93) );
  NAND2_X1 npu_inst_pe_1_2_0_U69 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_0_n52), .ZN(npu_inst_pe_1_2_0_n69) );
  OAI21_X1 npu_inst_pe_1_2_0_U68 ( .B1(npu_inst_pe_1_2_0_n61), .B2(
        npu_inst_pe_1_2_0_n52), .A(npu_inst_pe_1_2_0_n69), .ZN(
        npu_inst_pe_1_2_0_n92) );
  NAND2_X1 npu_inst_pe_1_2_0_U67 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_0_n48), .ZN(npu_inst_pe_1_2_0_n68) );
  OAI21_X1 npu_inst_pe_1_2_0_U66 ( .B1(npu_inst_pe_1_2_0_n63), .B2(
        npu_inst_pe_1_2_0_n48), .A(npu_inst_pe_1_2_0_n68), .ZN(
        npu_inst_pe_1_2_0_n91) );
  NAND2_X1 npu_inst_pe_1_2_0_U65 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_0_n48), .ZN(npu_inst_pe_1_2_0_n67) );
  OAI21_X1 npu_inst_pe_1_2_0_U64 ( .B1(npu_inst_pe_1_2_0_n61), .B2(
        npu_inst_pe_1_2_0_n48), .A(npu_inst_pe_1_2_0_n67), .ZN(
        npu_inst_pe_1_2_0_n90) );
  NAND2_X1 npu_inst_pe_1_2_0_U63 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_0_n44), .ZN(npu_inst_pe_1_2_0_n66) );
  OAI21_X1 npu_inst_pe_1_2_0_U62 ( .B1(npu_inst_pe_1_2_0_n63), .B2(
        npu_inst_pe_1_2_0_n44), .A(npu_inst_pe_1_2_0_n66), .ZN(
        npu_inst_pe_1_2_0_n89) );
  NAND2_X1 npu_inst_pe_1_2_0_U61 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_0_n44), .ZN(npu_inst_pe_1_2_0_n65) );
  OAI21_X1 npu_inst_pe_1_2_0_U60 ( .B1(npu_inst_pe_1_2_0_n61), .B2(
        npu_inst_pe_1_2_0_n44), .A(npu_inst_pe_1_2_0_n65), .ZN(
        npu_inst_pe_1_2_0_n88) );
  NAND2_X1 npu_inst_pe_1_2_0_U59 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_0_n40), .ZN(npu_inst_pe_1_2_0_n64) );
  OAI21_X1 npu_inst_pe_1_2_0_U58 ( .B1(npu_inst_pe_1_2_0_n63), .B2(
        npu_inst_pe_1_2_0_n40), .A(npu_inst_pe_1_2_0_n64), .ZN(
        npu_inst_pe_1_2_0_n87) );
  NAND2_X1 npu_inst_pe_1_2_0_U57 ( .A1(npu_inst_pe_1_2_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_0_n40), .ZN(npu_inst_pe_1_2_0_n62) );
  OAI21_X1 npu_inst_pe_1_2_0_U56 ( .B1(npu_inst_pe_1_2_0_n61), .B2(
        npu_inst_pe_1_2_0_n40), .A(npu_inst_pe_1_2_0_n62), .ZN(
        npu_inst_pe_1_2_0_n86) );
  AOI22_X1 npu_inst_pe_1_2_0_U55 ( .A1(npu_inst_pe_1_2_0_n38), .A2(
        npu_inst_int_data_y_3__0__0_), .B1(npu_inst_pe_1_2_0_n112), .B2(
        npu_inst_pe_1_2_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_0_n37) );
  INV_X1 npu_inst_pe_1_2_0_U54 ( .A(npu_inst_pe_1_2_0_n37), .ZN(
        npu_inst_pe_1_2_0_n111) );
  AND2_X1 npu_inst_pe_1_2_0_U53 ( .A1(npu_inst_n40), .A2(npu_inst_pe_1_2_0_N94), .ZN(npu_inst_int_data_y_2__0__1_) );
  AOI222_X1 npu_inst_pe_1_2_0_U52 ( .A1(npu_inst_int_data_res_3__0__0_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N73), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N65), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n84) );
  INV_X1 npu_inst_pe_1_2_0_U51 ( .A(npu_inst_pe_1_2_0_n84), .ZN(
        npu_inst_pe_1_2_0_n99) );
  AOI222_X1 npu_inst_pe_1_2_0_U50 ( .A1(npu_inst_pe_1_2_0_n1), .A2(
        npu_inst_int_data_res_3__0__7_), .B1(npu_inst_pe_1_2_0_N80), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N72), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n75) );
  INV_X1 npu_inst_pe_1_2_0_U49 ( .A(npu_inst_pe_1_2_0_n75), .ZN(
        npu_inst_pe_1_2_0_n31) );
  AOI222_X1 npu_inst_pe_1_2_0_U48 ( .A1(npu_inst_int_data_res_3__0__1_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N74), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N66), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n83) );
  INV_X1 npu_inst_pe_1_2_0_U47 ( .A(npu_inst_pe_1_2_0_n83), .ZN(
        npu_inst_pe_1_2_0_n98) );
  AOI222_X1 npu_inst_pe_1_2_0_U46 ( .A1(npu_inst_int_data_res_3__0__3_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N76), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N68), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n81) );
  INV_X1 npu_inst_pe_1_2_0_U45 ( .A(npu_inst_pe_1_2_0_n81), .ZN(
        npu_inst_pe_1_2_0_n35) );
  AOI222_X1 npu_inst_pe_1_2_0_U44 ( .A1(npu_inst_int_data_res_3__0__4_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N77), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N69), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n80) );
  INV_X1 npu_inst_pe_1_2_0_U43 ( .A(npu_inst_pe_1_2_0_n80), .ZN(
        npu_inst_pe_1_2_0_n34) );
  AOI222_X1 npu_inst_pe_1_2_0_U42 ( .A1(npu_inst_int_data_res_3__0__5_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N78), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N70), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n79) );
  INV_X1 npu_inst_pe_1_2_0_U41 ( .A(npu_inst_pe_1_2_0_n79), .ZN(
        npu_inst_pe_1_2_0_n33) );
  AOI222_X1 npu_inst_pe_1_2_0_U40 ( .A1(npu_inst_int_data_res_3__0__6_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N79), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N71), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n78) );
  INV_X1 npu_inst_pe_1_2_0_U39 ( .A(npu_inst_pe_1_2_0_n78), .ZN(
        npu_inst_pe_1_2_0_n32) );
  AND2_X1 npu_inst_pe_1_2_0_U38 ( .A1(npu_inst_pe_1_2_0_o_data_h_1_), .A2(
        npu_inst_pe_1_2_0_int_q_weight_1_), .ZN(npu_inst_pe_1_2_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_0_U37 ( .A1(npu_inst_pe_1_2_0_o_data_h_0_), .A2(
        npu_inst_pe_1_2_0_int_q_weight_1_), .ZN(npu_inst_pe_1_2_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_2_0_U36 ( .A(npu_inst_pe_1_2_0_int_data_1_), .ZN(
        npu_inst_pe_1_2_0_n12) );
  NOR3_X1 npu_inst_pe_1_2_0_U35 ( .A1(npu_inst_pe_1_2_0_n26), .A2(npu_inst_n40), .A3(npu_inst_int_ckg[47]), .ZN(npu_inst_pe_1_2_0_n85) );
  OR2_X1 npu_inst_pe_1_2_0_U34 ( .A1(npu_inst_pe_1_2_0_n85), .A2(
        npu_inst_pe_1_2_0_n1), .ZN(npu_inst_pe_1_2_0_N84) );
  AOI222_X1 npu_inst_pe_1_2_0_U33 ( .A1(npu_inst_int_data_res_3__0__2_), .A2(
        npu_inst_pe_1_2_0_n1), .B1(npu_inst_pe_1_2_0_N75), .B2(
        npu_inst_pe_1_2_0_n76), .C1(npu_inst_pe_1_2_0_N67), .C2(
        npu_inst_pe_1_2_0_n77), .ZN(npu_inst_pe_1_2_0_n82) );
  INV_X1 npu_inst_pe_1_2_0_U32 ( .A(npu_inst_pe_1_2_0_n82), .ZN(
        npu_inst_pe_1_2_0_n36) );
  AOI22_X1 npu_inst_pe_1_2_0_U31 ( .A1(npu_inst_n40), .A2(
        npu_inst_int_data_y_3__0__1_), .B1(npu_inst_pe_1_2_0_n2), .B2(
        npu_inst_int_data_x_2__1__1_), .ZN(npu_inst_pe_1_2_0_n63) );
  AOI22_X1 npu_inst_pe_1_2_0_U30 ( .A1(npu_inst_n40), .A2(
        npu_inst_int_data_y_3__0__0_), .B1(npu_inst_pe_1_2_0_n2), .B2(
        npu_inst_int_data_x_2__1__0_), .ZN(npu_inst_pe_1_2_0_n61) );
  INV_X1 npu_inst_pe_1_2_0_U29 ( .A(npu_inst_pe_1_2_0_int_data_0_), .ZN(
        npu_inst_pe_1_2_0_n11) );
  INV_X1 npu_inst_pe_1_2_0_U28 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_2_0_n4)
         );
  OR3_X1 npu_inst_pe_1_2_0_U27 ( .A1(npu_inst_n60), .A2(npu_inst_pe_1_2_0_n6), 
        .A3(npu_inst_pe_1_2_0_n4), .ZN(npu_inst_pe_1_2_0_n56) );
  OR3_X1 npu_inst_pe_1_2_0_U26 ( .A1(npu_inst_pe_1_2_0_n4), .A2(
        npu_inst_pe_1_2_0_n6), .A3(npu_inst_pe_1_2_0_n5), .ZN(
        npu_inst_pe_1_2_0_n48) );
  INV_X1 npu_inst_pe_1_2_0_U25 ( .A(npu_inst_pe_1_2_0_n4), .ZN(
        npu_inst_pe_1_2_0_n3) );
  OR3_X1 npu_inst_pe_1_2_0_U24 ( .A1(npu_inst_pe_1_2_0_n3), .A2(
        npu_inst_pe_1_2_0_n6), .A3(npu_inst_pe_1_2_0_n5), .ZN(
        npu_inst_pe_1_2_0_n52) );
  OR3_X1 npu_inst_pe_1_2_0_U23 ( .A1(npu_inst_n60), .A2(npu_inst_pe_1_2_0_n6), 
        .A3(npu_inst_pe_1_2_0_n3), .ZN(npu_inst_pe_1_2_0_n60) );
  BUF_X1 npu_inst_pe_1_2_0_U22 ( .A(npu_inst_n26), .Z(npu_inst_pe_1_2_0_n1) );
  NOR2_X1 npu_inst_pe_1_2_0_U21 ( .A1(npu_inst_pe_1_2_0_n60), .A2(
        npu_inst_pe_1_2_0_n2), .ZN(npu_inst_pe_1_2_0_n58) );
  NOR2_X1 npu_inst_pe_1_2_0_U20 ( .A1(npu_inst_pe_1_2_0_n56), .A2(
        npu_inst_pe_1_2_0_n2), .ZN(npu_inst_pe_1_2_0_n54) );
  NOR2_X1 npu_inst_pe_1_2_0_U19 ( .A1(npu_inst_pe_1_2_0_n52), .A2(
        npu_inst_pe_1_2_0_n2), .ZN(npu_inst_pe_1_2_0_n50) );
  NOR2_X1 npu_inst_pe_1_2_0_U18 ( .A1(npu_inst_pe_1_2_0_n48), .A2(
        npu_inst_pe_1_2_0_n2), .ZN(npu_inst_pe_1_2_0_n46) );
  NOR2_X1 npu_inst_pe_1_2_0_U17 ( .A1(npu_inst_pe_1_2_0_n40), .A2(
        npu_inst_pe_1_2_0_n2), .ZN(npu_inst_pe_1_2_0_n38) );
  NOR2_X1 npu_inst_pe_1_2_0_U16 ( .A1(npu_inst_pe_1_2_0_n44), .A2(
        npu_inst_pe_1_2_0_n2), .ZN(npu_inst_pe_1_2_0_n42) );
  BUF_X1 npu_inst_pe_1_2_0_U15 ( .A(npu_inst_n85), .Z(npu_inst_pe_1_2_0_n6) );
  INV_X1 npu_inst_pe_1_2_0_U14 ( .A(npu_inst_n107), .ZN(npu_inst_pe_1_2_0_n10)
         );
  INV_X1 npu_inst_pe_1_2_0_U13 ( .A(npu_inst_pe_1_2_0_n38), .ZN(
        npu_inst_pe_1_2_0_n112) );
  INV_X1 npu_inst_pe_1_2_0_U12 ( .A(npu_inst_pe_1_2_0_n58), .ZN(
        npu_inst_pe_1_2_0_n117) );
  INV_X1 npu_inst_pe_1_2_0_U11 ( .A(npu_inst_pe_1_2_0_n54), .ZN(
        npu_inst_pe_1_2_0_n116) );
  INV_X1 npu_inst_pe_1_2_0_U10 ( .A(npu_inst_pe_1_2_0_n50), .ZN(
        npu_inst_pe_1_2_0_n115) );
  INV_X1 npu_inst_pe_1_2_0_U9 ( .A(npu_inst_pe_1_2_0_n46), .ZN(
        npu_inst_pe_1_2_0_n114) );
  INV_X1 npu_inst_pe_1_2_0_U8 ( .A(npu_inst_pe_1_2_0_n42), .ZN(
        npu_inst_pe_1_2_0_n113) );
  BUF_X1 npu_inst_pe_1_2_0_U7 ( .A(npu_inst_pe_1_2_0_n10), .Z(
        npu_inst_pe_1_2_0_n9) );
  BUF_X1 npu_inst_pe_1_2_0_U6 ( .A(npu_inst_pe_1_2_0_n10), .Z(
        npu_inst_pe_1_2_0_n8) );
  BUF_X1 npu_inst_pe_1_2_0_U5 ( .A(npu_inst_pe_1_2_0_n10), .Z(
        npu_inst_pe_1_2_0_n7) );
  NOR2_X1 npu_inst_pe_1_2_0_U4 ( .A1(npu_inst_pe_1_2_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_0_n1), .ZN(npu_inst_pe_1_2_0_n76) );
  NOR2_X1 npu_inst_pe_1_2_0_U3 ( .A1(npu_inst_pe_1_2_0_n27), .A2(
        npu_inst_pe_1_2_0_n1), .ZN(npu_inst_pe_1_2_0_n77) );
  FA_X1 npu_inst_pe_1_2_0_sub_77_U2_1 ( .A(npu_inst_int_data_res_2__0__1_), 
        .B(npu_inst_pe_1_2_0_n12), .CI(npu_inst_pe_1_2_0_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_2_0_sub_77_carry_2_), .S(npu_inst_pe_1_2_0_N66) );
  FA_X1 npu_inst_pe_1_2_0_add_79_U1_1 ( .A(npu_inst_int_data_res_2__0__1_), 
        .B(npu_inst_pe_1_2_0_int_data_1_), .CI(
        npu_inst_pe_1_2_0_add_79_carry_1_), .CO(
        npu_inst_pe_1_2_0_add_79_carry_2_), .S(npu_inst_pe_1_2_0_N74) );
  NAND3_X1 npu_inst_pe_1_2_0_U101 ( .A1(npu_inst_pe_1_2_0_n4), .A2(
        npu_inst_pe_1_2_0_n5), .A3(npu_inst_pe_1_2_0_n6), .ZN(
        npu_inst_pe_1_2_0_n44) );
  NAND3_X1 npu_inst_pe_1_2_0_U100 ( .A1(npu_inst_pe_1_2_0_n3), .A2(
        npu_inst_pe_1_2_0_n5), .A3(npu_inst_pe_1_2_0_n6), .ZN(
        npu_inst_pe_1_2_0_n40) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_0_n32), .CK(
        npu_inst_pe_1_2_0_net4110), .RN(npu_inst_pe_1_2_0_n7), .Q(
        npu_inst_int_data_res_2__0__6_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_0_n33), .CK(
        npu_inst_pe_1_2_0_net4110), .RN(npu_inst_pe_1_2_0_n7), .Q(
        npu_inst_int_data_res_2__0__5_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_0_n34), .CK(
        npu_inst_pe_1_2_0_net4110), .RN(npu_inst_pe_1_2_0_n7), .Q(
        npu_inst_int_data_res_2__0__4_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_0_n35), .CK(
        npu_inst_pe_1_2_0_net4110), .RN(npu_inst_pe_1_2_0_n7), .Q(
        npu_inst_int_data_res_2__0__3_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_0_n36), .CK(
        npu_inst_pe_1_2_0_net4110), .RN(npu_inst_pe_1_2_0_n7), .Q(
        npu_inst_int_data_res_2__0__2_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_0_n98), .CK(
        npu_inst_pe_1_2_0_net4110), .RN(npu_inst_pe_1_2_0_n7), .Q(
        npu_inst_int_data_res_2__0__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_0_n31), .CK(
        npu_inst_pe_1_2_0_net4110), .RN(npu_inst_pe_1_2_0_n7), .Q(
        npu_inst_int_data_res_2__0__7_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_0_n99), .CK(
        npu_inst_pe_1_2_0_net4110), .RN(npu_inst_pe_1_2_0_n7), .Q(
        npu_inst_int_data_res_2__0__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_weight_reg_0_ ( .D(npu_inst_n93), .CK(
        npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n7), .Q(
        npu_inst_pe_1_2_0_int_q_weight_0_), .QN(npu_inst_pe_1_2_0_n27) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_weight_reg_1_ ( .D(npu_inst_n99), .CK(
        npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n7), .Q(
        npu_inst_pe_1_2_0_int_q_weight_1_), .QN(npu_inst_pe_1_2_0_n26) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_0_n111), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n7), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_0_n105), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n7), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_0_n110), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_0_n104), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_0_n109), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_0_n103), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_0_n108), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_0_n102), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_0_n107), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_0_n101), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_0_n106), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_0_n100), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_0_n86), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_0_n87), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n8), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_0_n88), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_0_n89), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_0_n90), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_0_n91), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_0_n92), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_0_n93), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_0_n94), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_0_n95), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_0_n96), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_0_n97), 
        .CK(npu_inst_pe_1_2_0_net4116), .RN(npu_inst_pe_1_2_0_n9), .Q(
        npu_inst_pe_1_2_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_0_net4110) );
  CLKGATETST_X1 npu_inst_pe_1_2_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n47), .SE(1'b0), .GCK(npu_inst_pe_1_2_0_net4116) );
  MUX2_X1 npu_inst_pe_1_2_1_U153 ( .A(npu_inst_pe_1_2_1_n31), .B(
        npu_inst_pe_1_2_1_n28), .S(npu_inst_pe_1_2_1_n7), .Z(
        npu_inst_pe_1_2_1_N93) );
  MUX2_X1 npu_inst_pe_1_2_1_U152 ( .A(npu_inst_pe_1_2_1_n30), .B(
        npu_inst_pe_1_2_1_n29), .S(npu_inst_pe_1_2_1_n5), .Z(
        npu_inst_pe_1_2_1_n31) );
  MUX2_X1 npu_inst_pe_1_2_1_U151 ( .A(npu_inst_pe_1_2_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_1_n3), .Z(
        npu_inst_pe_1_2_1_n30) );
  MUX2_X1 npu_inst_pe_1_2_1_U150 ( .A(npu_inst_pe_1_2_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_1_n3), .Z(
        npu_inst_pe_1_2_1_n29) );
  MUX2_X1 npu_inst_pe_1_2_1_U149 ( .A(npu_inst_pe_1_2_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_1_n3), .Z(
        npu_inst_pe_1_2_1_n28) );
  MUX2_X1 npu_inst_pe_1_2_1_U148 ( .A(npu_inst_pe_1_2_1_n25), .B(
        npu_inst_pe_1_2_1_n22), .S(npu_inst_pe_1_2_1_n7), .Z(
        npu_inst_pe_1_2_1_N94) );
  MUX2_X1 npu_inst_pe_1_2_1_U147 ( .A(npu_inst_pe_1_2_1_n24), .B(
        npu_inst_pe_1_2_1_n23), .S(npu_inst_pe_1_2_1_n5), .Z(
        npu_inst_pe_1_2_1_n25) );
  MUX2_X1 npu_inst_pe_1_2_1_U146 ( .A(npu_inst_pe_1_2_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_1_n3), .Z(
        npu_inst_pe_1_2_1_n24) );
  MUX2_X1 npu_inst_pe_1_2_1_U145 ( .A(npu_inst_pe_1_2_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_1_n3), .Z(
        npu_inst_pe_1_2_1_n23) );
  MUX2_X1 npu_inst_pe_1_2_1_U144 ( .A(npu_inst_pe_1_2_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_1_n3), .Z(
        npu_inst_pe_1_2_1_n22) );
  MUX2_X1 npu_inst_pe_1_2_1_U143 ( .A(npu_inst_pe_1_2_1_n21), .B(
        npu_inst_pe_1_2_1_n18), .S(npu_inst_pe_1_2_1_n7), .Z(
        npu_inst_int_data_x_2__1__1_) );
  MUX2_X1 npu_inst_pe_1_2_1_U142 ( .A(npu_inst_pe_1_2_1_n20), .B(
        npu_inst_pe_1_2_1_n19), .S(npu_inst_pe_1_2_1_n5), .Z(
        npu_inst_pe_1_2_1_n21) );
  MUX2_X1 npu_inst_pe_1_2_1_U141 ( .A(npu_inst_pe_1_2_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_1_n3), .Z(
        npu_inst_pe_1_2_1_n20) );
  MUX2_X1 npu_inst_pe_1_2_1_U140 ( .A(npu_inst_pe_1_2_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_1_n3), .Z(
        npu_inst_pe_1_2_1_n19) );
  MUX2_X1 npu_inst_pe_1_2_1_U139 ( .A(npu_inst_pe_1_2_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_1_n3), .Z(
        npu_inst_pe_1_2_1_n18) );
  MUX2_X1 npu_inst_pe_1_2_1_U138 ( .A(npu_inst_pe_1_2_1_n17), .B(
        npu_inst_pe_1_2_1_n14), .S(npu_inst_pe_1_2_1_n7), .Z(
        npu_inst_int_data_x_2__1__0_) );
  MUX2_X1 npu_inst_pe_1_2_1_U137 ( .A(npu_inst_pe_1_2_1_n16), .B(
        npu_inst_pe_1_2_1_n15), .S(npu_inst_pe_1_2_1_n5), .Z(
        npu_inst_pe_1_2_1_n17) );
  MUX2_X1 npu_inst_pe_1_2_1_U136 ( .A(npu_inst_pe_1_2_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_1_n3), .Z(
        npu_inst_pe_1_2_1_n16) );
  MUX2_X1 npu_inst_pe_1_2_1_U135 ( .A(npu_inst_pe_1_2_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_1_n3), .Z(
        npu_inst_pe_1_2_1_n15) );
  MUX2_X1 npu_inst_pe_1_2_1_U134 ( .A(npu_inst_pe_1_2_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_1_n3), .Z(
        npu_inst_pe_1_2_1_n14) );
  XOR2_X1 npu_inst_pe_1_2_1_U133 ( .A(npu_inst_pe_1_2_1_int_data_0_), .B(
        npu_inst_int_data_res_2__1__0_), .Z(npu_inst_pe_1_2_1_N73) );
  AND2_X1 npu_inst_pe_1_2_1_U132 ( .A1(npu_inst_int_data_res_2__1__0_), .A2(
        npu_inst_pe_1_2_1_int_data_0_), .ZN(npu_inst_pe_1_2_1_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_1_U131 ( .A(npu_inst_int_data_res_2__1__0_), .B(
        npu_inst_pe_1_2_1_n12), .ZN(npu_inst_pe_1_2_1_N65) );
  OR2_X1 npu_inst_pe_1_2_1_U130 ( .A1(npu_inst_pe_1_2_1_n12), .A2(
        npu_inst_int_data_res_2__1__0_), .ZN(npu_inst_pe_1_2_1_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_1_U129 ( .A(npu_inst_int_data_res_2__1__2_), .B(
        npu_inst_pe_1_2_1_add_79_carry_2_), .Z(npu_inst_pe_1_2_1_N75) );
  AND2_X1 npu_inst_pe_1_2_1_U128 ( .A1(npu_inst_pe_1_2_1_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_2__1__2_), .ZN(
        npu_inst_pe_1_2_1_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_1_U127 ( .A(npu_inst_int_data_res_2__1__3_), .B(
        npu_inst_pe_1_2_1_add_79_carry_3_), .Z(npu_inst_pe_1_2_1_N76) );
  AND2_X1 npu_inst_pe_1_2_1_U126 ( .A1(npu_inst_pe_1_2_1_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_2__1__3_), .ZN(
        npu_inst_pe_1_2_1_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_1_U125 ( .A(npu_inst_int_data_res_2__1__4_), .B(
        npu_inst_pe_1_2_1_add_79_carry_4_), .Z(npu_inst_pe_1_2_1_N77) );
  AND2_X1 npu_inst_pe_1_2_1_U124 ( .A1(npu_inst_pe_1_2_1_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_2__1__4_), .ZN(
        npu_inst_pe_1_2_1_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_1_U123 ( .A(npu_inst_int_data_res_2__1__5_), .B(
        npu_inst_pe_1_2_1_add_79_carry_5_), .Z(npu_inst_pe_1_2_1_N78) );
  AND2_X1 npu_inst_pe_1_2_1_U122 ( .A1(npu_inst_pe_1_2_1_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_2__1__5_), .ZN(
        npu_inst_pe_1_2_1_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_1_U121 ( .A(npu_inst_int_data_res_2__1__6_), .B(
        npu_inst_pe_1_2_1_add_79_carry_6_), .Z(npu_inst_pe_1_2_1_N79) );
  AND2_X1 npu_inst_pe_1_2_1_U120 ( .A1(npu_inst_pe_1_2_1_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_2__1__6_), .ZN(
        npu_inst_pe_1_2_1_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_1_U119 ( .A(npu_inst_int_data_res_2__1__7_), .B(
        npu_inst_pe_1_2_1_add_79_carry_7_), .Z(npu_inst_pe_1_2_1_N80) );
  XNOR2_X1 npu_inst_pe_1_2_1_U118 ( .A(npu_inst_pe_1_2_1_sub_77_carry_2_), .B(
        npu_inst_int_data_res_2__1__2_), .ZN(npu_inst_pe_1_2_1_N67) );
  OR2_X1 npu_inst_pe_1_2_1_U117 ( .A1(npu_inst_int_data_res_2__1__2_), .A2(
        npu_inst_pe_1_2_1_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_2_1_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_1_U116 ( .A(npu_inst_pe_1_2_1_sub_77_carry_3_), .B(
        npu_inst_int_data_res_2__1__3_), .ZN(npu_inst_pe_1_2_1_N68) );
  OR2_X1 npu_inst_pe_1_2_1_U115 ( .A1(npu_inst_int_data_res_2__1__3_), .A2(
        npu_inst_pe_1_2_1_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_2_1_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_1_U114 ( .A(npu_inst_pe_1_2_1_sub_77_carry_4_), .B(
        npu_inst_int_data_res_2__1__4_), .ZN(npu_inst_pe_1_2_1_N69) );
  OR2_X1 npu_inst_pe_1_2_1_U113 ( .A1(npu_inst_int_data_res_2__1__4_), .A2(
        npu_inst_pe_1_2_1_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_2_1_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_1_U112 ( .A(npu_inst_pe_1_2_1_sub_77_carry_5_), .B(
        npu_inst_int_data_res_2__1__5_), .ZN(npu_inst_pe_1_2_1_N70) );
  OR2_X1 npu_inst_pe_1_2_1_U111 ( .A1(npu_inst_int_data_res_2__1__5_), .A2(
        npu_inst_pe_1_2_1_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_2_1_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_1_U110 ( .A(npu_inst_pe_1_2_1_sub_77_carry_6_), .B(
        npu_inst_int_data_res_2__1__6_), .ZN(npu_inst_pe_1_2_1_N71) );
  OR2_X1 npu_inst_pe_1_2_1_U109 ( .A1(npu_inst_int_data_res_2__1__6_), .A2(
        npu_inst_pe_1_2_1_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_2_1_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_1_U108 ( .A(npu_inst_int_data_res_2__1__7_), .B(
        npu_inst_pe_1_2_1_sub_77_carry_7_), .ZN(npu_inst_pe_1_2_1_N72) );
  INV_X1 npu_inst_pe_1_2_1_U107 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_2_1_n6)
         );
  INV_X1 npu_inst_pe_1_2_1_U106 ( .A(npu_inst_pe_1_2_1_n6), .ZN(
        npu_inst_pe_1_2_1_n5) );
  INV_X1 npu_inst_pe_1_2_1_U105 ( .A(npu_inst_n40), .ZN(npu_inst_pe_1_2_1_n2)
         );
  AOI22_X1 npu_inst_pe_1_2_1_U104 ( .A1(npu_inst_int_data_y_3__1__0_), .A2(
        npu_inst_pe_1_2_1_n58), .B1(npu_inst_pe_1_2_1_n118), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_1_n57) );
  INV_X1 npu_inst_pe_1_2_1_U103 ( .A(npu_inst_pe_1_2_1_n57), .ZN(
        npu_inst_pe_1_2_1_n107) );
  AOI22_X1 npu_inst_pe_1_2_1_U102 ( .A1(npu_inst_int_data_y_3__1__0_), .A2(
        npu_inst_pe_1_2_1_n54), .B1(npu_inst_pe_1_2_1_n117), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_1_n53) );
  INV_X1 npu_inst_pe_1_2_1_U99 ( .A(npu_inst_pe_1_2_1_n53), .ZN(
        npu_inst_pe_1_2_1_n108) );
  AOI22_X1 npu_inst_pe_1_2_1_U98 ( .A1(npu_inst_int_data_y_3__1__0_), .A2(
        npu_inst_pe_1_2_1_n50), .B1(npu_inst_pe_1_2_1_n116), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_1_n49) );
  INV_X1 npu_inst_pe_1_2_1_U97 ( .A(npu_inst_pe_1_2_1_n49), .ZN(
        npu_inst_pe_1_2_1_n109) );
  AOI22_X1 npu_inst_pe_1_2_1_U96 ( .A1(npu_inst_int_data_y_3__1__0_), .A2(
        npu_inst_pe_1_2_1_n46), .B1(npu_inst_pe_1_2_1_n115), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_1_n45) );
  INV_X1 npu_inst_pe_1_2_1_U95 ( .A(npu_inst_pe_1_2_1_n45), .ZN(
        npu_inst_pe_1_2_1_n110) );
  AOI22_X1 npu_inst_pe_1_2_1_U94 ( .A1(npu_inst_int_data_y_3__1__0_), .A2(
        npu_inst_pe_1_2_1_n42), .B1(npu_inst_pe_1_2_1_n114), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_1_n41) );
  INV_X1 npu_inst_pe_1_2_1_U93 ( .A(npu_inst_pe_1_2_1_n41), .ZN(
        npu_inst_pe_1_2_1_n111) );
  AOI22_X1 npu_inst_pe_1_2_1_U92 ( .A1(npu_inst_int_data_y_3__1__1_), .A2(
        npu_inst_pe_1_2_1_n58), .B1(npu_inst_pe_1_2_1_n118), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_1_n59) );
  INV_X1 npu_inst_pe_1_2_1_U91 ( .A(npu_inst_pe_1_2_1_n59), .ZN(
        npu_inst_pe_1_2_1_n101) );
  AOI22_X1 npu_inst_pe_1_2_1_U90 ( .A1(npu_inst_int_data_y_3__1__1_), .A2(
        npu_inst_pe_1_2_1_n54), .B1(npu_inst_pe_1_2_1_n117), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_1_n55) );
  INV_X1 npu_inst_pe_1_2_1_U89 ( .A(npu_inst_pe_1_2_1_n55), .ZN(
        npu_inst_pe_1_2_1_n102) );
  AOI22_X1 npu_inst_pe_1_2_1_U88 ( .A1(npu_inst_int_data_y_3__1__1_), .A2(
        npu_inst_pe_1_2_1_n50), .B1(npu_inst_pe_1_2_1_n116), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_1_n51) );
  INV_X1 npu_inst_pe_1_2_1_U87 ( .A(npu_inst_pe_1_2_1_n51), .ZN(
        npu_inst_pe_1_2_1_n103) );
  AOI22_X1 npu_inst_pe_1_2_1_U86 ( .A1(npu_inst_int_data_y_3__1__1_), .A2(
        npu_inst_pe_1_2_1_n46), .B1(npu_inst_pe_1_2_1_n115), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_1_n47) );
  INV_X1 npu_inst_pe_1_2_1_U85 ( .A(npu_inst_pe_1_2_1_n47), .ZN(
        npu_inst_pe_1_2_1_n104) );
  AOI22_X1 npu_inst_pe_1_2_1_U84 ( .A1(npu_inst_int_data_y_3__1__1_), .A2(
        npu_inst_pe_1_2_1_n42), .B1(npu_inst_pe_1_2_1_n114), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_1_n43) );
  INV_X1 npu_inst_pe_1_2_1_U83 ( .A(npu_inst_pe_1_2_1_n43), .ZN(
        npu_inst_pe_1_2_1_n105) );
  AOI22_X1 npu_inst_pe_1_2_1_U82 ( .A1(npu_inst_pe_1_2_1_n38), .A2(
        npu_inst_int_data_y_3__1__1_), .B1(npu_inst_pe_1_2_1_n113), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_1_n39) );
  INV_X1 npu_inst_pe_1_2_1_U81 ( .A(npu_inst_pe_1_2_1_n39), .ZN(
        npu_inst_pe_1_2_1_n106) );
  AND2_X1 npu_inst_pe_1_2_1_U80 ( .A1(npu_inst_pe_1_2_1_N93), .A2(npu_inst_n40), .ZN(npu_inst_int_data_y_2__1__0_) );
  NAND2_X1 npu_inst_pe_1_2_1_U79 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_1_n60), .ZN(npu_inst_pe_1_2_1_n74) );
  OAI21_X1 npu_inst_pe_1_2_1_U78 ( .B1(npu_inst_pe_1_2_1_n63), .B2(
        npu_inst_pe_1_2_1_n60), .A(npu_inst_pe_1_2_1_n74), .ZN(
        npu_inst_pe_1_2_1_n97) );
  NAND2_X1 npu_inst_pe_1_2_1_U77 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_1_n60), .ZN(npu_inst_pe_1_2_1_n73) );
  OAI21_X1 npu_inst_pe_1_2_1_U76 ( .B1(npu_inst_pe_1_2_1_n61), .B2(
        npu_inst_pe_1_2_1_n60), .A(npu_inst_pe_1_2_1_n73), .ZN(
        npu_inst_pe_1_2_1_n96) );
  NAND2_X1 npu_inst_pe_1_2_1_U75 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_1_n56), .ZN(npu_inst_pe_1_2_1_n72) );
  OAI21_X1 npu_inst_pe_1_2_1_U74 ( .B1(npu_inst_pe_1_2_1_n63), .B2(
        npu_inst_pe_1_2_1_n56), .A(npu_inst_pe_1_2_1_n72), .ZN(
        npu_inst_pe_1_2_1_n95) );
  NAND2_X1 npu_inst_pe_1_2_1_U73 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_1_n56), .ZN(npu_inst_pe_1_2_1_n71) );
  OAI21_X1 npu_inst_pe_1_2_1_U72 ( .B1(npu_inst_pe_1_2_1_n61), .B2(
        npu_inst_pe_1_2_1_n56), .A(npu_inst_pe_1_2_1_n71), .ZN(
        npu_inst_pe_1_2_1_n94) );
  NAND2_X1 npu_inst_pe_1_2_1_U71 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_1_n52), .ZN(npu_inst_pe_1_2_1_n70) );
  OAI21_X1 npu_inst_pe_1_2_1_U70 ( .B1(npu_inst_pe_1_2_1_n63), .B2(
        npu_inst_pe_1_2_1_n52), .A(npu_inst_pe_1_2_1_n70), .ZN(
        npu_inst_pe_1_2_1_n93) );
  NAND2_X1 npu_inst_pe_1_2_1_U69 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_1_n52), .ZN(npu_inst_pe_1_2_1_n69) );
  OAI21_X1 npu_inst_pe_1_2_1_U68 ( .B1(npu_inst_pe_1_2_1_n61), .B2(
        npu_inst_pe_1_2_1_n52), .A(npu_inst_pe_1_2_1_n69), .ZN(
        npu_inst_pe_1_2_1_n92) );
  NAND2_X1 npu_inst_pe_1_2_1_U67 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_1_n48), .ZN(npu_inst_pe_1_2_1_n68) );
  OAI21_X1 npu_inst_pe_1_2_1_U66 ( .B1(npu_inst_pe_1_2_1_n63), .B2(
        npu_inst_pe_1_2_1_n48), .A(npu_inst_pe_1_2_1_n68), .ZN(
        npu_inst_pe_1_2_1_n91) );
  NAND2_X1 npu_inst_pe_1_2_1_U65 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_1_n48), .ZN(npu_inst_pe_1_2_1_n67) );
  OAI21_X1 npu_inst_pe_1_2_1_U64 ( .B1(npu_inst_pe_1_2_1_n61), .B2(
        npu_inst_pe_1_2_1_n48), .A(npu_inst_pe_1_2_1_n67), .ZN(
        npu_inst_pe_1_2_1_n90) );
  NAND2_X1 npu_inst_pe_1_2_1_U63 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_1_n44), .ZN(npu_inst_pe_1_2_1_n66) );
  OAI21_X1 npu_inst_pe_1_2_1_U62 ( .B1(npu_inst_pe_1_2_1_n63), .B2(
        npu_inst_pe_1_2_1_n44), .A(npu_inst_pe_1_2_1_n66), .ZN(
        npu_inst_pe_1_2_1_n89) );
  NAND2_X1 npu_inst_pe_1_2_1_U61 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_1_n44), .ZN(npu_inst_pe_1_2_1_n65) );
  OAI21_X1 npu_inst_pe_1_2_1_U60 ( .B1(npu_inst_pe_1_2_1_n61), .B2(
        npu_inst_pe_1_2_1_n44), .A(npu_inst_pe_1_2_1_n65), .ZN(
        npu_inst_pe_1_2_1_n88) );
  NAND2_X1 npu_inst_pe_1_2_1_U59 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_1_n40), .ZN(npu_inst_pe_1_2_1_n64) );
  OAI21_X1 npu_inst_pe_1_2_1_U58 ( .B1(npu_inst_pe_1_2_1_n63), .B2(
        npu_inst_pe_1_2_1_n40), .A(npu_inst_pe_1_2_1_n64), .ZN(
        npu_inst_pe_1_2_1_n87) );
  NAND2_X1 npu_inst_pe_1_2_1_U57 ( .A1(npu_inst_pe_1_2_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_1_n40), .ZN(npu_inst_pe_1_2_1_n62) );
  OAI21_X1 npu_inst_pe_1_2_1_U56 ( .B1(npu_inst_pe_1_2_1_n61), .B2(
        npu_inst_pe_1_2_1_n40), .A(npu_inst_pe_1_2_1_n62), .ZN(
        npu_inst_pe_1_2_1_n86) );
  AOI22_X1 npu_inst_pe_1_2_1_U55 ( .A1(npu_inst_pe_1_2_1_n38), .A2(
        npu_inst_int_data_y_3__1__0_), .B1(npu_inst_pe_1_2_1_n113), .B2(
        npu_inst_pe_1_2_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_1_n37) );
  INV_X1 npu_inst_pe_1_2_1_U54 ( .A(npu_inst_pe_1_2_1_n37), .ZN(
        npu_inst_pe_1_2_1_n112) );
  AND2_X1 npu_inst_pe_1_2_1_U53 ( .A1(npu_inst_n40), .A2(npu_inst_pe_1_2_1_N94), .ZN(npu_inst_int_data_y_2__1__1_) );
  AOI222_X1 npu_inst_pe_1_2_1_U52 ( .A1(npu_inst_int_data_res_3__1__0_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N73), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N65), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n84) );
  INV_X1 npu_inst_pe_1_2_1_U51 ( .A(npu_inst_pe_1_2_1_n84), .ZN(
        npu_inst_pe_1_2_1_n100) );
  AOI222_X1 npu_inst_pe_1_2_1_U50 ( .A1(npu_inst_pe_1_2_1_n1), .A2(
        npu_inst_int_data_res_3__1__7_), .B1(npu_inst_pe_1_2_1_N80), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N72), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n75) );
  INV_X1 npu_inst_pe_1_2_1_U49 ( .A(npu_inst_pe_1_2_1_n75), .ZN(
        npu_inst_pe_1_2_1_n32) );
  AOI222_X1 npu_inst_pe_1_2_1_U48 ( .A1(npu_inst_int_data_res_3__1__1_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N74), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N66), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n83) );
  INV_X1 npu_inst_pe_1_2_1_U47 ( .A(npu_inst_pe_1_2_1_n83), .ZN(
        npu_inst_pe_1_2_1_n99) );
  AOI222_X1 npu_inst_pe_1_2_1_U46 ( .A1(npu_inst_int_data_res_3__1__3_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N76), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N68), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n81) );
  INV_X1 npu_inst_pe_1_2_1_U45 ( .A(npu_inst_pe_1_2_1_n81), .ZN(
        npu_inst_pe_1_2_1_n36) );
  AOI222_X1 npu_inst_pe_1_2_1_U44 ( .A1(npu_inst_int_data_res_3__1__4_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N77), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N69), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n80) );
  INV_X1 npu_inst_pe_1_2_1_U43 ( .A(npu_inst_pe_1_2_1_n80), .ZN(
        npu_inst_pe_1_2_1_n35) );
  AOI222_X1 npu_inst_pe_1_2_1_U42 ( .A1(npu_inst_int_data_res_3__1__5_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N78), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N70), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n79) );
  INV_X1 npu_inst_pe_1_2_1_U41 ( .A(npu_inst_pe_1_2_1_n79), .ZN(
        npu_inst_pe_1_2_1_n34) );
  AOI222_X1 npu_inst_pe_1_2_1_U40 ( .A1(npu_inst_int_data_res_3__1__6_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N79), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N71), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n78) );
  INV_X1 npu_inst_pe_1_2_1_U39 ( .A(npu_inst_pe_1_2_1_n78), .ZN(
        npu_inst_pe_1_2_1_n33) );
  AND2_X1 npu_inst_pe_1_2_1_U38 ( .A1(npu_inst_int_data_x_2__1__1_), .A2(
        npu_inst_pe_1_2_1_int_q_weight_1_), .ZN(npu_inst_pe_1_2_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_1_U37 ( .A1(npu_inst_int_data_x_2__1__0_), .A2(
        npu_inst_pe_1_2_1_int_q_weight_1_), .ZN(npu_inst_pe_1_2_1_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_2_1_U36 ( .A(npu_inst_pe_1_2_1_int_data_1_), .ZN(
        npu_inst_pe_1_2_1_n13) );
  NOR3_X1 npu_inst_pe_1_2_1_U35 ( .A1(npu_inst_pe_1_2_1_n26), .A2(npu_inst_n40), .A3(npu_inst_int_ckg[46]), .ZN(npu_inst_pe_1_2_1_n85) );
  OR2_X1 npu_inst_pe_1_2_1_U34 ( .A1(npu_inst_pe_1_2_1_n85), .A2(
        npu_inst_pe_1_2_1_n1), .ZN(npu_inst_pe_1_2_1_N84) );
  AOI222_X1 npu_inst_pe_1_2_1_U33 ( .A1(npu_inst_int_data_res_3__1__2_), .A2(
        npu_inst_pe_1_2_1_n1), .B1(npu_inst_pe_1_2_1_N75), .B2(
        npu_inst_pe_1_2_1_n76), .C1(npu_inst_pe_1_2_1_N67), .C2(
        npu_inst_pe_1_2_1_n77), .ZN(npu_inst_pe_1_2_1_n82) );
  INV_X1 npu_inst_pe_1_2_1_U32 ( .A(npu_inst_pe_1_2_1_n82), .ZN(
        npu_inst_pe_1_2_1_n98) );
  AOI22_X1 npu_inst_pe_1_2_1_U31 ( .A1(npu_inst_n40), .A2(
        npu_inst_int_data_y_3__1__1_), .B1(npu_inst_pe_1_2_1_n2), .B2(
        npu_inst_int_data_x_2__2__1_), .ZN(npu_inst_pe_1_2_1_n63) );
  AOI22_X1 npu_inst_pe_1_2_1_U30 ( .A1(npu_inst_n40), .A2(
        npu_inst_int_data_y_3__1__0_), .B1(npu_inst_pe_1_2_1_n2), .B2(
        npu_inst_int_data_x_2__2__0_), .ZN(npu_inst_pe_1_2_1_n61) );
  INV_X1 npu_inst_pe_1_2_1_U29 ( .A(npu_inst_pe_1_2_1_int_data_0_), .ZN(
        npu_inst_pe_1_2_1_n12) );
  INV_X1 npu_inst_pe_1_2_1_U28 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_2_1_n4)
         );
  OR3_X1 npu_inst_pe_1_2_1_U27 ( .A1(npu_inst_pe_1_2_1_n5), .A2(
        npu_inst_pe_1_2_1_n7), .A3(npu_inst_pe_1_2_1_n4), .ZN(
        npu_inst_pe_1_2_1_n56) );
  OR3_X1 npu_inst_pe_1_2_1_U26 ( .A1(npu_inst_pe_1_2_1_n4), .A2(
        npu_inst_pe_1_2_1_n7), .A3(npu_inst_pe_1_2_1_n6), .ZN(
        npu_inst_pe_1_2_1_n48) );
  INV_X1 npu_inst_pe_1_2_1_U25 ( .A(npu_inst_pe_1_2_1_n4), .ZN(
        npu_inst_pe_1_2_1_n3) );
  OR3_X1 npu_inst_pe_1_2_1_U24 ( .A1(npu_inst_pe_1_2_1_n3), .A2(
        npu_inst_pe_1_2_1_n7), .A3(npu_inst_pe_1_2_1_n6), .ZN(
        npu_inst_pe_1_2_1_n52) );
  OR3_X1 npu_inst_pe_1_2_1_U23 ( .A1(npu_inst_pe_1_2_1_n5), .A2(
        npu_inst_pe_1_2_1_n7), .A3(npu_inst_pe_1_2_1_n3), .ZN(
        npu_inst_pe_1_2_1_n60) );
  BUF_X1 npu_inst_pe_1_2_1_U22 ( .A(npu_inst_n26), .Z(npu_inst_pe_1_2_1_n1) );
  NOR2_X1 npu_inst_pe_1_2_1_U21 ( .A1(npu_inst_pe_1_2_1_n60), .A2(
        npu_inst_pe_1_2_1_n2), .ZN(npu_inst_pe_1_2_1_n58) );
  NOR2_X1 npu_inst_pe_1_2_1_U20 ( .A1(npu_inst_pe_1_2_1_n56), .A2(
        npu_inst_pe_1_2_1_n2), .ZN(npu_inst_pe_1_2_1_n54) );
  NOR2_X1 npu_inst_pe_1_2_1_U19 ( .A1(npu_inst_pe_1_2_1_n52), .A2(
        npu_inst_pe_1_2_1_n2), .ZN(npu_inst_pe_1_2_1_n50) );
  NOR2_X1 npu_inst_pe_1_2_1_U18 ( .A1(npu_inst_pe_1_2_1_n48), .A2(
        npu_inst_pe_1_2_1_n2), .ZN(npu_inst_pe_1_2_1_n46) );
  NOR2_X1 npu_inst_pe_1_2_1_U17 ( .A1(npu_inst_pe_1_2_1_n40), .A2(
        npu_inst_pe_1_2_1_n2), .ZN(npu_inst_pe_1_2_1_n38) );
  NOR2_X1 npu_inst_pe_1_2_1_U16 ( .A1(npu_inst_pe_1_2_1_n44), .A2(
        npu_inst_pe_1_2_1_n2), .ZN(npu_inst_pe_1_2_1_n42) );
  BUF_X1 npu_inst_pe_1_2_1_U15 ( .A(npu_inst_n85), .Z(npu_inst_pe_1_2_1_n7) );
  INV_X1 npu_inst_pe_1_2_1_U14 ( .A(npu_inst_n107), .ZN(npu_inst_pe_1_2_1_n11)
         );
  INV_X1 npu_inst_pe_1_2_1_U13 ( .A(npu_inst_pe_1_2_1_n38), .ZN(
        npu_inst_pe_1_2_1_n113) );
  INV_X1 npu_inst_pe_1_2_1_U12 ( .A(npu_inst_pe_1_2_1_n58), .ZN(
        npu_inst_pe_1_2_1_n118) );
  INV_X1 npu_inst_pe_1_2_1_U11 ( .A(npu_inst_pe_1_2_1_n54), .ZN(
        npu_inst_pe_1_2_1_n117) );
  INV_X1 npu_inst_pe_1_2_1_U10 ( .A(npu_inst_pe_1_2_1_n50), .ZN(
        npu_inst_pe_1_2_1_n116) );
  INV_X1 npu_inst_pe_1_2_1_U9 ( .A(npu_inst_pe_1_2_1_n46), .ZN(
        npu_inst_pe_1_2_1_n115) );
  INV_X1 npu_inst_pe_1_2_1_U8 ( .A(npu_inst_pe_1_2_1_n42), .ZN(
        npu_inst_pe_1_2_1_n114) );
  BUF_X1 npu_inst_pe_1_2_1_U7 ( .A(npu_inst_pe_1_2_1_n11), .Z(
        npu_inst_pe_1_2_1_n10) );
  BUF_X1 npu_inst_pe_1_2_1_U6 ( .A(npu_inst_pe_1_2_1_n11), .Z(
        npu_inst_pe_1_2_1_n9) );
  BUF_X1 npu_inst_pe_1_2_1_U5 ( .A(npu_inst_pe_1_2_1_n11), .Z(
        npu_inst_pe_1_2_1_n8) );
  NOR2_X1 npu_inst_pe_1_2_1_U4 ( .A1(npu_inst_pe_1_2_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_1_n1), .ZN(npu_inst_pe_1_2_1_n76) );
  NOR2_X1 npu_inst_pe_1_2_1_U3 ( .A1(npu_inst_pe_1_2_1_n27), .A2(
        npu_inst_pe_1_2_1_n1), .ZN(npu_inst_pe_1_2_1_n77) );
  FA_X1 npu_inst_pe_1_2_1_sub_77_U2_1 ( .A(npu_inst_int_data_res_2__1__1_), 
        .B(npu_inst_pe_1_2_1_n13), .CI(npu_inst_pe_1_2_1_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_2_1_sub_77_carry_2_), .S(npu_inst_pe_1_2_1_N66) );
  FA_X1 npu_inst_pe_1_2_1_add_79_U1_1 ( .A(npu_inst_int_data_res_2__1__1_), 
        .B(npu_inst_pe_1_2_1_int_data_1_), .CI(
        npu_inst_pe_1_2_1_add_79_carry_1_), .CO(
        npu_inst_pe_1_2_1_add_79_carry_2_), .S(npu_inst_pe_1_2_1_N74) );
  NAND3_X1 npu_inst_pe_1_2_1_U101 ( .A1(npu_inst_pe_1_2_1_n4), .A2(
        npu_inst_pe_1_2_1_n6), .A3(npu_inst_pe_1_2_1_n7), .ZN(
        npu_inst_pe_1_2_1_n44) );
  NAND3_X1 npu_inst_pe_1_2_1_U100 ( .A1(npu_inst_pe_1_2_1_n3), .A2(
        npu_inst_pe_1_2_1_n6), .A3(npu_inst_pe_1_2_1_n7), .ZN(
        npu_inst_pe_1_2_1_n40) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_1_n33), .CK(
        npu_inst_pe_1_2_1_net4087), .RN(npu_inst_pe_1_2_1_n8), .Q(
        npu_inst_int_data_res_2__1__6_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_1_n34), .CK(
        npu_inst_pe_1_2_1_net4087), .RN(npu_inst_pe_1_2_1_n8), .Q(
        npu_inst_int_data_res_2__1__5_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_1_n35), .CK(
        npu_inst_pe_1_2_1_net4087), .RN(npu_inst_pe_1_2_1_n8), .Q(
        npu_inst_int_data_res_2__1__4_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_1_n36), .CK(
        npu_inst_pe_1_2_1_net4087), .RN(npu_inst_pe_1_2_1_n8), .Q(
        npu_inst_int_data_res_2__1__3_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_1_n98), .CK(
        npu_inst_pe_1_2_1_net4087), .RN(npu_inst_pe_1_2_1_n8), .Q(
        npu_inst_int_data_res_2__1__2_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_1_n99), .CK(
        npu_inst_pe_1_2_1_net4087), .RN(npu_inst_pe_1_2_1_n8), .Q(
        npu_inst_int_data_res_2__1__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_1_n32), .CK(
        npu_inst_pe_1_2_1_net4087), .RN(npu_inst_pe_1_2_1_n8), .Q(
        npu_inst_int_data_res_2__1__7_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_1_n100), 
        .CK(npu_inst_pe_1_2_1_net4087), .RN(npu_inst_pe_1_2_1_n8), .Q(
        npu_inst_int_data_res_2__1__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_weight_reg_0_ ( .D(npu_inst_n93), .CK(
        npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n8), .Q(
        npu_inst_pe_1_2_1_int_q_weight_0_), .QN(npu_inst_pe_1_2_1_n27) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_weight_reg_1_ ( .D(npu_inst_n99), .CK(
        npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n8), .Q(
        npu_inst_pe_1_2_1_int_q_weight_1_), .QN(npu_inst_pe_1_2_1_n26) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_1_n112), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n8), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_1_n106), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n8), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_1_n111), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_1_n105), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_1_n110), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_1_n104), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_1_n109), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_1_n103), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_1_n108), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_1_n102), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_1_n107), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_1_n101), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_1_n86), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_1_n87), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n9), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_1_n88), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_1_n89), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_1_n90), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_1_n91), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_1_n92), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_1_n93), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_1_n94), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_1_n95), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_1_n96), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_1_n97), 
        .CK(npu_inst_pe_1_2_1_net4093), .RN(npu_inst_pe_1_2_1_n10), .Q(
        npu_inst_pe_1_2_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_1_net4087) );
  CLKGATETST_X1 npu_inst_pe_1_2_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n47), .SE(1'b0), .GCK(npu_inst_pe_1_2_1_net4093) );
  MUX2_X1 npu_inst_pe_1_2_2_U153 ( .A(npu_inst_pe_1_2_2_n31), .B(
        npu_inst_pe_1_2_2_n28), .S(npu_inst_pe_1_2_2_n7), .Z(
        npu_inst_pe_1_2_2_N93) );
  MUX2_X1 npu_inst_pe_1_2_2_U152 ( .A(npu_inst_pe_1_2_2_n30), .B(
        npu_inst_pe_1_2_2_n29), .S(npu_inst_pe_1_2_2_n5), .Z(
        npu_inst_pe_1_2_2_n31) );
  MUX2_X1 npu_inst_pe_1_2_2_U151 ( .A(npu_inst_pe_1_2_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_2_n3), .Z(
        npu_inst_pe_1_2_2_n30) );
  MUX2_X1 npu_inst_pe_1_2_2_U150 ( .A(npu_inst_pe_1_2_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_2_n3), .Z(
        npu_inst_pe_1_2_2_n29) );
  MUX2_X1 npu_inst_pe_1_2_2_U149 ( .A(npu_inst_pe_1_2_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_2_n3), .Z(
        npu_inst_pe_1_2_2_n28) );
  MUX2_X1 npu_inst_pe_1_2_2_U148 ( .A(npu_inst_pe_1_2_2_n25), .B(
        npu_inst_pe_1_2_2_n22), .S(npu_inst_pe_1_2_2_n7), .Z(
        npu_inst_pe_1_2_2_N94) );
  MUX2_X1 npu_inst_pe_1_2_2_U147 ( .A(npu_inst_pe_1_2_2_n24), .B(
        npu_inst_pe_1_2_2_n23), .S(npu_inst_pe_1_2_2_n5), .Z(
        npu_inst_pe_1_2_2_n25) );
  MUX2_X1 npu_inst_pe_1_2_2_U146 ( .A(npu_inst_pe_1_2_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_2_n3), .Z(
        npu_inst_pe_1_2_2_n24) );
  MUX2_X1 npu_inst_pe_1_2_2_U145 ( .A(npu_inst_pe_1_2_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_2_n3), .Z(
        npu_inst_pe_1_2_2_n23) );
  MUX2_X1 npu_inst_pe_1_2_2_U144 ( .A(npu_inst_pe_1_2_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_2_n3), .Z(
        npu_inst_pe_1_2_2_n22) );
  MUX2_X1 npu_inst_pe_1_2_2_U143 ( .A(npu_inst_pe_1_2_2_n21), .B(
        npu_inst_pe_1_2_2_n18), .S(npu_inst_pe_1_2_2_n7), .Z(
        npu_inst_int_data_x_2__2__1_) );
  MUX2_X1 npu_inst_pe_1_2_2_U142 ( .A(npu_inst_pe_1_2_2_n20), .B(
        npu_inst_pe_1_2_2_n19), .S(npu_inst_pe_1_2_2_n5), .Z(
        npu_inst_pe_1_2_2_n21) );
  MUX2_X1 npu_inst_pe_1_2_2_U141 ( .A(npu_inst_pe_1_2_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_2_n3), .Z(
        npu_inst_pe_1_2_2_n20) );
  MUX2_X1 npu_inst_pe_1_2_2_U140 ( .A(npu_inst_pe_1_2_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_2_n3), .Z(
        npu_inst_pe_1_2_2_n19) );
  MUX2_X1 npu_inst_pe_1_2_2_U139 ( .A(npu_inst_pe_1_2_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_2_n3), .Z(
        npu_inst_pe_1_2_2_n18) );
  MUX2_X1 npu_inst_pe_1_2_2_U138 ( .A(npu_inst_pe_1_2_2_n17), .B(
        npu_inst_pe_1_2_2_n14), .S(npu_inst_pe_1_2_2_n7), .Z(
        npu_inst_int_data_x_2__2__0_) );
  MUX2_X1 npu_inst_pe_1_2_2_U137 ( .A(npu_inst_pe_1_2_2_n16), .B(
        npu_inst_pe_1_2_2_n15), .S(npu_inst_pe_1_2_2_n5), .Z(
        npu_inst_pe_1_2_2_n17) );
  MUX2_X1 npu_inst_pe_1_2_2_U136 ( .A(npu_inst_pe_1_2_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_2_n3), .Z(
        npu_inst_pe_1_2_2_n16) );
  MUX2_X1 npu_inst_pe_1_2_2_U135 ( .A(npu_inst_pe_1_2_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_2_n3), .Z(
        npu_inst_pe_1_2_2_n15) );
  MUX2_X1 npu_inst_pe_1_2_2_U134 ( .A(npu_inst_pe_1_2_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_2_n3), .Z(
        npu_inst_pe_1_2_2_n14) );
  XOR2_X1 npu_inst_pe_1_2_2_U133 ( .A(npu_inst_pe_1_2_2_int_data_0_), .B(
        npu_inst_int_data_res_2__2__0_), .Z(npu_inst_pe_1_2_2_N73) );
  AND2_X1 npu_inst_pe_1_2_2_U132 ( .A1(npu_inst_int_data_res_2__2__0_), .A2(
        npu_inst_pe_1_2_2_int_data_0_), .ZN(npu_inst_pe_1_2_2_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_2_U131 ( .A(npu_inst_int_data_res_2__2__0_), .B(
        npu_inst_pe_1_2_2_n12), .ZN(npu_inst_pe_1_2_2_N65) );
  OR2_X1 npu_inst_pe_1_2_2_U130 ( .A1(npu_inst_pe_1_2_2_n12), .A2(
        npu_inst_int_data_res_2__2__0_), .ZN(npu_inst_pe_1_2_2_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_2_U129 ( .A(npu_inst_int_data_res_2__2__2_), .B(
        npu_inst_pe_1_2_2_add_79_carry_2_), .Z(npu_inst_pe_1_2_2_N75) );
  AND2_X1 npu_inst_pe_1_2_2_U128 ( .A1(npu_inst_pe_1_2_2_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_2__2__2_), .ZN(
        npu_inst_pe_1_2_2_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_2_U127 ( .A(npu_inst_int_data_res_2__2__3_), .B(
        npu_inst_pe_1_2_2_add_79_carry_3_), .Z(npu_inst_pe_1_2_2_N76) );
  AND2_X1 npu_inst_pe_1_2_2_U126 ( .A1(npu_inst_pe_1_2_2_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_2__2__3_), .ZN(
        npu_inst_pe_1_2_2_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_2_U125 ( .A(npu_inst_int_data_res_2__2__4_), .B(
        npu_inst_pe_1_2_2_add_79_carry_4_), .Z(npu_inst_pe_1_2_2_N77) );
  AND2_X1 npu_inst_pe_1_2_2_U124 ( .A1(npu_inst_pe_1_2_2_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_2__2__4_), .ZN(
        npu_inst_pe_1_2_2_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_2_U123 ( .A(npu_inst_int_data_res_2__2__5_), .B(
        npu_inst_pe_1_2_2_add_79_carry_5_), .Z(npu_inst_pe_1_2_2_N78) );
  AND2_X1 npu_inst_pe_1_2_2_U122 ( .A1(npu_inst_pe_1_2_2_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_2__2__5_), .ZN(
        npu_inst_pe_1_2_2_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_2_U121 ( .A(npu_inst_int_data_res_2__2__6_), .B(
        npu_inst_pe_1_2_2_add_79_carry_6_), .Z(npu_inst_pe_1_2_2_N79) );
  AND2_X1 npu_inst_pe_1_2_2_U120 ( .A1(npu_inst_pe_1_2_2_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_2__2__6_), .ZN(
        npu_inst_pe_1_2_2_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_2_U119 ( .A(npu_inst_int_data_res_2__2__7_), .B(
        npu_inst_pe_1_2_2_add_79_carry_7_), .Z(npu_inst_pe_1_2_2_N80) );
  XNOR2_X1 npu_inst_pe_1_2_2_U118 ( .A(npu_inst_pe_1_2_2_sub_77_carry_2_), .B(
        npu_inst_int_data_res_2__2__2_), .ZN(npu_inst_pe_1_2_2_N67) );
  OR2_X1 npu_inst_pe_1_2_2_U117 ( .A1(npu_inst_int_data_res_2__2__2_), .A2(
        npu_inst_pe_1_2_2_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_2_2_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_2_U116 ( .A(npu_inst_pe_1_2_2_sub_77_carry_3_), .B(
        npu_inst_int_data_res_2__2__3_), .ZN(npu_inst_pe_1_2_2_N68) );
  OR2_X1 npu_inst_pe_1_2_2_U115 ( .A1(npu_inst_int_data_res_2__2__3_), .A2(
        npu_inst_pe_1_2_2_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_2_2_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_2_U114 ( .A(npu_inst_pe_1_2_2_sub_77_carry_4_), .B(
        npu_inst_int_data_res_2__2__4_), .ZN(npu_inst_pe_1_2_2_N69) );
  OR2_X1 npu_inst_pe_1_2_2_U113 ( .A1(npu_inst_int_data_res_2__2__4_), .A2(
        npu_inst_pe_1_2_2_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_2_2_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_2_U112 ( .A(npu_inst_pe_1_2_2_sub_77_carry_5_), .B(
        npu_inst_int_data_res_2__2__5_), .ZN(npu_inst_pe_1_2_2_N70) );
  OR2_X1 npu_inst_pe_1_2_2_U111 ( .A1(npu_inst_int_data_res_2__2__5_), .A2(
        npu_inst_pe_1_2_2_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_2_2_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_2_U110 ( .A(npu_inst_pe_1_2_2_sub_77_carry_6_), .B(
        npu_inst_int_data_res_2__2__6_), .ZN(npu_inst_pe_1_2_2_N71) );
  OR2_X1 npu_inst_pe_1_2_2_U109 ( .A1(npu_inst_int_data_res_2__2__6_), .A2(
        npu_inst_pe_1_2_2_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_2_2_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_2_U108 ( .A(npu_inst_int_data_res_2__2__7_), .B(
        npu_inst_pe_1_2_2_sub_77_carry_7_), .ZN(npu_inst_pe_1_2_2_N72) );
  INV_X1 npu_inst_pe_1_2_2_U107 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_2_2_n6)
         );
  INV_X1 npu_inst_pe_1_2_2_U106 ( .A(npu_inst_pe_1_2_2_n6), .ZN(
        npu_inst_pe_1_2_2_n5) );
  INV_X1 npu_inst_pe_1_2_2_U105 ( .A(npu_inst_n40), .ZN(npu_inst_pe_1_2_2_n2)
         );
  AOI22_X1 npu_inst_pe_1_2_2_U104 ( .A1(npu_inst_int_data_y_3__2__0_), .A2(
        npu_inst_pe_1_2_2_n58), .B1(npu_inst_pe_1_2_2_n118), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_2_n57) );
  INV_X1 npu_inst_pe_1_2_2_U103 ( .A(npu_inst_pe_1_2_2_n57), .ZN(
        npu_inst_pe_1_2_2_n107) );
  AOI22_X1 npu_inst_pe_1_2_2_U102 ( .A1(npu_inst_int_data_y_3__2__0_), .A2(
        npu_inst_pe_1_2_2_n54), .B1(npu_inst_pe_1_2_2_n117), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_2_n53) );
  INV_X1 npu_inst_pe_1_2_2_U99 ( .A(npu_inst_pe_1_2_2_n53), .ZN(
        npu_inst_pe_1_2_2_n108) );
  AOI22_X1 npu_inst_pe_1_2_2_U98 ( .A1(npu_inst_int_data_y_3__2__0_), .A2(
        npu_inst_pe_1_2_2_n50), .B1(npu_inst_pe_1_2_2_n116), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_2_n49) );
  INV_X1 npu_inst_pe_1_2_2_U97 ( .A(npu_inst_pe_1_2_2_n49), .ZN(
        npu_inst_pe_1_2_2_n109) );
  AOI22_X1 npu_inst_pe_1_2_2_U96 ( .A1(npu_inst_int_data_y_3__2__0_), .A2(
        npu_inst_pe_1_2_2_n46), .B1(npu_inst_pe_1_2_2_n115), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_2_n45) );
  INV_X1 npu_inst_pe_1_2_2_U95 ( .A(npu_inst_pe_1_2_2_n45), .ZN(
        npu_inst_pe_1_2_2_n110) );
  AOI22_X1 npu_inst_pe_1_2_2_U94 ( .A1(npu_inst_int_data_y_3__2__0_), .A2(
        npu_inst_pe_1_2_2_n42), .B1(npu_inst_pe_1_2_2_n114), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_2_n41) );
  INV_X1 npu_inst_pe_1_2_2_U93 ( .A(npu_inst_pe_1_2_2_n41), .ZN(
        npu_inst_pe_1_2_2_n111) );
  AOI22_X1 npu_inst_pe_1_2_2_U92 ( .A1(npu_inst_int_data_y_3__2__1_), .A2(
        npu_inst_pe_1_2_2_n58), .B1(npu_inst_pe_1_2_2_n118), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_2_n59) );
  INV_X1 npu_inst_pe_1_2_2_U91 ( .A(npu_inst_pe_1_2_2_n59), .ZN(
        npu_inst_pe_1_2_2_n101) );
  AOI22_X1 npu_inst_pe_1_2_2_U90 ( .A1(npu_inst_int_data_y_3__2__1_), .A2(
        npu_inst_pe_1_2_2_n54), .B1(npu_inst_pe_1_2_2_n117), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_2_n55) );
  INV_X1 npu_inst_pe_1_2_2_U89 ( .A(npu_inst_pe_1_2_2_n55), .ZN(
        npu_inst_pe_1_2_2_n102) );
  AOI22_X1 npu_inst_pe_1_2_2_U88 ( .A1(npu_inst_int_data_y_3__2__1_), .A2(
        npu_inst_pe_1_2_2_n50), .B1(npu_inst_pe_1_2_2_n116), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_2_n51) );
  INV_X1 npu_inst_pe_1_2_2_U87 ( .A(npu_inst_pe_1_2_2_n51), .ZN(
        npu_inst_pe_1_2_2_n103) );
  AOI22_X1 npu_inst_pe_1_2_2_U86 ( .A1(npu_inst_int_data_y_3__2__1_), .A2(
        npu_inst_pe_1_2_2_n46), .B1(npu_inst_pe_1_2_2_n115), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_2_n47) );
  INV_X1 npu_inst_pe_1_2_2_U85 ( .A(npu_inst_pe_1_2_2_n47), .ZN(
        npu_inst_pe_1_2_2_n104) );
  AOI22_X1 npu_inst_pe_1_2_2_U84 ( .A1(npu_inst_int_data_y_3__2__1_), .A2(
        npu_inst_pe_1_2_2_n42), .B1(npu_inst_pe_1_2_2_n114), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_2_n43) );
  INV_X1 npu_inst_pe_1_2_2_U83 ( .A(npu_inst_pe_1_2_2_n43), .ZN(
        npu_inst_pe_1_2_2_n105) );
  AOI22_X1 npu_inst_pe_1_2_2_U82 ( .A1(npu_inst_pe_1_2_2_n38), .A2(
        npu_inst_int_data_y_3__2__1_), .B1(npu_inst_pe_1_2_2_n113), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_2_n39) );
  INV_X1 npu_inst_pe_1_2_2_U81 ( .A(npu_inst_pe_1_2_2_n39), .ZN(
        npu_inst_pe_1_2_2_n106) );
  AND2_X1 npu_inst_pe_1_2_2_U80 ( .A1(npu_inst_pe_1_2_2_N93), .A2(npu_inst_n40), .ZN(npu_inst_int_data_y_2__2__0_) );
  NAND2_X1 npu_inst_pe_1_2_2_U79 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_2_n60), .ZN(npu_inst_pe_1_2_2_n74) );
  OAI21_X1 npu_inst_pe_1_2_2_U78 ( .B1(npu_inst_pe_1_2_2_n63), .B2(
        npu_inst_pe_1_2_2_n60), .A(npu_inst_pe_1_2_2_n74), .ZN(
        npu_inst_pe_1_2_2_n97) );
  NAND2_X1 npu_inst_pe_1_2_2_U77 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_2_n60), .ZN(npu_inst_pe_1_2_2_n73) );
  OAI21_X1 npu_inst_pe_1_2_2_U76 ( .B1(npu_inst_pe_1_2_2_n61), .B2(
        npu_inst_pe_1_2_2_n60), .A(npu_inst_pe_1_2_2_n73), .ZN(
        npu_inst_pe_1_2_2_n96) );
  NAND2_X1 npu_inst_pe_1_2_2_U75 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_2_n56), .ZN(npu_inst_pe_1_2_2_n72) );
  OAI21_X1 npu_inst_pe_1_2_2_U74 ( .B1(npu_inst_pe_1_2_2_n63), .B2(
        npu_inst_pe_1_2_2_n56), .A(npu_inst_pe_1_2_2_n72), .ZN(
        npu_inst_pe_1_2_2_n95) );
  NAND2_X1 npu_inst_pe_1_2_2_U73 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_2_n56), .ZN(npu_inst_pe_1_2_2_n71) );
  OAI21_X1 npu_inst_pe_1_2_2_U72 ( .B1(npu_inst_pe_1_2_2_n61), .B2(
        npu_inst_pe_1_2_2_n56), .A(npu_inst_pe_1_2_2_n71), .ZN(
        npu_inst_pe_1_2_2_n94) );
  NAND2_X1 npu_inst_pe_1_2_2_U71 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_2_n52), .ZN(npu_inst_pe_1_2_2_n70) );
  OAI21_X1 npu_inst_pe_1_2_2_U70 ( .B1(npu_inst_pe_1_2_2_n63), .B2(
        npu_inst_pe_1_2_2_n52), .A(npu_inst_pe_1_2_2_n70), .ZN(
        npu_inst_pe_1_2_2_n93) );
  NAND2_X1 npu_inst_pe_1_2_2_U69 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_2_n52), .ZN(npu_inst_pe_1_2_2_n69) );
  OAI21_X1 npu_inst_pe_1_2_2_U68 ( .B1(npu_inst_pe_1_2_2_n61), .B2(
        npu_inst_pe_1_2_2_n52), .A(npu_inst_pe_1_2_2_n69), .ZN(
        npu_inst_pe_1_2_2_n92) );
  NAND2_X1 npu_inst_pe_1_2_2_U67 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_2_n48), .ZN(npu_inst_pe_1_2_2_n68) );
  OAI21_X1 npu_inst_pe_1_2_2_U66 ( .B1(npu_inst_pe_1_2_2_n63), .B2(
        npu_inst_pe_1_2_2_n48), .A(npu_inst_pe_1_2_2_n68), .ZN(
        npu_inst_pe_1_2_2_n91) );
  NAND2_X1 npu_inst_pe_1_2_2_U65 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_2_n48), .ZN(npu_inst_pe_1_2_2_n67) );
  OAI21_X1 npu_inst_pe_1_2_2_U64 ( .B1(npu_inst_pe_1_2_2_n61), .B2(
        npu_inst_pe_1_2_2_n48), .A(npu_inst_pe_1_2_2_n67), .ZN(
        npu_inst_pe_1_2_2_n90) );
  NAND2_X1 npu_inst_pe_1_2_2_U63 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_2_n44), .ZN(npu_inst_pe_1_2_2_n66) );
  OAI21_X1 npu_inst_pe_1_2_2_U62 ( .B1(npu_inst_pe_1_2_2_n63), .B2(
        npu_inst_pe_1_2_2_n44), .A(npu_inst_pe_1_2_2_n66), .ZN(
        npu_inst_pe_1_2_2_n89) );
  NAND2_X1 npu_inst_pe_1_2_2_U61 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_2_n44), .ZN(npu_inst_pe_1_2_2_n65) );
  OAI21_X1 npu_inst_pe_1_2_2_U60 ( .B1(npu_inst_pe_1_2_2_n61), .B2(
        npu_inst_pe_1_2_2_n44), .A(npu_inst_pe_1_2_2_n65), .ZN(
        npu_inst_pe_1_2_2_n88) );
  NAND2_X1 npu_inst_pe_1_2_2_U59 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_2_n40), .ZN(npu_inst_pe_1_2_2_n64) );
  OAI21_X1 npu_inst_pe_1_2_2_U58 ( .B1(npu_inst_pe_1_2_2_n63), .B2(
        npu_inst_pe_1_2_2_n40), .A(npu_inst_pe_1_2_2_n64), .ZN(
        npu_inst_pe_1_2_2_n87) );
  NAND2_X1 npu_inst_pe_1_2_2_U57 ( .A1(npu_inst_pe_1_2_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_2_n40), .ZN(npu_inst_pe_1_2_2_n62) );
  OAI21_X1 npu_inst_pe_1_2_2_U56 ( .B1(npu_inst_pe_1_2_2_n61), .B2(
        npu_inst_pe_1_2_2_n40), .A(npu_inst_pe_1_2_2_n62), .ZN(
        npu_inst_pe_1_2_2_n86) );
  AOI22_X1 npu_inst_pe_1_2_2_U55 ( .A1(npu_inst_pe_1_2_2_n38), .A2(
        npu_inst_int_data_y_3__2__0_), .B1(npu_inst_pe_1_2_2_n113), .B2(
        npu_inst_pe_1_2_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_2_n37) );
  INV_X1 npu_inst_pe_1_2_2_U54 ( .A(npu_inst_pe_1_2_2_n37), .ZN(
        npu_inst_pe_1_2_2_n112) );
  AND2_X1 npu_inst_pe_1_2_2_U53 ( .A1(npu_inst_n40), .A2(npu_inst_pe_1_2_2_N94), .ZN(npu_inst_int_data_y_2__2__1_) );
  AOI222_X1 npu_inst_pe_1_2_2_U52 ( .A1(npu_inst_int_data_res_3__2__0_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N73), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N65), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n84) );
  INV_X1 npu_inst_pe_1_2_2_U51 ( .A(npu_inst_pe_1_2_2_n84), .ZN(
        npu_inst_pe_1_2_2_n100) );
  AOI222_X1 npu_inst_pe_1_2_2_U50 ( .A1(npu_inst_pe_1_2_2_n1), .A2(
        npu_inst_int_data_res_3__2__7_), .B1(npu_inst_pe_1_2_2_N80), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N72), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n75) );
  INV_X1 npu_inst_pe_1_2_2_U49 ( .A(npu_inst_pe_1_2_2_n75), .ZN(
        npu_inst_pe_1_2_2_n32) );
  AOI222_X1 npu_inst_pe_1_2_2_U48 ( .A1(npu_inst_int_data_res_3__2__1_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N74), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N66), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n83) );
  INV_X1 npu_inst_pe_1_2_2_U47 ( .A(npu_inst_pe_1_2_2_n83), .ZN(
        npu_inst_pe_1_2_2_n99) );
  AOI222_X1 npu_inst_pe_1_2_2_U46 ( .A1(npu_inst_int_data_res_3__2__3_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N76), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N68), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n81) );
  INV_X1 npu_inst_pe_1_2_2_U45 ( .A(npu_inst_pe_1_2_2_n81), .ZN(
        npu_inst_pe_1_2_2_n36) );
  AOI222_X1 npu_inst_pe_1_2_2_U44 ( .A1(npu_inst_int_data_res_3__2__4_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N77), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N69), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n80) );
  INV_X1 npu_inst_pe_1_2_2_U43 ( .A(npu_inst_pe_1_2_2_n80), .ZN(
        npu_inst_pe_1_2_2_n35) );
  AOI222_X1 npu_inst_pe_1_2_2_U42 ( .A1(npu_inst_int_data_res_3__2__5_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N78), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N70), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n79) );
  INV_X1 npu_inst_pe_1_2_2_U41 ( .A(npu_inst_pe_1_2_2_n79), .ZN(
        npu_inst_pe_1_2_2_n34) );
  AOI222_X1 npu_inst_pe_1_2_2_U40 ( .A1(npu_inst_int_data_res_3__2__6_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N79), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N71), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n78) );
  INV_X1 npu_inst_pe_1_2_2_U39 ( .A(npu_inst_pe_1_2_2_n78), .ZN(
        npu_inst_pe_1_2_2_n33) );
  AND2_X1 npu_inst_pe_1_2_2_U38 ( .A1(npu_inst_int_data_x_2__2__1_), .A2(
        npu_inst_pe_1_2_2_int_q_weight_1_), .ZN(npu_inst_pe_1_2_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_2_U37 ( .A1(npu_inst_int_data_x_2__2__0_), .A2(
        npu_inst_pe_1_2_2_int_q_weight_1_), .ZN(npu_inst_pe_1_2_2_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_2_2_U36 ( .A(npu_inst_pe_1_2_2_int_data_1_), .ZN(
        npu_inst_pe_1_2_2_n13) );
  NOR3_X1 npu_inst_pe_1_2_2_U35 ( .A1(npu_inst_pe_1_2_2_n26), .A2(npu_inst_n40), .A3(npu_inst_int_ckg[45]), .ZN(npu_inst_pe_1_2_2_n85) );
  OR2_X1 npu_inst_pe_1_2_2_U34 ( .A1(npu_inst_pe_1_2_2_n85), .A2(
        npu_inst_pe_1_2_2_n1), .ZN(npu_inst_pe_1_2_2_N84) );
  AOI222_X1 npu_inst_pe_1_2_2_U33 ( .A1(npu_inst_int_data_res_3__2__2_), .A2(
        npu_inst_pe_1_2_2_n1), .B1(npu_inst_pe_1_2_2_N75), .B2(
        npu_inst_pe_1_2_2_n76), .C1(npu_inst_pe_1_2_2_N67), .C2(
        npu_inst_pe_1_2_2_n77), .ZN(npu_inst_pe_1_2_2_n82) );
  INV_X1 npu_inst_pe_1_2_2_U32 ( .A(npu_inst_pe_1_2_2_n82), .ZN(
        npu_inst_pe_1_2_2_n98) );
  AOI22_X1 npu_inst_pe_1_2_2_U31 ( .A1(npu_inst_n40), .A2(
        npu_inst_int_data_y_3__2__1_), .B1(npu_inst_pe_1_2_2_n2), .B2(
        npu_inst_int_data_x_2__3__1_), .ZN(npu_inst_pe_1_2_2_n63) );
  AOI22_X1 npu_inst_pe_1_2_2_U30 ( .A1(npu_inst_n40), .A2(
        npu_inst_int_data_y_3__2__0_), .B1(npu_inst_pe_1_2_2_n2), .B2(
        npu_inst_int_data_x_2__3__0_), .ZN(npu_inst_pe_1_2_2_n61) );
  INV_X1 npu_inst_pe_1_2_2_U29 ( .A(npu_inst_pe_1_2_2_int_data_0_), .ZN(
        npu_inst_pe_1_2_2_n12) );
  INV_X1 npu_inst_pe_1_2_2_U28 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_2_2_n4)
         );
  OR3_X1 npu_inst_pe_1_2_2_U27 ( .A1(npu_inst_pe_1_2_2_n5), .A2(
        npu_inst_pe_1_2_2_n7), .A3(npu_inst_pe_1_2_2_n4), .ZN(
        npu_inst_pe_1_2_2_n56) );
  OR3_X1 npu_inst_pe_1_2_2_U26 ( .A1(npu_inst_pe_1_2_2_n4), .A2(
        npu_inst_pe_1_2_2_n7), .A3(npu_inst_pe_1_2_2_n6), .ZN(
        npu_inst_pe_1_2_2_n48) );
  INV_X1 npu_inst_pe_1_2_2_U25 ( .A(npu_inst_pe_1_2_2_n4), .ZN(
        npu_inst_pe_1_2_2_n3) );
  OR3_X1 npu_inst_pe_1_2_2_U24 ( .A1(npu_inst_pe_1_2_2_n3), .A2(
        npu_inst_pe_1_2_2_n7), .A3(npu_inst_pe_1_2_2_n6), .ZN(
        npu_inst_pe_1_2_2_n52) );
  OR3_X1 npu_inst_pe_1_2_2_U23 ( .A1(npu_inst_pe_1_2_2_n5), .A2(
        npu_inst_pe_1_2_2_n7), .A3(npu_inst_pe_1_2_2_n3), .ZN(
        npu_inst_pe_1_2_2_n60) );
  BUF_X1 npu_inst_pe_1_2_2_U22 ( .A(npu_inst_n26), .Z(npu_inst_pe_1_2_2_n1) );
  NOR2_X1 npu_inst_pe_1_2_2_U21 ( .A1(npu_inst_pe_1_2_2_n60), .A2(
        npu_inst_pe_1_2_2_n2), .ZN(npu_inst_pe_1_2_2_n58) );
  NOR2_X1 npu_inst_pe_1_2_2_U20 ( .A1(npu_inst_pe_1_2_2_n56), .A2(
        npu_inst_pe_1_2_2_n2), .ZN(npu_inst_pe_1_2_2_n54) );
  NOR2_X1 npu_inst_pe_1_2_2_U19 ( .A1(npu_inst_pe_1_2_2_n52), .A2(
        npu_inst_pe_1_2_2_n2), .ZN(npu_inst_pe_1_2_2_n50) );
  NOR2_X1 npu_inst_pe_1_2_2_U18 ( .A1(npu_inst_pe_1_2_2_n48), .A2(
        npu_inst_pe_1_2_2_n2), .ZN(npu_inst_pe_1_2_2_n46) );
  NOR2_X1 npu_inst_pe_1_2_2_U17 ( .A1(npu_inst_pe_1_2_2_n40), .A2(
        npu_inst_pe_1_2_2_n2), .ZN(npu_inst_pe_1_2_2_n38) );
  NOR2_X1 npu_inst_pe_1_2_2_U16 ( .A1(npu_inst_pe_1_2_2_n44), .A2(
        npu_inst_pe_1_2_2_n2), .ZN(npu_inst_pe_1_2_2_n42) );
  BUF_X1 npu_inst_pe_1_2_2_U15 ( .A(npu_inst_n85), .Z(npu_inst_pe_1_2_2_n7) );
  INV_X1 npu_inst_pe_1_2_2_U14 ( .A(npu_inst_n107), .ZN(npu_inst_pe_1_2_2_n11)
         );
  INV_X1 npu_inst_pe_1_2_2_U13 ( .A(npu_inst_pe_1_2_2_n38), .ZN(
        npu_inst_pe_1_2_2_n113) );
  INV_X1 npu_inst_pe_1_2_2_U12 ( .A(npu_inst_pe_1_2_2_n58), .ZN(
        npu_inst_pe_1_2_2_n118) );
  INV_X1 npu_inst_pe_1_2_2_U11 ( .A(npu_inst_pe_1_2_2_n54), .ZN(
        npu_inst_pe_1_2_2_n117) );
  INV_X1 npu_inst_pe_1_2_2_U10 ( .A(npu_inst_pe_1_2_2_n50), .ZN(
        npu_inst_pe_1_2_2_n116) );
  INV_X1 npu_inst_pe_1_2_2_U9 ( .A(npu_inst_pe_1_2_2_n46), .ZN(
        npu_inst_pe_1_2_2_n115) );
  INV_X1 npu_inst_pe_1_2_2_U8 ( .A(npu_inst_pe_1_2_2_n42), .ZN(
        npu_inst_pe_1_2_2_n114) );
  BUF_X1 npu_inst_pe_1_2_2_U7 ( .A(npu_inst_pe_1_2_2_n11), .Z(
        npu_inst_pe_1_2_2_n10) );
  BUF_X1 npu_inst_pe_1_2_2_U6 ( .A(npu_inst_pe_1_2_2_n11), .Z(
        npu_inst_pe_1_2_2_n9) );
  BUF_X1 npu_inst_pe_1_2_2_U5 ( .A(npu_inst_pe_1_2_2_n11), .Z(
        npu_inst_pe_1_2_2_n8) );
  NOR2_X1 npu_inst_pe_1_2_2_U4 ( .A1(npu_inst_pe_1_2_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_2_n1), .ZN(npu_inst_pe_1_2_2_n76) );
  NOR2_X1 npu_inst_pe_1_2_2_U3 ( .A1(npu_inst_pe_1_2_2_n27), .A2(
        npu_inst_pe_1_2_2_n1), .ZN(npu_inst_pe_1_2_2_n77) );
  FA_X1 npu_inst_pe_1_2_2_sub_77_U2_1 ( .A(npu_inst_int_data_res_2__2__1_), 
        .B(npu_inst_pe_1_2_2_n13), .CI(npu_inst_pe_1_2_2_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_2_2_sub_77_carry_2_), .S(npu_inst_pe_1_2_2_N66) );
  FA_X1 npu_inst_pe_1_2_2_add_79_U1_1 ( .A(npu_inst_int_data_res_2__2__1_), 
        .B(npu_inst_pe_1_2_2_int_data_1_), .CI(
        npu_inst_pe_1_2_2_add_79_carry_1_), .CO(
        npu_inst_pe_1_2_2_add_79_carry_2_), .S(npu_inst_pe_1_2_2_N74) );
  NAND3_X1 npu_inst_pe_1_2_2_U101 ( .A1(npu_inst_pe_1_2_2_n4), .A2(
        npu_inst_pe_1_2_2_n6), .A3(npu_inst_pe_1_2_2_n7), .ZN(
        npu_inst_pe_1_2_2_n44) );
  NAND3_X1 npu_inst_pe_1_2_2_U100 ( .A1(npu_inst_pe_1_2_2_n3), .A2(
        npu_inst_pe_1_2_2_n6), .A3(npu_inst_pe_1_2_2_n7), .ZN(
        npu_inst_pe_1_2_2_n40) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_2_n33), .CK(
        npu_inst_pe_1_2_2_net4064), .RN(npu_inst_pe_1_2_2_n8), .Q(
        npu_inst_int_data_res_2__2__6_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_2_n34), .CK(
        npu_inst_pe_1_2_2_net4064), .RN(npu_inst_pe_1_2_2_n8), .Q(
        npu_inst_int_data_res_2__2__5_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_2_n35), .CK(
        npu_inst_pe_1_2_2_net4064), .RN(npu_inst_pe_1_2_2_n8), .Q(
        npu_inst_int_data_res_2__2__4_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_2_n36), .CK(
        npu_inst_pe_1_2_2_net4064), .RN(npu_inst_pe_1_2_2_n8), .Q(
        npu_inst_int_data_res_2__2__3_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_2_n98), .CK(
        npu_inst_pe_1_2_2_net4064), .RN(npu_inst_pe_1_2_2_n8), .Q(
        npu_inst_int_data_res_2__2__2_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_2_n99), .CK(
        npu_inst_pe_1_2_2_net4064), .RN(npu_inst_pe_1_2_2_n8), .Q(
        npu_inst_int_data_res_2__2__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_2_n32), .CK(
        npu_inst_pe_1_2_2_net4064), .RN(npu_inst_pe_1_2_2_n8), .Q(
        npu_inst_int_data_res_2__2__7_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_2_n100), 
        .CK(npu_inst_pe_1_2_2_net4064), .RN(npu_inst_pe_1_2_2_n8), .Q(
        npu_inst_int_data_res_2__2__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_weight_reg_0_ ( .D(npu_inst_n93), .CK(
        npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n8), .Q(
        npu_inst_pe_1_2_2_int_q_weight_0_), .QN(npu_inst_pe_1_2_2_n27) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_weight_reg_1_ ( .D(npu_inst_n99), .CK(
        npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n8), .Q(
        npu_inst_pe_1_2_2_int_q_weight_1_), .QN(npu_inst_pe_1_2_2_n26) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_2_n112), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n8), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_2_n106), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n8), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_2_n111), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_2_n105), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_2_n110), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_2_n104), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_2_n109), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_2_n103), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_2_n108), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_2_n102), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_2_n107), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_2_n101), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_2_n86), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_2_n87), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n9), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_2_n88), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_2_n89), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_2_n90), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_2_n91), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_2_n92), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_2_n93), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_2_n94), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_2_n95), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_2_n96), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_2_n97), 
        .CK(npu_inst_pe_1_2_2_net4070), .RN(npu_inst_pe_1_2_2_n10), .Q(
        npu_inst_pe_1_2_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_2_net4064) );
  CLKGATETST_X1 npu_inst_pe_1_2_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n47), .SE(1'b0), .GCK(npu_inst_pe_1_2_2_net4070) );
  MUX2_X1 npu_inst_pe_1_2_3_U153 ( .A(npu_inst_pe_1_2_3_n31), .B(
        npu_inst_pe_1_2_3_n28), .S(npu_inst_pe_1_2_3_n7), .Z(
        npu_inst_pe_1_2_3_N93) );
  MUX2_X1 npu_inst_pe_1_2_3_U152 ( .A(npu_inst_pe_1_2_3_n30), .B(
        npu_inst_pe_1_2_3_n29), .S(npu_inst_pe_1_2_3_n5), .Z(
        npu_inst_pe_1_2_3_n31) );
  MUX2_X1 npu_inst_pe_1_2_3_U151 ( .A(npu_inst_pe_1_2_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_3_n3), .Z(
        npu_inst_pe_1_2_3_n30) );
  MUX2_X1 npu_inst_pe_1_2_3_U150 ( .A(npu_inst_pe_1_2_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_3_n3), .Z(
        npu_inst_pe_1_2_3_n29) );
  MUX2_X1 npu_inst_pe_1_2_3_U149 ( .A(npu_inst_pe_1_2_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_3_n3), .Z(
        npu_inst_pe_1_2_3_n28) );
  MUX2_X1 npu_inst_pe_1_2_3_U148 ( .A(npu_inst_pe_1_2_3_n25), .B(
        npu_inst_pe_1_2_3_n22), .S(npu_inst_pe_1_2_3_n7), .Z(
        npu_inst_pe_1_2_3_N94) );
  MUX2_X1 npu_inst_pe_1_2_3_U147 ( .A(npu_inst_pe_1_2_3_n24), .B(
        npu_inst_pe_1_2_3_n23), .S(npu_inst_pe_1_2_3_n5), .Z(
        npu_inst_pe_1_2_3_n25) );
  MUX2_X1 npu_inst_pe_1_2_3_U146 ( .A(npu_inst_pe_1_2_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_3_n3), .Z(
        npu_inst_pe_1_2_3_n24) );
  MUX2_X1 npu_inst_pe_1_2_3_U145 ( .A(npu_inst_pe_1_2_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_3_n3), .Z(
        npu_inst_pe_1_2_3_n23) );
  MUX2_X1 npu_inst_pe_1_2_3_U144 ( .A(npu_inst_pe_1_2_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_3_n3), .Z(
        npu_inst_pe_1_2_3_n22) );
  MUX2_X1 npu_inst_pe_1_2_3_U143 ( .A(npu_inst_pe_1_2_3_n21), .B(
        npu_inst_pe_1_2_3_n18), .S(npu_inst_pe_1_2_3_n7), .Z(
        npu_inst_int_data_x_2__3__1_) );
  MUX2_X1 npu_inst_pe_1_2_3_U142 ( .A(npu_inst_pe_1_2_3_n20), .B(
        npu_inst_pe_1_2_3_n19), .S(npu_inst_pe_1_2_3_n5), .Z(
        npu_inst_pe_1_2_3_n21) );
  MUX2_X1 npu_inst_pe_1_2_3_U141 ( .A(npu_inst_pe_1_2_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_3_n3), .Z(
        npu_inst_pe_1_2_3_n20) );
  MUX2_X1 npu_inst_pe_1_2_3_U140 ( .A(npu_inst_pe_1_2_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_3_n3), .Z(
        npu_inst_pe_1_2_3_n19) );
  MUX2_X1 npu_inst_pe_1_2_3_U139 ( .A(npu_inst_pe_1_2_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_3_n3), .Z(
        npu_inst_pe_1_2_3_n18) );
  MUX2_X1 npu_inst_pe_1_2_3_U138 ( .A(npu_inst_pe_1_2_3_n17), .B(
        npu_inst_pe_1_2_3_n14), .S(npu_inst_pe_1_2_3_n7), .Z(
        npu_inst_int_data_x_2__3__0_) );
  MUX2_X1 npu_inst_pe_1_2_3_U137 ( .A(npu_inst_pe_1_2_3_n16), .B(
        npu_inst_pe_1_2_3_n15), .S(npu_inst_pe_1_2_3_n5), .Z(
        npu_inst_pe_1_2_3_n17) );
  MUX2_X1 npu_inst_pe_1_2_3_U136 ( .A(npu_inst_pe_1_2_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_3_n3), .Z(
        npu_inst_pe_1_2_3_n16) );
  MUX2_X1 npu_inst_pe_1_2_3_U135 ( .A(npu_inst_pe_1_2_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_3_n3), .Z(
        npu_inst_pe_1_2_3_n15) );
  MUX2_X1 npu_inst_pe_1_2_3_U134 ( .A(npu_inst_pe_1_2_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_3_n3), .Z(
        npu_inst_pe_1_2_3_n14) );
  XOR2_X1 npu_inst_pe_1_2_3_U133 ( .A(npu_inst_pe_1_2_3_int_data_0_), .B(
        npu_inst_int_data_res_2__3__0_), .Z(npu_inst_pe_1_2_3_N73) );
  AND2_X1 npu_inst_pe_1_2_3_U132 ( .A1(npu_inst_int_data_res_2__3__0_), .A2(
        npu_inst_pe_1_2_3_int_data_0_), .ZN(npu_inst_pe_1_2_3_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_3_U131 ( .A(npu_inst_int_data_res_2__3__0_), .B(
        npu_inst_pe_1_2_3_n12), .ZN(npu_inst_pe_1_2_3_N65) );
  OR2_X1 npu_inst_pe_1_2_3_U130 ( .A1(npu_inst_pe_1_2_3_n12), .A2(
        npu_inst_int_data_res_2__3__0_), .ZN(npu_inst_pe_1_2_3_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_3_U129 ( .A(npu_inst_int_data_res_2__3__2_), .B(
        npu_inst_pe_1_2_3_add_79_carry_2_), .Z(npu_inst_pe_1_2_3_N75) );
  AND2_X1 npu_inst_pe_1_2_3_U128 ( .A1(npu_inst_pe_1_2_3_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_2__3__2_), .ZN(
        npu_inst_pe_1_2_3_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_3_U127 ( .A(npu_inst_int_data_res_2__3__3_), .B(
        npu_inst_pe_1_2_3_add_79_carry_3_), .Z(npu_inst_pe_1_2_3_N76) );
  AND2_X1 npu_inst_pe_1_2_3_U126 ( .A1(npu_inst_pe_1_2_3_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_2__3__3_), .ZN(
        npu_inst_pe_1_2_3_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_3_U125 ( .A(npu_inst_int_data_res_2__3__4_), .B(
        npu_inst_pe_1_2_3_add_79_carry_4_), .Z(npu_inst_pe_1_2_3_N77) );
  AND2_X1 npu_inst_pe_1_2_3_U124 ( .A1(npu_inst_pe_1_2_3_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_2__3__4_), .ZN(
        npu_inst_pe_1_2_3_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_3_U123 ( .A(npu_inst_int_data_res_2__3__5_), .B(
        npu_inst_pe_1_2_3_add_79_carry_5_), .Z(npu_inst_pe_1_2_3_N78) );
  AND2_X1 npu_inst_pe_1_2_3_U122 ( .A1(npu_inst_pe_1_2_3_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_2__3__5_), .ZN(
        npu_inst_pe_1_2_3_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_3_U121 ( .A(npu_inst_int_data_res_2__3__6_), .B(
        npu_inst_pe_1_2_3_add_79_carry_6_), .Z(npu_inst_pe_1_2_3_N79) );
  AND2_X1 npu_inst_pe_1_2_3_U120 ( .A1(npu_inst_pe_1_2_3_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_2__3__6_), .ZN(
        npu_inst_pe_1_2_3_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_3_U119 ( .A(npu_inst_int_data_res_2__3__7_), .B(
        npu_inst_pe_1_2_3_add_79_carry_7_), .Z(npu_inst_pe_1_2_3_N80) );
  XNOR2_X1 npu_inst_pe_1_2_3_U118 ( .A(npu_inst_pe_1_2_3_sub_77_carry_2_), .B(
        npu_inst_int_data_res_2__3__2_), .ZN(npu_inst_pe_1_2_3_N67) );
  OR2_X1 npu_inst_pe_1_2_3_U117 ( .A1(npu_inst_int_data_res_2__3__2_), .A2(
        npu_inst_pe_1_2_3_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_2_3_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_3_U116 ( .A(npu_inst_pe_1_2_3_sub_77_carry_3_), .B(
        npu_inst_int_data_res_2__3__3_), .ZN(npu_inst_pe_1_2_3_N68) );
  OR2_X1 npu_inst_pe_1_2_3_U115 ( .A1(npu_inst_int_data_res_2__3__3_), .A2(
        npu_inst_pe_1_2_3_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_2_3_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_3_U114 ( .A(npu_inst_pe_1_2_3_sub_77_carry_4_), .B(
        npu_inst_int_data_res_2__3__4_), .ZN(npu_inst_pe_1_2_3_N69) );
  OR2_X1 npu_inst_pe_1_2_3_U113 ( .A1(npu_inst_int_data_res_2__3__4_), .A2(
        npu_inst_pe_1_2_3_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_2_3_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_3_U112 ( .A(npu_inst_pe_1_2_3_sub_77_carry_5_), .B(
        npu_inst_int_data_res_2__3__5_), .ZN(npu_inst_pe_1_2_3_N70) );
  OR2_X1 npu_inst_pe_1_2_3_U111 ( .A1(npu_inst_int_data_res_2__3__5_), .A2(
        npu_inst_pe_1_2_3_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_2_3_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_3_U110 ( .A(npu_inst_pe_1_2_3_sub_77_carry_6_), .B(
        npu_inst_int_data_res_2__3__6_), .ZN(npu_inst_pe_1_2_3_N71) );
  OR2_X1 npu_inst_pe_1_2_3_U109 ( .A1(npu_inst_int_data_res_2__3__6_), .A2(
        npu_inst_pe_1_2_3_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_2_3_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_3_U108 ( .A(npu_inst_int_data_res_2__3__7_), .B(
        npu_inst_pe_1_2_3_sub_77_carry_7_), .ZN(npu_inst_pe_1_2_3_N72) );
  INV_X1 npu_inst_pe_1_2_3_U107 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_2_3_n6)
         );
  INV_X1 npu_inst_pe_1_2_3_U106 ( .A(npu_inst_pe_1_2_3_n6), .ZN(
        npu_inst_pe_1_2_3_n5) );
  INV_X1 npu_inst_pe_1_2_3_U105 ( .A(npu_inst_n40), .ZN(npu_inst_pe_1_2_3_n2)
         );
  AOI22_X1 npu_inst_pe_1_2_3_U104 ( .A1(npu_inst_int_data_y_3__3__0_), .A2(
        npu_inst_pe_1_2_3_n58), .B1(npu_inst_pe_1_2_3_n118), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_3_n57) );
  INV_X1 npu_inst_pe_1_2_3_U103 ( .A(npu_inst_pe_1_2_3_n57), .ZN(
        npu_inst_pe_1_2_3_n107) );
  AOI22_X1 npu_inst_pe_1_2_3_U102 ( .A1(npu_inst_int_data_y_3__3__0_), .A2(
        npu_inst_pe_1_2_3_n54), .B1(npu_inst_pe_1_2_3_n117), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_3_n53) );
  INV_X1 npu_inst_pe_1_2_3_U99 ( .A(npu_inst_pe_1_2_3_n53), .ZN(
        npu_inst_pe_1_2_3_n108) );
  AOI22_X1 npu_inst_pe_1_2_3_U98 ( .A1(npu_inst_int_data_y_3__3__0_), .A2(
        npu_inst_pe_1_2_3_n50), .B1(npu_inst_pe_1_2_3_n116), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_3_n49) );
  INV_X1 npu_inst_pe_1_2_3_U97 ( .A(npu_inst_pe_1_2_3_n49), .ZN(
        npu_inst_pe_1_2_3_n109) );
  AOI22_X1 npu_inst_pe_1_2_3_U96 ( .A1(npu_inst_int_data_y_3__3__0_), .A2(
        npu_inst_pe_1_2_3_n46), .B1(npu_inst_pe_1_2_3_n115), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_3_n45) );
  INV_X1 npu_inst_pe_1_2_3_U95 ( .A(npu_inst_pe_1_2_3_n45), .ZN(
        npu_inst_pe_1_2_3_n110) );
  AOI22_X1 npu_inst_pe_1_2_3_U94 ( .A1(npu_inst_int_data_y_3__3__0_), .A2(
        npu_inst_pe_1_2_3_n42), .B1(npu_inst_pe_1_2_3_n114), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_3_n41) );
  INV_X1 npu_inst_pe_1_2_3_U93 ( .A(npu_inst_pe_1_2_3_n41), .ZN(
        npu_inst_pe_1_2_3_n111) );
  AOI22_X1 npu_inst_pe_1_2_3_U92 ( .A1(npu_inst_int_data_y_3__3__1_), .A2(
        npu_inst_pe_1_2_3_n58), .B1(npu_inst_pe_1_2_3_n118), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_3_n59) );
  INV_X1 npu_inst_pe_1_2_3_U91 ( .A(npu_inst_pe_1_2_3_n59), .ZN(
        npu_inst_pe_1_2_3_n101) );
  AOI22_X1 npu_inst_pe_1_2_3_U90 ( .A1(npu_inst_int_data_y_3__3__1_), .A2(
        npu_inst_pe_1_2_3_n54), .B1(npu_inst_pe_1_2_3_n117), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_3_n55) );
  INV_X1 npu_inst_pe_1_2_3_U89 ( .A(npu_inst_pe_1_2_3_n55), .ZN(
        npu_inst_pe_1_2_3_n102) );
  AOI22_X1 npu_inst_pe_1_2_3_U88 ( .A1(npu_inst_int_data_y_3__3__1_), .A2(
        npu_inst_pe_1_2_3_n50), .B1(npu_inst_pe_1_2_3_n116), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_3_n51) );
  INV_X1 npu_inst_pe_1_2_3_U87 ( .A(npu_inst_pe_1_2_3_n51), .ZN(
        npu_inst_pe_1_2_3_n103) );
  AOI22_X1 npu_inst_pe_1_2_3_U86 ( .A1(npu_inst_int_data_y_3__3__1_), .A2(
        npu_inst_pe_1_2_3_n46), .B1(npu_inst_pe_1_2_3_n115), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_3_n47) );
  INV_X1 npu_inst_pe_1_2_3_U85 ( .A(npu_inst_pe_1_2_3_n47), .ZN(
        npu_inst_pe_1_2_3_n104) );
  AOI22_X1 npu_inst_pe_1_2_3_U84 ( .A1(npu_inst_int_data_y_3__3__1_), .A2(
        npu_inst_pe_1_2_3_n42), .B1(npu_inst_pe_1_2_3_n114), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_3_n43) );
  INV_X1 npu_inst_pe_1_2_3_U83 ( .A(npu_inst_pe_1_2_3_n43), .ZN(
        npu_inst_pe_1_2_3_n105) );
  AOI22_X1 npu_inst_pe_1_2_3_U82 ( .A1(npu_inst_pe_1_2_3_n38), .A2(
        npu_inst_int_data_y_3__3__1_), .B1(npu_inst_pe_1_2_3_n113), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_3_n39) );
  INV_X1 npu_inst_pe_1_2_3_U81 ( .A(npu_inst_pe_1_2_3_n39), .ZN(
        npu_inst_pe_1_2_3_n106) );
  AND2_X1 npu_inst_pe_1_2_3_U80 ( .A1(npu_inst_pe_1_2_3_N93), .A2(npu_inst_n40), .ZN(npu_inst_int_data_y_2__3__0_) );
  NAND2_X1 npu_inst_pe_1_2_3_U79 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_3_n60), .ZN(npu_inst_pe_1_2_3_n74) );
  OAI21_X1 npu_inst_pe_1_2_3_U78 ( .B1(npu_inst_pe_1_2_3_n63), .B2(
        npu_inst_pe_1_2_3_n60), .A(npu_inst_pe_1_2_3_n74), .ZN(
        npu_inst_pe_1_2_3_n97) );
  NAND2_X1 npu_inst_pe_1_2_3_U77 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_3_n60), .ZN(npu_inst_pe_1_2_3_n73) );
  OAI21_X1 npu_inst_pe_1_2_3_U76 ( .B1(npu_inst_pe_1_2_3_n61), .B2(
        npu_inst_pe_1_2_3_n60), .A(npu_inst_pe_1_2_3_n73), .ZN(
        npu_inst_pe_1_2_3_n96) );
  NAND2_X1 npu_inst_pe_1_2_3_U75 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_3_n56), .ZN(npu_inst_pe_1_2_3_n72) );
  OAI21_X1 npu_inst_pe_1_2_3_U74 ( .B1(npu_inst_pe_1_2_3_n63), .B2(
        npu_inst_pe_1_2_3_n56), .A(npu_inst_pe_1_2_3_n72), .ZN(
        npu_inst_pe_1_2_3_n95) );
  NAND2_X1 npu_inst_pe_1_2_3_U73 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_3_n56), .ZN(npu_inst_pe_1_2_3_n71) );
  OAI21_X1 npu_inst_pe_1_2_3_U72 ( .B1(npu_inst_pe_1_2_3_n61), .B2(
        npu_inst_pe_1_2_3_n56), .A(npu_inst_pe_1_2_3_n71), .ZN(
        npu_inst_pe_1_2_3_n94) );
  NAND2_X1 npu_inst_pe_1_2_3_U71 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_3_n52), .ZN(npu_inst_pe_1_2_3_n70) );
  OAI21_X1 npu_inst_pe_1_2_3_U70 ( .B1(npu_inst_pe_1_2_3_n63), .B2(
        npu_inst_pe_1_2_3_n52), .A(npu_inst_pe_1_2_3_n70), .ZN(
        npu_inst_pe_1_2_3_n93) );
  NAND2_X1 npu_inst_pe_1_2_3_U69 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_3_n52), .ZN(npu_inst_pe_1_2_3_n69) );
  OAI21_X1 npu_inst_pe_1_2_3_U68 ( .B1(npu_inst_pe_1_2_3_n61), .B2(
        npu_inst_pe_1_2_3_n52), .A(npu_inst_pe_1_2_3_n69), .ZN(
        npu_inst_pe_1_2_3_n92) );
  NAND2_X1 npu_inst_pe_1_2_3_U67 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_3_n48), .ZN(npu_inst_pe_1_2_3_n68) );
  OAI21_X1 npu_inst_pe_1_2_3_U66 ( .B1(npu_inst_pe_1_2_3_n63), .B2(
        npu_inst_pe_1_2_3_n48), .A(npu_inst_pe_1_2_3_n68), .ZN(
        npu_inst_pe_1_2_3_n91) );
  NAND2_X1 npu_inst_pe_1_2_3_U65 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_3_n48), .ZN(npu_inst_pe_1_2_3_n67) );
  OAI21_X1 npu_inst_pe_1_2_3_U64 ( .B1(npu_inst_pe_1_2_3_n61), .B2(
        npu_inst_pe_1_2_3_n48), .A(npu_inst_pe_1_2_3_n67), .ZN(
        npu_inst_pe_1_2_3_n90) );
  NAND2_X1 npu_inst_pe_1_2_3_U63 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_3_n44), .ZN(npu_inst_pe_1_2_3_n66) );
  OAI21_X1 npu_inst_pe_1_2_3_U62 ( .B1(npu_inst_pe_1_2_3_n63), .B2(
        npu_inst_pe_1_2_3_n44), .A(npu_inst_pe_1_2_3_n66), .ZN(
        npu_inst_pe_1_2_3_n89) );
  NAND2_X1 npu_inst_pe_1_2_3_U61 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_3_n44), .ZN(npu_inst_pe_1_2_3_n65) );
  OAI21_X1 npu_inst_pe_1_2_3_U60 ( .B1(npu_inst_pe_1_2_3_n61), .B2(
        npu_inst_pe_1_2_3_n44), .A(npu_inst_pe_1_2_3_n65), .ZN(
        npu_inst_pe_1_2_3_n88) );
  NAND2_X1 npu_inst_pe_1_2_3_U59 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_3_n40), .ZN(npu_inst_pe_1_2_3_n64) );
  OAI21_X1 npu_inst_pe_1_2_3_U58 ( .B1(npu_inst_pe_1_2_3_n63), .B2(
        npu_inst_pe_1_2_3_n40), .A(npu_inst_pe_1_2_3_n64), .ZN(
        npu_inst_pe_1_2_3_n87) );
  NAND2_X1 npu_inst_pe_1_2_3_U57 ( .A1(npu_inst_pe_1_2_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_3_n40), .ZN(npu_inst_pe_1_2_3_n62) );
  OAI21_X1 npu_inst_pe_1_2_3_U56 ( .B1(npu_inst_pe_1_2_3_n61), .B2(
        npu_inst_pe_1_2_3_n40), .A(npu_inst_pe_1_2_3_n62), .ZN(
        npu_inst_pe_1_2_3_n86) );
  AOI22_X1 npu_inst_pe_1_2_3_U55 ( .A1(npu_inst_pe_1_2_3_n38), .A2(
        npu_inst_int_data_y_3__3__0_), .B1(npu_inst_pe_1_2_3_n113), .B2(
        npu_inst_pe_1_2_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_3_n37) );
  INV_X1 npu_inst_pe_1_2_3_U54 ( .A(npu_inst_pe_1_2_3_n37), .ZN(
        npu_inst_pe_1_2_3_n112) );
  AND2_X1 npu_inst_pe_1_2_3_U53 ( .A1(npu_inst_n40), .A2(npu_inst_pe_1_2_3_N94), .ZN(npu_inst_int_data_y_2__3__1_) );
  AOI222_X1 npu_inst_pe_1_2_3_U52 ( .A1(npu_inst_int_data_res_3__3__0_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N73), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N65), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n84) );
  INV_X1 npu_inst_pe_1_2_3_U51 ( .A(npu_inst_pe_1_2_3_n84), .ZN(
        npu_inst_pe_1_2_3_n100) );
  AOI222_X1 npu_inst_pe_1_2_3_U50 ( .A1(npu_inst_pe_1_2_3_n1), .A2(
        npu_inst_int_data_res_3__3__7_), .B1(npu_inst_pe_1_2_3_N80), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N72), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n75) );
  INV_X1 npu_inst_pe_1_2_3_U49 ( .A(npu_inst_pe_1_2_3_n75), .ZN(
        npu_inst_pe_1_2_3_n32) );
  AOI222_X1 npu_inst_pe_1_2_3_U48 ( .A1(npu_inst_int_data_res_3__3__1_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N74), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N66), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n83) );
  INV_X1 npu_inst_pe_1_2_3_U47 ( .A(npu_inst_pe_1_2_3_n83), .ZN(
        npu_inst_pe_1_2_3_n99) );
  AOI222_X1 npu_inst_pe_1_2_3_U46 ( .A1(npu_inst_int_data_res_3__3__3_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N76), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N68), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n81) );
  INV_X1 npu_inst_pe_1_2_3_U45 ( .A(npu_inst_pe_1_2_3_n81), .ZN(
        npu_inst_pe_1_2_3_n36) );
  AOI222_X1 npu_inst_pe_1_2_3_U44 ( .A1(npu_inst_int_data_res_3__3__4_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N77), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N69), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n80) );
  INV_X1 npu_inst_pe_1_2_3_U43 ( .A(npu_inst_pe_1_2_3_n80), .ZN(
        npu_inst_pe_1_2_3_n35) );
  AOI222_X1 npu_inst_pe_1_2_3_U42 ( .A1(npu_inst_int_data_res_3__3__5_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N78), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N70), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n79) );
  INV_X1 npu_inst_pe_1_2_3_U41 ( .A(npu_inst_pe_1_2_3_n79), .ZN(
        npu_inst_pe_1_2_3_n34) );
  AOI222_X1 npu_inst_pe_1_2_3_U40 ( .A1(npu_inst_int_data_res_3__3__6_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N79), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N71), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n78) );
  INV_X1 npu_inst_pe_1_2_3_U39 ( .A(npu_inst_pe_1_2_3_n78), .ZN(
        npu_inst_pe_1_2_3_n33) );
  AND2_X1 npu_inst_pe_1_2_3_U38 ( .A1(npu_inst_int_data_x_2__3__1_), .A2(
        npu_inst_pe_1_2_3_int_q_weight_1_), .ZN(npu_inst_pe_1_2_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_3_U37 ( .A1(npu_inst_int_data_x_2__3__0_), .A2(
        npu_inst_pe_1_2_3_int_q_weight_1_), .ZN(npu_inst_pe_1_2_3_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_2_3_U36 ( .A(npu_inst_pe_1_2_3_int_data_1_), .ZN(
        npu_inst_pe_1_2_3_n13) );
  NOR3_X1 npu_inst_pe_1_2_3_U35 ( .A1(npu_inst_pe_1_2_3_n26), .A2(npu_inst_n40), .A3(npu_inst_int_ckg[44]), .ZN(npu_inst_pe_1_2_3_n85) );
  OR2_X1 npu_inst_pe_1_2_3_U34 ( .A1(npu_inst_pe_1_2_3_n85), .A2(
        npu_inst_pe_1_2_3_n1), .ZN(npu_inst_pe_1_2_3_N84) );
  AOI222_X1 npu_inst_pe_1_2_3_U33 ( .A1(npu_inst_int_data_res_3__3__2_), .A2(
        npu_inst_pe_1_2_3_n1), .B1(npu_inst_pe_1_2_3_N75), .B2(
        npu_inst_pe_1_2_3_n76), .C1(npu_inst_pe_1_2_3_N67), .C2(
        npu_inst_pe_1_2_3_n77), .ZN(npu_inst_pe_1_2_3_n82) );
  INV_X1 npu_inst_pe_1_2_3_U32 ( .A(npu_inst_pe_1_2_3_n82), .ZN(
        npu_inst_pe_1_2_3_n98) );
  AOI22_X1 npu_inst_pe_1_2_3_U31 ( .A1(npu_inst_n40), .A2(
        npu_inst_int_data_y_3__3__1_), .B1(npu_inst_pe_1_2_3_n2), .B2(
        npu_inst_int_data_x_2__4__1_), .ZN(npu_inst_pe_1_2_3_n63) );
  AOI22_X1 npu_inst_pe_1_2_3_U30 ( .A1(npu_inst_n40), .A2(
        npu_inst_int_data_y_3__3__0_), .B1(npu_inst_pe_1_2_3_n2), .B2(
        npu_inst_int_data_x_2__4__0_), .ZN(npu_inst_pe_1_2_3_n61) );
  INV_X1 npu_inst_pe_1_2_3_U29 ( .A(npu_inst_pe_1_2_3_int_data_0_), .ZN(
        npu_inst_pe_1_2_3_n12) );
  INV_X1 npu_inst_pe_1_2_3_U28 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_2_3_n4)
         );
  OR3_X1 npu_inst_pe_1_2_3_U27 ( .A1(npu_inst_pe_1_2_3_n5), .A2(
        npu_inst_pe_1_2_3_n7), .A3(npu_inst_pe_1_2_3_n4), .ZN(
        npu_inst_pe_1_2_3_n56) );
  OR3_X1 npu_inst_pe_1_2_3_U26 ( .A1(npu_inst_pe_1_2_3_n4), .A2(
        npu_inst_pe_1_2_3_n7), .A3(npu_inst_pe_1_2_3_n6), .ZN(
        npu_inst_pe_1_2_3_n48) );
  INV_X1 npu_inst_pe_1_2_3_U25 ( .A(npu_inst_pe_1_2_3_n4), .ZN(
        npu_inst_pe_1_2_3_n3) );
  OR3_X1 npu_inst_pe_1_2_3_U24 ( .A1(npu_inst_pe_1_2_3_n3), .A2(
        npu_inst_pe_1_2_3_n7), .A3(npu_inst_pe_1_2_3_n6), .ZN(
        npu_inst_pe_1_2_3_n52) );
  OR3_X1 npu_inst_pe_1_2_3_U23 ( .A1(npu_inst_pe_1_2_3_n5), .A2(
        npu_inst_pe_1_2_3_n7), .A3(npu_inst_pe_1_2_3_n3), .ZN(
        npu_inst_pe_1_2_3_n60) );
  BUF_X1 npu_inst_pe_1_2_3_U22 ( .A(npu_inst_n25), .Z(npu_inst_pe_1_2_3_n1) );
  NOR2_X1 npu_inst_pe_1_2_3_U21 ( .A1(npu_inst_pe_1_2_3_n60), .A2(
        npu_inst_pe_1_2_3_n2), .ZN(npu_inst_pe_1_2_3_n58) );
  NOR2_X1 npu_inst_pe_1_2_3_U20 ( .A1(npu_inst_pe_1_2_3_n56), .A2(
        npu_inst_pe_1_2_3_n2), .ZN(npu_inst_pe_1_2_3_n54) );
  NOR2_X1 npu_inst_pe_1_2_3_U19 ( .A1(npu_inst_pe_1_2_3_n52), .A2(
        npu_inst_pe_1_2_3_n2), .ZN(npu_inst_pe_1_2_3_n50) );
  NOR2_X1 npu_inst_pe_1_2_3_U18 ( .A1(npu_inst_pe_1_2_3_n48), .A2(
        npu_inst_pe_1_2_3_n2), .ZN(npu_inst_pe_1_2_3_n46) );
  NOR2_X1 npu_inst_pe_1_2_3_U17 ( .A1(npu_inst_pe_1_2_3_n40), .A2(
        npu_inst_pe_1_2_3_n2), .ZN(npu_inst_pe_1_2_3_n38) );
  NOR2_X1 npu_inst_pe_1_2_3_U16 ( .A1(npu_inst_pe_1_2_3_n44), .A2(
        npu_inst_pe_1_2_3_n2), .ZN(npu_inst_pe_1_2_3_n42) );
  BUF_X1 npu_inst_pe_1_2_3_U15 ( .A(npu_inst_n85), .Z(npu_inst_pe_1_2_3_n7) );
  INV_X1 npu_inst_pe_1_2_3_U14 ( .A(npu_inst_n107), .ZN(npu_inst_pe_1_2_3_n11)
         );
  INV_X1 npu_inst_pe_1_2_3_U13 ( .A(npu_inst_pe_1_2_3_n38), .ZN(
        npu_inst_pe_1_2_3_n113) );
  INV_X1 npu_inst_pe_1_2_3_U12 ( .A(npu_inst_pe_1_2_3_n58), .ZN(
        npu_inst_pe_1_2_3_n118) );
  INV_X1 npu_inst_pe_1_2_3_U11 ( .A(npu_inst_pe_1_2_3_n54), .ZN(
        npu_inst_pe_1_2_3_n117) );
  INV_X1 npu_inst_pe_1_2_3_U10 ( .A(npu_inst_pe_1_2_3_n50), .ZN(
        npu_inst_pe_1_2_3_n116) );
  INV_X1 npu_inst_pe_1_2_3_U9 ( .A(npu_inst_pe_1_2_3_n46), .ZN(
        npu_inst_pe_1_2_3_n115) );
  INV_X1 npu_inst_pe_1_2_3_U8 ( .A(npu_inst_pe_1_2_3_n42), .ZN(
        npu_inst_pe_1_2_3_n114) );
  BUF_X1 npu_inst_pe_1_2_3_U7 ( .A(npu_inst_pe_1_2_3_n11), .Z(
        npu_inst_pe_1_2_3_n10) );
  BUF_X1 npu_inst_pe_1_2_3_U6 ( .A(npu_inst_pe_1_2_3_n11), .Z(
        npu_inst_pe_1_2_3_n9) );
  BUF_X1 npu_inst_pe_1_2_3_U5 ( .A(npu_inst_pe_1_2_3_n11), .Z(
        npu_inst_pe_1_2_3_n8) );
  NOR2_X1 npu_inst_pe_1_2_3_U4 ( .A1(npu_inst_pe_1_2_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_3_n1), .ZN(npu_inst_pe_1_2_3_n76) );
  NOR2_X1 npu_inst_pe_1_2_3_U3 ( .A1(npu_inst_pe_1_2_3_n27), .A2(
        npu_inst_pe_1_2_3_n1), .ZN(npu_inst_pe_1_2_3_n77) );
  FA_X1 npu_inst_pe_1_2_3_sub_77_U2_1 ( .A(npu_inst_int_data_res_2__3__1_), 
        .B(npu_inst_pe_1_2_3_n13), .CI(npu_inst_pe_1_2_3_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_2_3_sub_77_carry_2_), .S(npu_inst_pe_1_2_3_N66) );
  FA_X1 npu_inst_pe_1_2_3_add_79_U1_1 ( .A(npu_inst_int_data_res_2__3__1_), 
        .B(npu_inst_pe_1_2_3_int_data_1_), .CI(
        npu_inst_pe_1_2_3_add_79_carry_1_), .CO(
        npu_inst_pe_1_2_3_add_79_carry_2_), .S(npu_inst_pe_1_2_3_N74) );
  NAND3_X1 npu_inst_pe_1_2_3_U101 ( .A1(npu_inst_pe_1_2_3_n4), .A2(
        npu_inst_pe_1_2_3_n6), .A3(npu_inst_pe_1_2_3_n7), .ZN(
        npu_inst_pe_1_2_3_n44) );
  NAND3_X1 npu_inst_pe_1_2_3_U100 ( .A1(npu_inst_pe_1_2_3_n3), .A2(
        npu_inst_pe_1_2_3_n6), .A3(npu_inst_pe_1_2_3_n7), .ZN(
        npu_inst_pe_1_2_3_n40) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_3_n33), .CK(
        npu_inst_pe_1_2_3_net4041), .RN(npu_inst_pe_1_2_3_n8), .Q(
        npu_inst_int_data_res_2__3__6_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_3_n34), .CK(
        npu_inst_pe_1_2_3_net4041), .RN(npu_inst_pe_1_2_3_n8), .Q(
        npu_inst_int_data_res_2__3__5_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_3_n35), .CK(
        npu_inst_pe_1_2_3_net4041), .RN(npu_inst_pe_1_2_3_n8), .Q(
        npu_inst_int_data_res_2__3__4_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_3_n36), .CK(
        npu_inst_pe_1_2_3_net4041), .RN(npu_inst_pe_1_2_3_n8), .Q(
        npu_inst_int_data_res_2__3__3_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_3_n98), .CK(
        npu_inst_pe_1_2_3_net4041), .RN(npu_inst_pe_1_2_3_n8), .Q(
        npu_inst_int_data_res_2__3__2_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_3_n99), .CK(
        npu_inst_pe_1_2_3_net4041), .RN(npu_inst_pe_1_2_3_n8), .Q(
        npu_inst_int_data_res_2__3__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_3_n32), .CK(
        npu_inst_pe_1_2_3_net4041), .RN(npu_inst_pe_1_2_3_n8), .Q(
        npu_inst_int_data_res_2__3__7_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_3_n100), 
        .CK(npu_inst_pe_1_2_3_net4041), .RN(npu_inst_pe_1_2_3_n8), .Q(
        npu_inst_int_data_res_2__3__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_weight_reg_0_ ( .D(npu_inst_n93), .CK(
        npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n8), .Q(
        npu_inst_pe_1_2_3_int_q_weight_0_), .QN(npu_inst_pe_1_2_3_n27) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_weight_reg_1_ ( .D(npu_inst_n99), .CK(
        npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n8), .Q(
        npu_inst_pe_1_2_3_int_q_weight_1_), .QN(npu_inst_pe_1_2_3_n26) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_3_n112), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n8), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_3_n106), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n8), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_3_n111), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_3_n105), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_3_n110), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_3_n104), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_3_n109), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_3_n103), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_3_n108), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_3_n102), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_3_n107), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_3_n101), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_3_n86), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_3_n87), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n9), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_3_n88), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_3_n89), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_3_n90), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_3_n91), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_3_n92), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_3_n93), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_3_n94), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_3_n95), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_3_n96), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_3_n97), 
        .CK(npu_inst_pe_1_2_3_net4047), .RN(npu_inst_pe_1_2_3_n10), .Q(
        npu_inst_pe_1_2_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_3_net4041) );
  CLKGATETST_X1 npu_inst_pe_1_2_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n47), .SE(1'b0), .GCK(npu_inst_pe_1_2_3_net4047) );
  MUX2_X1 npu_inst_pe_1_2_4_U153 ( .A(npu_inst_pe_1_2_4_n31), .B(
        npu_inst_pe_1_2_4_n28), .S(npu_inst_pe_1_2_4_n7), .Z(
        npu_inst_pe_1_2_4_N93) );
  MUX2_X1 npu_inst_pe_1_2_4_U152 ( .A(npu_inst_pe_1_2_4_n30), .B(
        npu_inst_pe_1_2_4_n29), .S(npu_inst_pe_1_2_4_n5), .Z(
        npu_inst_pe_1_2_4_n31) );
  MUX2_X1 npu_inst_pe_1_2_4_U151 ( .A(npu_inst_pe_1_2_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_4_n3), .Z(
        npu_inst_pe_1_2_4_n30) );
  MUX2_X1 npu_inst_pe_1_2_4_U150 ( .A(npu_inst_pe_1_2_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_4_n3), .Z(
        npu_inst_pe_1_2_4_n29) );
  MUX2_X1 npu_inst_pe_1_2_4_U149 ( .A(npu_inst_pe_1_2_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_4_n3), .Z(
        npu_inst_pe_1_2_4_n28) );
  MUX2_X1 npu_inst_pe_1_2_4_U148 ( .A(npu_inst_pe_1_2_4_n25), .B(
        npu_inst_pe_1_2_4_n22), .S(npu_inst_pe_1_2_4_n7), .Z(
        npu_inst_pe_1_2_4_N94) );
  MUX2_X1 npu_inst_pe_1_2_4_U147 ( .A(npu_inst_pe_1_2_4_n24), .B(
        npu_inst_pe_1_2_4_n23), .S(npu_inst_pe_1_2_4_n5), .Z(
        npu_inst_pe_1_2_4_n25) );
  MUX2_X1 npu_inst_pe_1_2_4_U146 ( .A(npu_inst_pe_1_2_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_4_n3), .Z(
        npu_inst_pe_1_2_4_n24) );
  MUX2_X1 npu_inst_pe_1_2_4_U145 ( .A(npu_inst_pe_1_2_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_4_n3), .Z(
        npu_inst_pe_1_2_4_n23) );
  MUX2_X1 npu_inst_pe_1_2_4_U144 ( .A(npu_inst_pe_1_2_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_4_n3), .Z(
        npu_inst_pe_1_2_4_n22) );
  MUX2_X1 npu_inst_pe_1_2_4_U143 ( .A(npu_inst_pe_1_2_4_n21), .B(
        npu_inst_pe_1_2_4_n18), .S(npu_inst_pe_1_2_4_n7), .Z(
        npu_inst_int_data_x_2__4__1_) );
  MUX2_X1 npu_inst_pe_1_2_4_U142 ( .A(npu_inst_pe_1_2_4_n20), .B(
        npu_inst_pe_1_2_4_n19), .S(npu_inst_pe_1_2_4_n5), .Z(
        npu_inst_pe_1_2_4_n21) );
  MUX2_X1 npu_inst_pe_1_2_4_U141 ( .A(npu_inst_pe_1_2_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_4_n3), .Z(
        npu_inst_pe_1_2_4_n20) );
  MUX2_X1 npu_inst_pe_1_2_4_U140 ( .A(npu_inst_pe_1_2_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_4_n3), .Z(
        npu_inst_pe_1_2_4_n19) );
  MUX2_X1 npu_inst_pe_1_2_4_U139 ( .A(npu_inst_pe_1_2_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_4_n3), .Z(
        npu_inst_pe_1_2_4_n18) );
  MUX2_X1 npu_inst_pe_1_2_4_U138 ( .A(npu_inst_pe_1_2_4_n17), .B(
        npu_inst_pe_1_2_4_n14), .S(npu_inst_pe_1_2_4_n7), .Z(
        npu_inst_int_data_x_2__4__0_) );
  MUX2_X1 npu_inst_pe_1_2_4_U137 ( .A(npu_inst_pe_1_2_4_n16), .B(
        npu_inst_pe_1_2_4_n15), .S(npu_inst_pe_1_2_4_n5), .Z(
        npu_inst_pe_1_2_4_n17) );
  MUX2_X1 npu_inst_pe_1_2_4_U136 ( .A(npu_inst_pe_1_2_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_4_n3), .Z(
        npu_inst_pe_1_2_4_n16) );
  MUX2_X1 npu_inst_pe_1_2_4_U135 ( .A(npu_inst_pe_1_2_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_4_n3), .Z(
        npu_inst_pe_1_2_4_n15) );
  MUX2_X1 npu_inst_pe_1_2_4_U134 ( .A(npu_inst_pe_1_2_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_4_n3), .Z(
        npu_inst_pe_1_2_4_n14) );
  XOR2_X1 npu_inst_pe_1_2_4_U133 ( .A(npu_inst_pe_1_2_4_int_data_0_), .B(
        npu_inst_int_data_res_2__4__0_), .Z(npu_inst_pe_1_2_4_N73) );
  AND2_X1 npu_inst_pe_1_2_4_U132 ( .A1(npu_inst_int_data_res_2__4__0_), .A2(
        npu_inst_pe_1_2_4_int_data_0_), .ZN(npu_inst_pe_1_2_4_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_4_U131 ( .A(npu_inst_int_data_res_2__4__0_), .B(
        npu_inst_pe_1_2_4_n12), .ZN(npu_inst_pe_1_2_4_N65) );
  OR2_X1 npu_inst_pe_1_2_4_U130 ( .A1(npu_inst_pe_1_2_4_n12), .A2(
        npu_inst_int_data_res_2__4__0_), .ZN(npu_inst_pe_1_2_4_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_4_U129 ( .A(npu_inst_int_data_res_2__4__2_), .B(
        npu_inst_pe_1_2_4_add_79_carry_2_), .Z(npu_inst_pe_1_2_4_N75) );
  AND2_X1 npu_inst_pe_1_2_4_U128 ( .A1(npu_inst_pe_1_2_4_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_2__4__2_), .ZN(
        npu_inst_pe_1_2_4_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_4_U127 ( .A(npu_inst_int_data_res_2__4__3_), .B(
        npu_inst_pe_1_2_4_add_79_carry_3_), .Z(npu_inst_pe_1_2_4_N76) );
  AND2_X1 npu_inst_pe_1_2_4_U126 ( .A1(npu_inst_pe_1_2_4_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_2__4__3_), .ZN(
        npu_inst_pe_1_2_4_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_4_U125 ( .A(npu_inst_int_data_res_2__4__4_), .B(
        npu_inst_pe_1_2_4_add_79_carry_4_), .Z(npu_inst_pe_1_2_4_N77) );
  AND2_X1 npu_inst_pe_1_2_4_U124 ( .A1(npu_inst_pe_1_2_4_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_2__4__4_), .ZN(
        npu_inst_pe_1_2_4_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_4_U123 ( .A(npu_inst_int_data_res_2__4__5_), .B(
        npu_inst_pe_1_2_4_add_79_carry_5_), .Z(npu_inst_pe_1_2_4_N78) );
  AND2_X1 npu_inst_pe_1_2_4_U122 ( .A1(npu_inst_pe_1_2_4_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_2__4__5_), .ZN(
        npu_inst_pe_1_2_4_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_4_U121 ( .A(npu_inst_int_data_res_2__4__6_), .B(
        npu_inst_pe_1_2_4_add_79_carry_6_), .Z(npu_inst_pe_1_2_4_N79) );
  AND2_X1 npu_inst_pe_1_2_4_U120 ( .A1(npu_inst_pe_1_2_4_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_2__4__6_), .ZN(
        npu_inst_pe_1_2_4_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_4_U119 ( .A(npu_inst_int_data_res_2__4__7_), .B(
        npu_inst_pe_1_2_4_add_79_carry_7_), .Z(npu_inst_pe_1_2_4_N80) );
  XNOR2_X1 npu_inst_pe_1_2_4_U118 ( .A(npu_inst_pe_1_2_4_sub_77_carry_2_), .B(
        npu_inst_int_data_res_2__4__2_), .ZN(npu_inst_pe_1_2_4_N67) );
  OR2_X1 npu_inst_pe_1_2_4_U117 ( .A1(npu_inst_int_data_res_2__4__2_), .A2(
        npu_inst_pe_1_2_4_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_2_4_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_4_U116 ( .A(npu_inst_pe_1_2_4_sub_77_carry_3_), .B(
        npu_inst_int_data_res_2__4__3_), .ZN(npu_inst_pe_1_2_4_N68) );
  OR2_X1 npu_inst_pe_1_2_4_U115 ( .A1(npu_inst_int_data_res_2__4__3_), .A2(
        npu_inst_pe_1_2_4_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_2_4_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_4_U114 ( .A(npu_inst_pe_1_2_4_sub_77_carry_4_), .B(
        npu_inst_int_data_res_2__4__4_), .ZN(npu_inst_pe_1_2_4_N69) );
  OR2_X1 npu_inst_pe_1_2_4_U113 ( .A1(npu_inst_int_data_res_2__4__4_), .A2(
        npu_inst_pe_1_2_4_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_2_4_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_4_U112 ( .A(npu_inst_pe_1_2_4_sub_77_carry_5_), .B(
        npu_inst_int_data_res_2__4__5_), .ZN(npu_inst_pe_1_2_4_N70) );
  OR2_X1 npu_inst_pe_1_2_4_U111 ( .A1(npu_inst_int_data_res_2__4__5_), .A2(
        npu_inst_pe_1_2_4_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_2_4_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_4_U110 ( .A(npu_inst_pe_1_2_4_sub_77_carry_6_), .B(
        npu_inst_int_data_res_2__4__6_), .ZN(npu_inst_pe_1_2_4_N71) );
  OR2_X1 npu_inst_pe_1_2_4_U109 ( .A1(npu_inst_int_data_res_2__4__6_), .A2(
        npu_inst_pe_1_2_4_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_2_4_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_4_U108 ( .A(npu_inst_int_data_res_2__4__7_), .B(
        npu_inst_pe_1_2_4_sub_77_carry_7_), .ZN(npu_inst_pe_1_2_4_N72) );
  INV_X1 npu_inst_pe_1_2_4_U107 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_2_4_n6)
         );
  INV_X1 npu_inst_pe_1_2_4_U106 ( .A(npu_inst_pe_1_2_4_n6), .ZN(
        npu_inst_pe_1_2_4_n5) );
  INV_X1 npu_inst_pe_1_2_4_U105 ( .A(npu_inst_n40), .ZN(npu_inst_pe_1_2_4_n2)
         );
  AOI22_X1 npu_inst_pe_1_2_4_U104 ( .A1(npu_inst_int_data_y_3__4__0_), .A2(
        npu_inst_pe_1_2_4_n58), .B1(npu_inst_pe_1_2_4_n118), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_4_n57) );
  INV_X1 npu_inst_pe_1_2_4_U103 ( .A(npu_inst_pe_1_2_4_n57), .ZN(
        npu_inst_pe_1_2_4_n107) );
  AOI22_X1 npu_inst_pe_1_2_4_U102 ( .A1(npu_inst_int_data_y_3__4__0_), .A2(
        npu_inst_pe_1_2_4_n54), .B1(npu_inst_pe_1_2_4_n117), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_4_n53) );
  INV_X1 npu_inst_pe_1_2_4_U99 ( .A(npu_inst_pe_1_2_4_n53), .ZN(
        npu_inst_pe_1_2_4_n108) );
  AOI22_X1 npu_inst_pe_1_2_4_U98 ( .A1(npu_inst_int_data_y_3__4__0_), .A2(
        npu_inst_pe_1_2_4_n50), .B1(npu_inst_pe_1_2_4_n116), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_4_n49) );
  INV_X1 npu_inst_pe_1_2_4_U97 ( .A(npu_inst_pe_1_2_4_n49), .ZN(
        npu_inst_pe_1_2_4_n109) );
  AOI22_X1 npu_inst_pe_1_2_4_U96 ( .A1(npu_inst_int_data_y_3__4__0_), .A2(
        npu_inst_pe_1_2_4_n46), .B1(npu_inst_pe_1_2_4_n115), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_4_n45) );
  INV_X1 npu_inst_pe_1_2_4_U95 ( .A(npu_inst_pe_1_2_4_n45), .ZN(
        npu_inst_pe_1_2_4_n110) );
  AOI22_X1 npu_inst_pe_1_2_4_U94 ( .A1(npu_inst_int_data_y_3__4__0_), .A2(
        npu_inst_pe_1_2_4_n42), .B1(npu_inst_pe_1_2_4_n114), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_4_n41) );
  INV_X1 npu_inst_pe_1_2_4_U93 ( .A(npu_inst_pe_1_2_4_n41), .ZN(
        npu_inst_pe_1_2_4_n111) );
  AOI22_X1 npu_inst_pe_1_2_4_U92 ( .A1(npu_inst_int_data_y_3__4__1_), .A2(
        npu_inst_pe_1_2_4_n58), .B1(npu_inst_pe_1_2_4_n118), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_4_n59) );
  INV_X1 npu_inst_pe_1_2_4_U91 ( .A(npu_inst_pe_1_2_4_n59), .ZN(
        npu_inst_pe_1_2_4_n101) );
  AOI22_X1 npu_inst_pe_1_2_4_U90 ( .A1(npu_inst_int_data_y_3__4__1_), .A2(
        npu_inst_pe_1_2_4_n54), .B1(npu_inst_pe_1_2_4_n117), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_4_n55) );
  INV_X1 npu_inst_pe_1_2_4_U89 ( .A(npu_inst_pe_1_2_4_n55), .ZN(
        npu_inst_pe_1_2_4_n102) );
  AOI22_X1 npu_inst_pe_1_2_4_U88 ( .A1(npu_inst_int_data_y_3__4__1_), .A2(
        npu_inst_pe_1_2_4_n50), .B1(npu_inst_pe_1_2_4_n116), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_4_n51) );
  INV_X1 npu_inst_pe_1_2_4_U87 ( .A(npu_inst_pe_1_2_4_n51), .ZN(
        npu_inst_pe_1_2_4_n103) );
  AOI22_X1 npu_inst_pe_1_2_4_U86 ( .A1(npu_inst_int_data_y_3__4__1_), .A2(
        npu_inst_pe_1_2_4_n46), .B1(npu_inst_pe_1_2_4_n115), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_4_n47) );
  INV_X1 npu_inst_pe_1_2_4_U85 ( .A(npu_inst_pe_1_2_4_n47), .ZN(
        npu_inst_pe_1_2_4_n104) );
  AOI22_X1 npu_inst_pe_1_2_4_U84 ( .A1(npu_inst_int_data_y_3__4__1_), .A2(
        npu_inst_pe_1_2_4_n42), .B1(npu_inst_pe_1_2_4_n114), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_4_n43) );
  INV_X1 npu_inst_pe_1_2_4_U83 ( .A(npu_inst_pe_1_2_4_n43), .ZN(
        npu_inst_pe_1_2_4_n105) );
  AOI22_X1 npu_inst_pe_1_2_4_U82 ( .A1(npu_inst_pe_1_2_4_n38), .A2(
        npu_inst_int_data_y_3__4__1_), .B1(npu_inst_pe_1_2_4_n113), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_4_n39) );
  INV_X1 npu_inst_pe_1_2_4_U81 ( .A(npu_inst_pe_1_2_4_n39), .ZN(
        npu_inst_pe_1_2_4_n106) );
  AND2_X1 npu_inst_pe_1_2_4_U80 ( .A1(npu_inst_pe_1_2_4_N93), .A2(npu_inst_n40), .ZN(npu_inst_int_data_y_2__4__0_) );
  NAND2_X1 npu_inst_pe_1_2_4_U79 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_4_n60), .ZN(npu_inst_pe_1_2_4_n74) );
  OAI21_X1 npu_inst_pe_1_2_4_U78 ( .B1(npu_inst_pe_1_2_4_n63), .B2(
        npu_inst_pe_1_2_4_n60), .A(npu_inst_pe_1_2_4_n74), .ZN(
        npu_inst_pe_1_2_4_n97) );
  NAND2_X1 npu_inst_pe_1_2_4_U77 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_4_n60), .ZN(npu_inst_pe_1_2_4_n73) );
  OAI21_X1 npu_inst_pe_1_2_4_U76 ( .B1(npu_inst_pe_1_2_4_n61), .B2(
        npu_inst_pe_1_2_4_n60), .A(npu_inst_pe_1_2_4_n73), .ZN(
        npu_inst_pe_1_2_4_n96) );
  NAND2_X1 npu_inst_pe_1_2_4_U75 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_4_n56), .ZN(npu_inst_pe_1_2_4_n72) );
  OAI21_X1 npu_inst_pe_1_2_4_U74 ( .B1(npu_inst_pe_1_2_4_n63), .B2(
        npu_inst_pe_1_2_4_n56), .A(npu_inst_pe_1_2_4_n72), .ZN(
        npu_inst_pe_1_2_4_n95) );
  NAND2_X1 npu_inst_pe_1_2_4_U73 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_4_n56), .ZN(npu_inst_pe_1_2_4_n71) );
  OAI21_X1 npu_inst_pe_1_2_4_U72 ( .B1(npu_inst_pe_1_2_4_n61), .B2(
        npu_inst_pe_1_2_4_n56), .A(npu_inst_pe_1_2_4_n71), .ZN(
        npu_inst_pe_1_2_4_n94) );
  NAND2_X1 npu_inst_pe_1_2_4_U71 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_4_n52), .ZN(npu_inst_pe_1_2_4_n70) );
  OAI21_X1 npu_inst_pe_1_2_4_U70 ( .B1(npu_inst_pe_1_2_4_n63), .B2(
        npu_inst_pe_1_2_4_n52), .A(npu_inst_pe_1_2_4_n70), .ZN(
        npu_inst_pe_1_2_4_n93) );
  NAND2_X1 npu_inst_pe_1_2_4_U69 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_4_n52), .ZN(npu_inst_pe_1_2_4_n69) );
  OAI21_X1 npu_inst_pe_1_2_4_U68 ( .B1(npu_inst_pe_1_2_4_n61), .B2(
        npu_inst_pe_1_2_4_n52), .A(npu_inst_pe_1_2_4_n69), .ZN(
        npu_inst_pe_1_2_4_n92) );
  NAND2_X1 npu_inst_pe_1_2_4_U67 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_4_n48), .ZN(npu_inst_pe_1_2_4_n68) );
  OAI21_X1 npu_inst_pe_1_2_4_U66 ( .B1(npu_inst_pe_1_2_4_n63), .B2(
        npu_inst_pe_1_2_4_n48), .A(npu_inst_pe_1_2_4_n68), .ZN(
        npu_inst_pe_1_2_4_n91) );
  NAND2_X1 npu_inst_pe_1_2_4_U65 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_4_n48), .ZN(npu_inst_pe_1_2_4_n67) );
  OAI21_X1 npu_inst_pe_1_2_4_U64 ( .B1(npu_inst_pe_1_2_4_n61), .B2(
        npu_inst_pe_1_2_4_n48), .A(npu_inst_pe_1_2_4_n67), .ZN(
        npu_inst_pe_1_2_4_n90) );
  NAND2_X1 npu_inst_pe_1_2_4_U63 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_4_n44), .ZN(npu_inst_pe_1_2_4_n66) );
  OAI21_X1 npu_inst_pe_1_2_4_U62 ( .B1(npu_inst_pe_1_2_4_n63), .B2(
        npu_inst_pe_1_2_4_n44), .A(npu_inst_pe_1_2_4_n66), .ZN(
        npu_inst_pe_1_2_4_n89) );
  NAND2_X1 npu_inst_pe_1_2_4_U61 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_4_n44), .ZN(npu_inst_pe_1_2_4_n65) );
  OAI21_X1 npu_inst_pe_1_2_4_U60 ( .B1(npu_inst_pe_1_2_4_n61), .B2(
        npu_inst_pe_1_2_4_n44), .A(npu_inst_pe_1_2_4_n65), .ZN(
        npu_inst_pe_1_2_4_n88) );
  NAND2_X1 npu_inst_pe_1_2_4_U59 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_4_n40), .ZN(npu_inst_pe_1_2_4_n64) );
  OAI21_X1 npu_inst_pe_1_2_4_U58 ( .B1(npu_inst_pe_1_2_4_n63), .B2(
        npu_inst_pe_1_2_4_n40), .A(npu_inst_pe_1_2_4_n64), .ZN(
        npu_inst_pe_1_2_4_n87) );
  NAND2_X1 npu_inst_pe_1_2_4_U57 ( .A1(npu_inst_pe_1_2_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_4_n40), .ZN(npu_inst_pe_1_2_4_n62) );
  OAI21_X1 npu_inst_pe_1_2_4_U56 ( .B1(npu_inst_pe_1_2_4_n61), .B2(
        npu_inst_pe_1_2_4_n40), .A(npu_inst_pe_1_2_4_n62), .ZN(
        npu_inst_pe_1_2_4_n86) );
  AOI22_X1 npu_inst_pe_1_2_4_U55 ( .A1(npu_inst_pe_1_2_4_n38), .A2(
        npu_inst_int_data_y_3__4__0_), .B1(npu_inst_pe_1_2_4_n113), .B2(
        npu_inst_pe_1_2_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_4_n37) );
  INV_X1 npu_inst_pe_1_2_4_U54 ( .A(npu_inst_pe_1_2_4_n37), .ZN(
        npu_inst_pe_1_2_4_n112) );
  AND2_X1 npu_inst_pe_1_2_4_U53 ( .A1(npu_inst_n40), .A2(npu_inst_pe_1_2_4_N94), .ZN(npu_inst_int_data_y_2__4__1_) );
  AOI222_X1 npu_inst_pe_1_2_4_U52 ( .A1(npu_inst_int_data_res_3__4__0_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N73), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N65), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n84) );
  INV_X1 npu_inst_pe_1_2_4_U51 ( .A(npu_inst_pe_1_2_4_n84), .ZN(
        npu_inst_pe_1_2_4_n100) );
  AOI222_X1 npu_inst_pe_1_2_4_U50 ( .A1(npu_inst_pe_1_2_4_n1), .A2(
        npu_inst_int_data_res_3__4__7_), .B1(npu_inst_pe_1_2_4_N80), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N72), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n75) );
  INV_X1 npu_inst_pe_1_2_4_U49 ( .A(npu_inst_pe_1_2_4_n75), .ZN(
        npu_inst_pe_1_2_4_n32) );
  AOI222_X1 npu_inst_pe_1_2_4_U48 ( .A1(npu_inst_int_data_res_3__4__1_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N74), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N66), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n83) );
  INV_X1 npu_inst_pe_1_2_4_U47 ( .A(npu_inst_pe_1_2_4_n83), .ZN(
        npu_inst_pe_1_2_4_n99) );
  AOI222_X1 npu_inst_pe_1_2_4_U46 ( .A1(npu_inst_int_data_res_3__4__3_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N76), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N68), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n81) );
  INV_X1 npu_inst_pe_1_2_4_U45 ( .A(npu_inst_pe_1_2_4_n81), .ZN(
        npu_inst_pe_1_2_4_n36) );
  AOI222_X1 npu_inst_pe_1_2_4_U44 ( .A1(npu_inst_int_data_res_3__4__4_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N77), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N69), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n80) );
  INV_X1 npu_inst_pe_1_2_4_U43 ( .A(npu_inst_pe_1_2_4_n80), .ZN(
        npu_inst_pe_1_2_4_n35) );
  AOI222_X1 npu_inst_pe_1_2_4_U42 ( .A1(npu_inst_int_data_res_3__4__5_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N78), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N70), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n79) );
  INV_X1 npu_inst_pe_1_2_4_U41 ( .A(npu_inst_pe_1_2_4_n79), .ZN(
        npu_inst_pe_1_2_4_n34) );
  AOI222_X1 npu_inst_pe_1_2_4_U40 ( .A1(npu_inst_int_data_res_3__4__6_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N79), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N71), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n78) );
  INV_X1 npu_inst_pe_1_2_4_U39 ( .A(npu_inst_pe_1_2_4_n78), .ZN(
        npu_inst_pe_1_2_4_n33) );
  AND2_X1 npu_inst_pe_1_2_4_U38 ( .A1(npu_inst_int_data_x_2__4__1_), .A2(
        npu_inst_pe_1_2_4_int_q_weight_1_), .ZN(npu_inst_pe_1_2_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_4_U37 ( .A1(npu_inst_int_data_x_2__4__0_), .A2(
        npu_inst_pe_1_2_4_int_q_weight_1_), .ZN(npu_inst_pe_1_2_4_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_2_4_U36 ( .A(npu_inst_pe_1_2_4_int_data_1_), .ZN(
        npu_inst_pe_1_2_4_n13) );
  NOR3_X1 npu_inst_pe_1_2_4_U35 ( .A1(npu_inst_pe_1_2_4_n26), .A2(npu_inst_n40), .A3(npu_inst_int_ckg[43]), .ZN(npu_inst_pe_1_2_4_n85) );
  OR2_X1 npu_inst_pe_1_2_4_U34 ( .A1(npu_inst_pe_1_2_4_n85), .A2(
        npu_inst_pe_1_2_4_n1), .ZN(npu_inst_pe_1_2_4_N84) );
  AOI222_X1 npu_inst_pe_1_2_4_U33 ( .A1(npu_inst_int_data_res_3__4__2_), .A2(
        npu_inst_pe_1_2_4_n1), .B1(npu_inst_pe_1_2_4_N75), .B2(
        npu_inst_pe_1_2_4_n76), .C1(npu_inst_pe_1_2_4_N67), .C2(
        npu_inst_pe_1_2_4_n77), .ZN(npu_inst_pe_1_2_4_n82) );
  INV_X1 npu_inst_pe_1_2_4_U32 ( .A(npu_inst_pe_1_2_4_n82), .ZN(
        npu_inst_pe_1_2_4_n98) );
  AOI22_X1 npu_inst_pe_1_2_4_U31 ( .A1(npu_inst_n40), .A2(
        npu_inst_int_data_y_3__4__1_), .B1(npu_inst_pe_1_2_4_n2), .B2(
        npu_inst_int_data_x_2__5__1_), .ZN(npu_inst_pe_1_2_4_n63) );
  AOI22_X1 npu_inst_pe_1_2_4_U30 ( .A1(npu_inst_n40), .A2(
        npu_inst_int_data_y_3__4__0_), .B1(npu_inst_pe_1_2_4_n2), .B2(
        npu_inst_int_data_x_2__5__0_), .ZN(npu_inst_pe_1_2_4_n61) );
  INV_X1 npu_inst_pe_1_2_4_U29 ( .A(npu_inst_pe_1_2_4_int_data_0_), .ZN(
        npu_inst_pe_1_2_4_n12) );
  INV_X1 npu_inst_pe_1_2_4_U28 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_2_4_n4)
         );
  OR3_X1 npu_inst_pe_1_2_4_U27 ( .A1(npu_inst_pe_1_2_4_n5), .A2(
        npu_inst_pe_1_2_4_n7), .A3(npu_inst_pe_1_2_4_n4), .ZN(
        npu_inst_pe_1_2_4_n56) );
  OR3_X1 npu_inst_pe_1_2_4_U26 ( .A1(npu_inst_pe_1_2_4_n4), .A2(
        npu_inst_pe_1_2_4_n7), .A3(npu_inst_pe_1_2_4_n6), .ZN(
        npu_inst_pe_1_2_4_n48) );
  INV_X1 npu_inst_pe_1_2_4_U25 ( .A(npu_inst_pe_1_2_4_n4), .ZN(
        npu_inst_pe_1_2_4_n3) );
  OR3_X1 npu_inst_pe_1_2_4_U24 ( .A1(npu_inst_pe_1_2_4_n3), .A2(
        npu_inst_pe_1_2_4_n7), .A3(npu_inst_pe_1_2_4_n6), .ZN(
        npu_inst_pe_1_2_4_n52) );
  OR3_X1 npu_inst_pe_1_2_4_U23 ( .A1(npu_inst_pe_1_2_4_n5), .A2(
        npu_inst_pe_1_2_4_n7), .A3(npu_inst_pe_1_2_4_n3), .ZN(
        npu_inst_pe_1_2_4_n60) );
  BUF_X1 npu_inst_pe_1_2_4_U22 ( .A(npu_inst_n25), .Z(npu_inst_pe_1_2_4_n1) );
  NOR2_X1 npu_inst_pe_1_2_4_U21 ( .A1(npu_inst_pe_1_2_4_n60), .A2(
        npu_inst_pe_1_2_4_n2), .ZN(npu_inst_pe_1_2_4_n58) );
  NOR2_X1 npu_inst_pe_1_2_4_U20 ( .A1(npu_inst_pe_1_2_4_n56), .A2(
        npu_inst_pe_1_2_4_n2), .ZN(npu_inst_pe_1_2_4_n54) );
  NOR2_X1 npu_inst_pe_1_2_4_U19 ( .A1(npu_inst_pe_1_2_4_n52), .A2(
        npu_inst_pe_1_2_4_n2), .ZN(npu_inst_pe_1_2_4_n50) );
  NOR2_X1 npu_inst_pe_1_2_4_U18 ( .A1(npu_inst_pe_1_2_4_n48), .A2(
        npu_inst_pe_1_2_4_n2), .ZN(npu_inst_pe_1_2_4_n46) );
  NOR2_X1 npu_inst_pe_1_2_4_U17 ( .A1(npu_inst_pe_1_2_4_n40), .A2(
        npu_inst_pe_1_2_4_n2), .ZN(npu_inst_pe_1_2_4_n38) );
  NOR2_X1 npu_inst_pe_1_2_4_U16 ( .A1(npu_inst_pe_1_2_4_n44), .A2(
        npu_inst_pe_1_2_4_n2), .ZN(npu_inst_pe_1_2_4_n42) );
  BUF_X1 npu_inst_pe_1_2_4_U15 ( .A(npu_inst_n84), .Z(npu_inst_pe_1_2_4_n7) );
  INV_X1 npu_inst_pe_1_2_4_U14 ( .A(npu_inst_n107), .ZN(npu_inst_pe_1_2_4_n11)
         );
  INV_X1 npu_inst_pe_1_2_4_U13 ( .A(npu_inst_pe_1_2_4_n38), .ZN(
        npu_inst_pe_1_2_4_n113) );
  INV_X1 npu_inst_pe_1_2_4_U12 ( .A(npu_inst_pe_1_2_4_n58), .ZN(
        npu_inst_pe_1_2_4_n118) );
  INV_X1 npu_inst_pe_1_2_4_U11 ( .A(npu_inst_pe_1_2_4_n54), .ZN(
        npu_inst_pe_1_2_4_n117) );
  INV_X1 npu_inst_pe_1_2_4_U10 ( .A(npu_inst_pe_1_2_4_n50), .ZN(
        npu_inst_pe_1_2_4_n116) );
  INV_X1 npu_inst_pe_1_2_4_U9 ( .A(npu_inst_pe_1_2_4_n46), .ZN(
        npu_inst_pe_1_2_4_n115) );
  INV_X1 npu_inst_pe_1_2_4_U8 ( .A(npu_inst_pe_1_2_4_n42), .ZN(
        npu_inst_pe_1_2_4_n114) );
  BUF_X1 npu_inst_pe_1_2_4_U7 ( .A(npu_inst_pe_1_2_4_n11), .Z(
        npu_inst_pe_1_2_4_n10) );
  BUF_X1 npu_inst_pe_1_2_4_U6 ( .A(npu_inst_pe_1_2_4_n11), .Z(
        npu_inst_pe_1_2_4_n9) );
  BUF_X1 npu_inst_pe_1_2_4_U5 ( .A(npu_inst_pe_1_2_4_n11), .Z(
        npu_inst_pe_1_2_4_n8) );
  NOR2_X1 npu_inst_pe_1_2_4_U4 ( .A1(npu_inst_pe_1_2_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_4_n1), .ZN(npu_inst_pe_1_2_4_n76) );
  NOR2_X1 npu_inst_pe_1_2_4_U3 ( .A1(npu_inst_pe_1_2_4_n27), .A2(
        npu_inst_pe_1_2_4_n1), .ZN(npu_inst_pe_1_2_4_n77) );
  FA_X1 npu_inst_pe_1_2_4_sub_77_U2_1 ( .A(npu_inst_int_data_res_2__4__1_), 
        .B(npu_inst_pe_1_2_4_n13), .CI(npu_inst_pe_1_2_4_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_2_4_sub_77_carry_2_), .S(npu_inst_pe_1_2_4_N66) );
  FA_X1 npu_inst_pe_1_2_4_add_79_U1_1 ( .A(npu_inst_int_data_res_2__4__1_), 
        .B(npu_inst_pe_1_2_4_int_data_1_), .CI(
        npu_inst_pe_1_2_4_add_79_carry_1_), .CO(
        npu_inst_pe_1_2_4_add_79_carry_2_), .S(npu_inst_pe_1_2_4_N74) );
  NAND3_X1 npu_inst_pe_1_2_4_U101 ( .A1(npu_inst_pe_1_2_4_n4), .A2(
        npu_inst_pe_1_2_4_n6), .A3(npu_inst_pe_1_2_4_n7), .ZN(
        npu_inst_pe_1_2_4_n44) );
  NAND3_X1 npu_inst_pe_1_2_4_U100 ( .A1(npu_inst_pe_1_2_4_n3), .A2(
        npu_inst_pe_1_2_4_n6), .A3(npu_inst_pe_1_2_4_n7), .ZN(
        npu_inst_pe_1_2_4_n40) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_4_n33), .CK(
        npu_inst_pe_1_2_4_net4018), .RN(npu_inst_pe_1_2_4_n8), .Q(
        npu_inst_int_data_res_2__4__6_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_4_n34), .CK(
        npu_inst_pe_1_2_4_net4018), .RN(npu_inst_pe_1_2_4_n8), .Q(
        npu_inst_int_data_res_2__4__5_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_4_n35), .CK(
        npu_inst_pe_1_2_4_net4018), .RN(npu_inst_pe_1_2_4_n8), .Q(
        npu_inst_int_data_res_2__4__4_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_4_n36), .CK(
        npu_inst_pe_1_2_4_net4018), .RN(npu_inst_pe_1_2_4_n8), .Q(
        npu_inst_int_data_res_2__4__3_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_4_n98), .CK(
        npu_inst_pe_1_2_4_net4018), .RN(npu_inst_pe_1_2_4_n8), .Q(
        npu_inst_int_data_res_2__4__2_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_4_n99), .CK(
        npu_inst_pe_1_2_4_net4018), .RN(npu_inst_pe_1_2_4_n8), .Q(
        npu_inst_int_data_res_2__4__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_4_n32), .CK(
        npu_inst_pe_1_2_4_net4018), .RN(npu_inst_pe_1_2_4_n8), .Q(
        npu_inst_int_data_res_2__4__7_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_4_n100), 
        .CK(npu_inst_pe_1_2_4_net4018), .RN(npu_inst_pe_1_2_4_n8), .Q(
        npu_inst_int_data_res_2__4__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_weight_reg_0_ ( .D(npu_inst_n93), .CK(
        npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n8), .Q(
        npu_inst_pe_1_2_4_int_q_weight_0_), .QN(npu_inst_pe_1_2_4_n27) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_weight_reg_1_ ( .D(npu_inst_n99), .CK(
        npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n8), .Q(
        npu_inst_pe_1_2_4_int_q_weight_1_), .QN(npu_inst_pe_1_2_4_n26) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_4_n112), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n8), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_4_n106), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n8), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_4_n111), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_4_n105), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_4_n110), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_4_n104), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_4_n109), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_4_n103), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_4_n108), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_4_n102), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_4_n107), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_4_n101), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_4_n86), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_4_n87), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n9), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_4_n88), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_4_n89), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_4_n90), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_4_n91), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_4_n92), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_4_n93), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_4_n94), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_4_n95), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_4_n96), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_4_n97), 
        .CK(npu_inst_pe_1_2_4_net4024), .RN(npu_inst_pe_1_2_4_n10), .Q(
        npu_inst_pe_1_2_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_4_net4018) );
  CLKGATETST_X1 npu_inst_pe_1_2_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n46), .SE(1'b0), .GCK(npu_inst_pe_1_2_4_net4024) );
  MUX2_X1 npu_inst_pe_1_2_5_U153 ( .A(npu_inst_pe_1_2_5_n31), .B(
        npu_inst_pe_1_2_5_n28), .S(npu_inst_pe_1_2_5_n7), .Z(
        npu_inst_pe_1_2_5_N93) );
  MUX2_X1 npu_inst_pe_1_2_5_U152 ( .A(npu_inst_pe_1_2_5_n30), .B(
        npu_inst_pe_1_2_5_n29), .S(npu_inst_pe_1_2_5_n5), .Z(
        npu_inst_pe_1_2_5_n31) );
  MUX2_X1 npu_inst_pe_1_2_5_U151 ( .A(npu_inst_pe_1_2_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_5_n3), .Z(
        npu_inst_pe_1_2_5_n30) );
  MUX2_X1 npu_inst_pe_1_2_5_U150 ( .A(npu_inst_pe_1_2_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_5_n3), .Z(
        npu_inst_pe_1_2_5_n29) );
  MUX2_X1 npu_inst_pe_1_2_5_U149 ( .A(npu_inst_pe_1_2_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_5_n3), .Z(
        npu_inst_pe_1_2_5_n28) );
  MUX2_X1 npu_inst_pe_1_2_5_U148 ( .A(npu_inst_pe_1_2_5_n25), .B(
        npu_inst_pe_1_2_5_n22), .S(npu_inst_pe_1_2_5_n7), .Z(
        npu_inst_pe_1_2_5_N94) );
  MUX2_X1 npu_inst_pe_1_2_5_U147 ( .A(npu_inst_pe_1_2_5_n24), .B(
        npu_inst_pe_1_2_5_n23), .S(npu_inst_pe_1_2_5_n5), .Z(
        npu_inst_pe_1_2_5_n25) );
  MUX2_X1 npu_inst_pe_1_2_5_U146 ( .A(npu_inst_pe_1_2_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_5_n3), .Z(
        npu_inst_pe_1_2_5_n24) );
  MUX2_X1 npu_inst_pe_1_2_5_U145 ( .A(npu_inst_pe_1_2_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_5_n3), .Z(
        npu_inst_pe_1_2_5_n23) );
  MUX2_X1 npu_inst_pe_1_2_5_U144 ( .A(npu_inst_pe_1_2_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_5_n3), .Z(
        npu_inst_pe_1_2_5_n22) );
  MUX2_X1 npu_inst_pe_1_2_5_U143 ( .A(npu_inst_pe_1_2_5_n21), .B(
        npu_inst_pe_1_2_5_n18), .S(npu_inst_pe_1_2_5_n7), .Z(
        npu_inst_int_data_x_2__5__1_) );
  MUX2_X1 npu_inst_pe_1_2_5_U142 ( .A(npu_inst_pe_1_2_5_n20), .B(
        npu_inst_pe_1_2_5_n19), .S(npu_inst_pe_1_2_5_n5), .Z(
        npu_inst_pe_1_2_5_n21) );
  MUX2_X1 npu_inst_pe_1_2_5_U141 ( .A(npu_inst_pe_1_2_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_5_n3), .Z(
        npu_inst_pe_1_2_5_n20) );
  MUX2_X1 npu_inst_pe_1_2_5_U140 ( .A(npu_inst_pe_1_2_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_5_n3), .Z(
        npu_inst_pe_1_2_5_n19) );
  MUX2_X1 npu_inst_pe_1_2_5_U139 ( .A(npu_inst_pe_1_2_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_5_n3), .Z(
        npu_inst_pe_1_2_5_n18) );
  MUX2_X1 npu_inst_pe_1_2_5_U138 ( .A(npu_inst_pe_1_2_5_n17), .B(
        npu_inst_pe_1_2_5_n14), .S(npu_inst_pe_1_2_5_n7), .Z(
        npu_inst_int_data_x_2__5__0_) );
  MUX2_X1 npu_inst_pe_1_2_5_U137 ( .A(npu_inst_pe_1_2_5_n16), .B(
        npu_inst_pe_1_2_5_n15), .S(npu_inst_pe_1_2_5_n5), .Z(
        npu_inst_pe_1_2_5_n17) );
  MUX2_X1 npu_inst_pe_1_2_5_U136 ( .A(npu_inst_pe_1_2_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_5_n3), .Z(
        npu_inst_pe_1_2_5_n16) );
  MUX2_X1 npu_inst_pe_1_2_5_U135 ( .A(npu_inst_pe_1_2_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_5_n3), .Z(
        npu_inst_pe_1_2_5_n15) );
  MUX2_X1 npu_inst_pe_1_2_5_U134 ( .A(npu_inst_pe_1_2_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_5_n3), .Z(
        npu_inst_pe_1_2_5_n14) );
  XOR2_X1 npu_inst_pe_1_2_5_U133 ( .A(npu_inst_pe_1_2_5_int_data_0_), .B(
        npu_inst_int_data_res_2__5__0_), .Z(npu_inst_pe_1_2_5_N73) );
  AND2_X1 npu_inst_pe_1_2_5_U132 ( .A1(npu_inst_int_data_res_2__5__0_), .A2(
        npu_inst_pe_1_2_5_int_data_0_), .ZN(npu_inst_pe_1_2_5_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_5_U131 ( .A(npu_inst_int_data_res_2__5__0_), .B(
        npu_inst_pe_1_2_5_n12), .ZN(npu_inst_pe_1_2_5_N65) );
  OR2_X1 npu_inst_pe_1_2_5_U130 ( .A1(npu_inst_pe_1_2_5_n12), .A2(
        npu_inst_int_data_res_2__5__0_), .ZN(npu_inst_pe_1_2_5_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_5_U129 ( .A(npu_inst_int_data_res_2__5__2_), .B(
        npu_inst_pe_1_2_5_add_79_carry_2_), .Z(npu_inst_pe_1_2_5_N75) );
  AND2_X1 npu_inst_pe_1_2_5_U128 ( .A1(npu_inst_pe_1_2_5_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_2__5__2_), .ZN(
        npu_inst_pe_1_2_5_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_5_U127 ( .A(npu_inst_int_data_res_2__5__3_), .B(
        npu_inst_pe_1_2_5_add_79_carry_3_), .Z(npu_inst_pe_1_2_5_N76) );
  AND2_X1 npu_inst_pe_1_2_5_U126 ( .A1(npu_inst_pe_1_2_5_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_2__5__3_), .ZN(
        npu_inst_pe_1_2_5_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_5_U125 ( .A(npu_inst_int_data_res_2__5__4_), .B(
        npu_inst_pe_1_2_5_add_79_carry_4_), .Z(npu_inst_pe_1_2_5_N77) );
  AND2_X1 npu_inst_pe_1_2_5_U124 ( .A1(npu_inst_pe_1_2_5_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_2__5__4_), .ZN(
        npu_inst_pe_1_2_5_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_5_U123 ( .A(npu_inst_int_data_res_2__5__5_), .B(
        npu_inst_pe_1_2_5_add_79_carry_5_), .Z(npu_inst_pe_1_2_5_N78) );
  AND2_X1 npu_inst_pe_1_2_5_U122 ( .A1(npu_inst_pe_1_2_5_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_2__5__5_), .ZN(
        npu_inst_pe_1_2_5_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_5_U121 ( .A(npu_inst_int_data_res_2__5__6_), .B(
        npu_inst_pe_1_2_5_add_79_carry_6_), .Z(npu_inst_pe_1_2_5_N79) );
  AND2_X1 npu_inst_pe_1_2_5_U120 ( .A1(npu_inst_pe_1_2_5_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_2__5__6_), .ZN(
        npu_inst_pe_1_2_5_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_5_U119 ( .A(npu_inst_int_data_res_2__5__7_), .B(
        npu_inst_pe_1_2_5_add_79_carry_7_), .Z(npu_inst_pe_1_2_5_N80) );
  XNOR2_X1 npu_inst_pe_1_2_5_U118 ( .A(npu_inst_pe_1_2_5_sub_77_carry_2_), .B(
        npu_inst_int_data_res_2__5__2_), .ZN(npu_inst_pe_1_2_5_N67) );
  OR2_X1 npu_inst_pe_1_2_5_U117 ( .A1(npu_inst_int_data_res_2__5__2_), .A2(
        npu_inst_pe_1_2_5_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_2_5_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_5_U116 ( .A(npu_inst_pe_1_2_5_sub_77_carry_3_), .B(
        npu_inst_int_data_res_2__5__3_), .ZN(npu_inst_pe_1_2_5_N68) );
  OR2_X1 npu_inst_pe_1_2_5_U115 ( .A1(npu_inst_int_data_res_2__5__3_), .A2(
        npu_inst_pe_1_2_5_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_2_5_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_5_U114 ( .A(npu_inst_pe_1_2_5_sub_77_carry_4_), .B(
        npu_inst_int_data_res_2__5__4_), .ZN(npu_inst_pe_1_2_5_N69) );
  OR2_X1 npu_inst_pe_1_2_5_U113 ( .A1(npu_inst_int_data_res_2__5__4_), .A2(
        npu_inst_pe_1_2_5_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_2_5_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_5_U112 ( .A(npu_inst_pe_1_2_5_sub_77_carry_5_), .B(
        npu_inst_int_data_res_2__5__5_), .ZN(npu_inst_pe_1_2_5_N70) );
  OR2_X1 npu_inst_pe_1_2_5_U111 ( .A1(npu_inst_int_data_res_2__5__5_), .A2(
        npu_inst_pe_1_2_5_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_2_5_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_5_U110 ( .A(npu_inst_pe_1_2_5_sub_77_carry_6_), .B(
        npu_inst_int_data_res_2__5__6_), .ZN(npu_inst_pe_1_2_5_N71) );
  OR2_X1 npu_inst_pe_1_2_5_U109 ( .A1(npu_inst_int_data_res_2__5__6_), .A2(
        npu_inst_pe_1_2_5_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_2_5_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_5_U108 ( .A(npu_inst_int_data_res_2__5__7_), .B(
        npu_inst_pe_1_2_5_sub_77_carry_7_), .ZN(npu_inst_pe_1_2_5_N72) );
  INV_X1 npu_inst_pe_1_2_5_U107 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_2_5_n6)
         );
  INV_X1 npu_inst_pe_1_2_5_U106 ( .A(npu_inst_pe_1_2_5_n6), .ZN(
        npu_inst_pe_1_2_5_n5) );
  INV_X1 npu_inst_pe_1_2_5_U105 ( .A(npu_inst_n40), .ZN(npu_inst_pe_1_2_5_n2)
         );
  AOI22_X1 npu_inst_pe_1_2_5_U104 ( .A1(npu_inst_int_data_y_3__5__0_), .A2(
        npu_inst_pe_1_2_5_n58), .B1(npu_inst_pe_1_2_5_n118), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_5_n57) );
  INV_X1 npu_inst_pe_1_2_5_U103 ( .A(npu_inst_pe_1_2_5_n57), .ZN(
        npu_inst_pe_1_2_5_n107) );
  AOI22_X1 npu_inst_pe_1_2_5_U102 ( .A1(npu_inst_int_data_y_3__5__0_), .A2(
        npu_inst_pe_1_2_5_n54), .B1(npu_inst_pe_1_2_5_n117), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_5_n53) );
  INV_X1 npu_inst_pe_1_2_5_U99 ( .A(npu_inst_pe_1_2_5_n53), .ZN(
        npu_inst_pe_1_2_5_n108) );
  AOI22_X1 npu_inst_pe_1_2_5_U98 ( .A1(npu_inst_int_data_y_3__5__0_), .A2(
        npu_inst_pe_1_2_5_n50), .B1(npu_inst_pe_1_2_5_n116), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_5_n49) );
  INV_X1 npu_inst_pe_1_2_5_U97 ( .A(npu_inst_pe_1_2_5_n49), .ZN(
        npu_inst_pe_1_2_5_n109) );
  AOI22_X1 npu_inst_pe_1_2_5_U96 ( .A1(npu_inst_int_data_y_3__5__0_), .A2(
        npu_inst_pe_1_2_5_n46), .B1(npu_inst_pe_1_2_5_n115), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_5_n45) );
  INV_X1 npu_inst_pe_1_2_5_U95 ( .A(npu_inst_pe_1_2_5_n45), .ZN(
        npu_inst_pe_1_2_5_n110) );
  AOI22_X1 npu_inst_pe_1_2_5_U94 ( .A1(npu_inst_int_data_y_3__5__0_), .A2(
        npu_inst_pe_1_2_5_n42), .B1(npu_inst_pe_1_2_5_n114), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_5_n41) );
  INV_X1 npu_inst_pe_1_2_5_U93 ( .A(npu_inst_pe_1_2_5_n41), .ZN(
        npu_inst_pe_1_2_5_n111) );
  AOI22_X1 npu_inst_pe_1_2_5_U92 ( .A1(npu_inst_int_data_y_3__5__1_), .A2(
        npu_inst_pe_1_2_5_n58), .B1(npu_inst_pe_1_2_5_n118), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_5_n59) );
  INV_X1 npu_inst_pe_1_2_5_U91 ( .A(npu_inst_pe_1_2_5_n59), .ZN(
        npu_inst_pe_1_2_5_n101) );
  AOI22_X1 npu_inst_pe_1_2_5_U90 ( .A1(npu_inst_int_data_y_3__5__1_), .A2(
        npu_inst_pe_1_2_5_n54), .B1(npu_inst_pe_1_2_5_n117), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_5_n55) );
  INV_X1 npu_inst_pe_1_2_5_U89 ( .A(npu_inst_pe_1_2_5_n55), .ZN(
        npu_inst_pe_1_2_5_n102) );
  AOI22_X1 npu_inst_pe_1_2_5_U88 ( .A1(npu_inst_int_data_y_3__5__1_), .A2(
        npu_inst_pe_1_2_5_n50), .B1(npu_inst_pe_1_2_5_n116), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_5_n51) );
  INV_X1 npu_inst_pe_1_2_5_U87 ( .A(npu_inst_pe_1_2_5_n51), .ZN(
        npu_inst_pe_1_2_5_n103) );
  AOI22_X1 npu_inst_pe_1_2_5_U86 ( .A1(npu_inst_int_data_y_3__5__1_), .A2(
        npu_inst_pe_1_2_5_n46), .B1(npu_inst_pe_1_2_5_n115), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_5_n47) );
  INV_X1 npu_inst_pe_1_2_5_U85 ( .A(npu_inst_pe_1_2_5_n47), .ZN(
        npu_inst_pe_1_2_5_n104) );
  AOI22_X1 npu_inst_pe_1_2_5_U84 ( .A1(npu_inst_int_data_y_3__5__1_), .A2(
        npu_inst_pe_1_2_5_n42), .B1(npu_inst_pe_1_2_5_n114), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_5_n43) );
  INV_X1 npu_inst_pe_1_2_5_U83 ( .A(npu_inst_pe_1_2_5_n43), .ZN(
        npu_inst_pe_1_2_5_n105) );
  AOI22_X1 npu_inst_pe_1_2_5_U82 ( .A1(npu_inst_pe_1_2_5_n38), .A2(
        npu_inst_int_data_y_3__5__1_), .B1(npu_inst_pe_1_2_5_n113), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_5_n39) );
  INV_X1 npu_inst_pe_1_2_5_U81 ( .A(npu_inst_pe_1_2_5_n39), .ZN(
        npu_inst_pe_1_2_5_n106) );
  AND2_X1 npu_inst_pe_1_2_5_U80 ( .A1(npu_inst_pe_1_2_5_N93), .A2(npu_inst_n40), .ZN(npu_inst_int_data_y_2__5__0_) );
  NAND2_X1 npu_inst_pe_1_2_5_U79 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_5_n60), .ZN(npu_inst_pe_1_2_5_n74) );
  OAI21_X1 npu_inst_pe_1_2_5_U78 ( .B1(npu_inst_pe_1_2_5_n63), .B2(
        npu_inst_pe_1_2_5_n60), .A(npu_inst_pe_1_2_5_n74), .ZN(
        npu_inst_pe_1_2_5_n97) );
  NAND2_X1 npu_inst_pe_1_2_5_U77 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_5_n60), .ZN(npu_inst_pe_1_2_5_n73) );
  OAI21_X1 npu_inst_pe_1_2_5_U76 ( .B1(npu_inst_pe_1_2_5_n61), .B2(
        npu_inst_pe_1_2_5_n60), .A(npu_inst_pe_1_2_5_n73), .ZN(
        npu_inst_pe_1_2_5_n96) );
  NAND2_X1 npu_inst_pe_1_2_5_U75 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_5_n56), .ZN(npu_inst_pe_1_2_5_n72) );
  OAI21_X1 npu_inst_pe_1_2_5_U74 ( .B1(npu_inst_pe_1_2_5_n63), .B2(
        npu_inst_pe_1_2_5_n56), .A(npu_inst_pe_1_2_5_n72), .ZN(
        npu_inst_pe_1_2_5_n95) );
  NAND2_X1 npu_inst_pe_1_2_5_U73 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_5_n56), .ZN(npu_inst_pe_1_2_5_n71) );
  OAI21_X1 npu_inst_pe_1_2_5_U72 ( .B1(npu_inst_pe_1_2_5_n61), .B2(
        npu_inst_pe_1_2_5_n56), .A(npu_inst_pe_1_2_5_n71), .ZN(
        npu_inst_pe_1_2_5_n94) );
  NAND2_X1 npu_inst_pe_1_2_5_U71 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_5_n52), .ZN(npu_inst_pe_1_2_5_n70) );
  OAI21_X1 npu_inst_pe_1_2_5_U70 ( .B1(npu_inst_pe_1_2_5_n63), .B2(
        npu_inst_pe_1_2_5_n52), .A(npu_inst_pe_1_2_5_n70), .ZN(
        npu_inst_pe_1_2_5_n93) );
  NAND2_X1 npu_inst_pe_1_2_5_U69 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_5_n52), .ZN(npu_inst_pe_1_2_5_n69) );
  OAI21_X1 npu_inst_pe_1_2_5_U68 ( .B1(npu_inst_pe_1_2_5_n61), .B2(
        npu_inst_pe_1_2_5_n52), .A(npu_inst_pe_1_2_5_n69), .ZN(
        npu_inst_pe_1_2_5_n92) );
  NAND2_X1 npu_inst_pe_1_2_5_U67 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_5_n48), .ZN(npu_inst_pe_1_2_5_n68) );
  OAI21_X1 npu_inst_pe_1_2_5_U66 ( .B1(npu_inst_pe_1_2_5_n63), .B2(
        npu_inst_pe_1_2_5_n48), .A(npu_inst_pe_1_2_5_n68), .ZN(
        npu_inst_pe_1_2_5_n91) );
  NAND2_X1 npu_inst_pe_1_2_5_U65 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_5_n48), .ZN(npu_inst_pe_1_2_5_n67) );
  OAI21_X1 npu_inst_pe_1_2_5_U64 ( .B1(npu_inst_pe_1_2_5_n61), .B2(
        npu_inst_pe_1_2_5_n48), .A(npu_inst_pe_1_2_5_n67), .ZN(
        npu_inst_pe_1_2_5_n90) );
  NAND2_X1 npu_inst_pe_1_2_5_U63 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_5_n44), .ZN(npu_inst_pe_1_2_5_n66) );
  OAI21_X1 npu_inst_pe_1_2_5_U62 ( .B1(npu_inst_pe_1_2_5_n63), .B2(
        npu_inst_pe_1_2_5_n44), .A(npu_inst_pe_1_2_5_n66), .ZN(
        npu_inst_pe_1_2_5_n89) );
  NAND2_X1 npu_inst_pe_1_2_5_U61 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_5_n44), .ZN(npu_inst_pe_1_2_5_n65) );
  OAI21_X1 npu_inst_pe_1_2_5_U60 ( .B1(npu_inst_pe_1_2_5_n61), .B2(
        npu_inst_pe_1_2_5_n44), .A(npu_inst_pe_1_2_5_n65), .ZN(
        npu_inst_pe_1_2_5_n88) );
  NAND2_X1 npu_inst_pe_1_2_5_U59 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_5_n40), .ZN(npu_inst_pe_1_2_5_n64) );
  OAI21_X1 npu_inst_pe_1_2_5_U58 ( .B1(npu_inst_pe_1_2_5_n63), .B2(
        npu_inst_pe_1_2_5_n40), .A(npu_inst_pe_1_2_5_n64), .ZN(
        npu_inst_pe_1_2_5_n87) );
  NAND2_X1 npu_inst_pe_1_2_5_U57 ( .A1(npu_inst_pe_1_2_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_5_n40), .ZN(npu_inst_pe_1_2_5_n62) );
  OAI21_X1 npu_inst_pe_1_2_5_U56 ( .B1(npu_inst_pe_1_2_5_n61), .B2(
        npu_inst_pe_1_2_5_n40), .A(npu_inst_pe_1_2_5_n62), .ZN(
        npu_inst_pe_1_2_5_n86) );
  AOI22_X1 npu_inst_pe_1_2_5_U55 ( .A1(npu_inst_pe_1_2_5_n38), .A2(
        npu_inst_int_data_y_3__5__0_), .B1(npu_inst_pe_1_2_5_n113), .B2(
        npu_inst_pe_1_2_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_5_n37) );
  INV_X1 npu_inst_pe_1_2_5_U54 ( .A(npu_inst_pe_1_2_5_n37), .ZN(
        npu_inst_pe_1_2_5_n112) );
  AND2_X1 npu_inst_pe_1_2_5_U53 ( .A1(npu_inst_n40), .A2(npu_inst_pe_1_2_5_N94), .ZN(npu_inst_int_data_y_2__5__1_) );
  AOI222_X1 npu_inst_pe_1_2_5_U52 ( .A1(npu_inst_int_data_res_3__5__0_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N73), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N65), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n84) );
  INV_X1 npu_inst_pe_1_2_5_U51 ( .A(npu_inst_pe_1_2_5_n84), .ZN(
        npu_inst_pe_1_2_5_n100) );
  AOI222_X1 npu_inst_pe_1_2_5_U50 ( .A1(npu_inst_pe_1_2_5_n1), .A2(
        npu_inst_int_data_res_3__5__7_), .B1(npu_inst_pe_1_2_5_N80), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N72), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n75) );
  INV_X1 npu_inst_pe_1_2_5_U49 ( .A(npu_inst_pe_1_2_5_n75), .ZN(
        npu_inst_pe_1_2_5_n32) );
  AOI222_X1 npu_inst_pe_1_2_5_U48 ( .A1(npu_inst_int_data_res_3__5__1_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N74), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N66), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n83) );
  INV_X1 npu_inst_pe_1_2_5_U47 ( .A(npu_inst_pe_1_2_5_n83), .ZN(
        npu_inst_pe_1_2_5_n99) );
  AOI222_X1 npu_inst_pe_1_2_5_U46 ( .A1(npu_inst_int_data_res_3__5__3_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N76), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N68), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n81) );
  INV_X1 npu_inst_pe_1_2_5_U45 ( .A(npu_inst_pe_1_2_5_n81), .ZN(
        npu_inst_pe_1_2_5_n36) );
  AOI222_X1 npu_inst_pe_1_2_5_U44 ( .A1(npu_inst_int_data_res_3__5__4_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N77), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N69), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n80) );
  INV_X1 npu_inst_pe_1_2_5_U43 ( .A(npu_inst_pe_1_2_5_n80), .ZN(
        npu_inst_pe_1_2_5_n35) );
  AOI222_X1 npu_inst_pe_1_2_5_U42 ( .A1(npu_inst_int_data_res_3__5__5_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N78), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N70), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n79) );
  INV_X1 npu_inst_pe_1_2_5_U41 ( .A(npu_inst_pe_1_2_5_n79), .ZN(
        npu_inst_pe_1_2_5_n34) );
  AOI222_X1 npu_inst_pe_1_2_5_U40 ( .A1(npu_inst_int_data_res_3__5__6_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N79), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N71), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n78) );
  INV_X1 npu_inst_pe_1_2_5_U39 ( .A(npu_inst_pe_1_2_5_n78), .ZN(
        npu_inst_pe_1_2_5_n33) );
  AND2_X1 npu_inst_pe_1_2_5_U38 ( .A1(npu_inst_int_data_x_2__5__1_), .A2(
        npu_inst_pe_1_2_5_int_q_weight_1_), .ZN(npu_inst_pe_1_2_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_5_U37 ( .A1(npu_inst_int_data_x_2__5__0_), .A2(
        npu_inst_pe_1_2_5_int_q_weight_1_), .ZN(npu_inst_pe_1_2_5_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_2_5_U36 ( .A(npu_inst_pe_1_2_5_int_data_1_), .ZN(
        npu_inst_pe_1_2_5_n13) );
  NOR3_X1 npu_inst_pe_1_2_5_U35 ( .A1(npu_inst_pe_1_2_5_n26), .A2(npu_inst_n40), .A3(npu_inst_int_ckg[42]), .ZN(npu_inst_pe_1_2_5_n85) );
  OR2_X1 npu_inst_pe_1_2_5_U34 ( .A1(npu_inst_pe_1_2_5_n85), .A2(
        npu_inst_pe_1_2_5_n1), .ZN(npu_inst_pe_1_2_5_N84) );
  AOI222_X1 npu_inst_pe_1_2_5_U33 ( .A1(npu_inst_int_data_res_3__5__2_), .A2(
        npu_inst_pe_1_2_5_n1), .B1(npu_inst_pe_1_2_5_N75), .B2(
        npu_inst_pe_1_2_5_n76), .C1(npu_inst_pe_1_2_5_N67), .C2(
        npu_inst_pe_1_2_5_n77), .ZN(npu_inst_pe_1_2_5_n82) );
  INV_X1 npu_inst_pe_1_2_5_U32 ( .A(npu_inst_pe_1_2_5_n82), .ZN(
        npu_inst_pe_1_2_5_n98) );
  AOI22_X1 npu_inst_pe_1_2_5_U31 ( .A1(npu_inst_n40), .A2(
        npu_inst_int_data_y_3__5__1_), .B1(npu_inst_pe_1_2_5_n2), .B2(
        npu_inst_int_data_x_2__6__1_), .ZN(npu_inst_pe_1_2_5_n63) );
  AOI22_X1 npu_inst_pe_1_2_5_U30 ( .A1(npu_inst_n40), .A2(
        npu_inst_int_data_y_3__5__0_), .B1(npu_inst_pe_1_2_5_n2), .B2(
        npu_inst_int_data_x_2__6__0_), .ZN(npu_inst_pe_1_2_5_n61) );
  INV_X1 npu_inst_pe_1_2_5_U29 ( .A(npu_inst_pe_1_2_5_int_data_0_), .ZN(
        npu_inst_pe_1_2_5_n12) );
  INV_X1 npu_inst_pe_1_2_5_U28 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_2_5_n4)
         );
  OR3_X1 npu_inst_pe_1_2_5_U27 ( .A1(npu_inst_pe_1_2_5_n5), .A2(
        npu_inst_pe_1_2_5_n7), .A3(npu_inst_pe_1_2_5_n4), .ZN(
        npu_inst_pe_1_2_5_n56) );
  OR3_X1 npu_inst_pe_1_2_5_U26 ( .A1(npu_inst_pe_1_2_5_n4), .A2(
        npu_inst_pe_1_2_5_n7), .A3(npu_inst_pe_1_2_5_n6), .ZN(
        npu_inst_pe_1_2_5_n48) );
  INV_X1 npu_inst_pe_1_2_5_U25 ( .A(npu_inst_pe_1_2_5_n4), .ZN(
        npu_inst_pe_1_2_5_n3) );
  OR3_X1 npu_inst_pe_1_2_5_U24 ( .A1(npu_inst_pe_1_2_5_n3), .A2(
        npu_inst_pe_1_2_5_n7), .A3(npu_inst_pe_1_2_5_n6), .ZN(
        npu_inst_pe_1_2_5_n52) );
  OR3_X1 npu_inst_pe_1_2_5_U23 ( .A1(npu_inst_pe_1_2_5_n5), .A2(
        npu_inst_pe_1_2_5_n7), .A3(npu_inst_pe_1_2_5_n3), .ZN(
        npu_inst_pe_1_2_5_n60) );
  BUF_X1 npu_inst_pe_1_2_5_U22 ( .A(npu_inst_n25), .Z(npu_inst_pe_1_2_5_n1) );
  NOR2_X1 npu_inst_pe_1_2_5_U21 ( .A1(npu_inst_pe_1_2_5_n60), .A2(
        npu_inst_pe_1_2_5_n2), .ZN(npu_inst_pe_1_2_5_n58) );
  NOR2_X1 npu_inst_pe_1_2_5_U20 ( .A1(npu_inst_pe_1_2_5_n56), .A2(
        npu_inst_pe_1_2_5_n2), .ZN(npu_inst_pe_1_2_5_n54) );
  NOR2_X1 npu_inst_pe_1_2_5_U19 ( .A1(npu_inst_pe_1_2_5_n52), .A2(
        npu_inst_pe_1_2_5_n2), .ZN(npu_inst_pe_1_2_5_n50) );
  NOR2_X1 npu_inst_pe_1_2_5_U18 ( .A1(npu_inst_pe_1_2_5_n48), .A2(
        npu_inst_pe_1_2_5_n2), .ZN(npu_inst_pe_1_2_5_n46) );
  NOR2_X1 npu_inst_pe_1_2_5_U17 ( .A1(npu_inst_pe_1_2_5_n40), .A2(
        npu_inst_pe_1_2_5_n2), .ZN(npu_inst_pe_1_2_5_n38) );
  NOR2_X1 npu_inst_pe_1_2_5_U16 ( .A1(npu_inst_pe_1_2_5_n44), .A2(
        npu_inst_pe_1_2_5_n2), .ZN(npu_inst_pe_1_2_5_n42) );
  BUF_X1 npu_inst_pe_1_2_5_U15 ( .A(npu_inst_n84), .Z(npu_inst_pe_1_2_5_n7) );
  INV_X1 npu_inst_pe_1_2_5_U14 ( .A(npu_inst_n107), .ZN(npu_inst_pe_1_2_5_n11)
         );
  INV_X1 npu_inst_pe_1_2_5_U13 ( .A(npu_inst_pe_1_2_5_n38), .ZN(
        npu_inst_pe_1_2_5_n113) );
  INV_X1 npu_inst_pe_1_2_5_U12 ( .A(npu_inst_pe_1_2_5_n58), .ZN(
        npu_inst_pe_1_2_5_n118) );
  INV_X1 npu_inst_pe_1_2_5_U11 ( .A(npu_inst_pe_1_2_5_n54), .ZN(
        npu_inst_pe_1_2_5_n117) );
  INV_X1 npu_inst_pe_1_2_5_U10 ( .A(npu_inst_pe_1_2_5_n50), .ZN(
        npu_inst_pe_1_2_5_n116) );
  INV_X1 npu_inst_pe_1_2_5_U9 ( .A(npu_inst_pe_1_2_5_n46), .ZN(
        npu_inst_pe_1_2_5_n115) );
  INV_X1 npu_inst_pe_1_2_5_U8 ( .A(npu_inst_pe_1_2_5_n42), .ZN(
        npu_inst_pe_1_2_5_n114) );
  BUF_X1 npu_inst_pe_1_2_5_U7 ( .A(npu_inst_pe_1_2_5_n11), .Z(
        npu_inst_pe_1_2_5_n10) );
  BUF_X1 npu_inst_pe_1_2_5_U6 ( .A(npu_inst_pe_1_2_5_n11), .Z(
        npu_inst_pe_1_2_5_n9) );
  BUF_X1 npu_inst_pe_1_2_5_U5 ( .A(npu_inst_pe_1_2_5_n11), .Z(
        npu_inst_pe_1_2_5_n8) );
  NOR2_X1 npu_inst_pe_1_2_5_U4 ( .A1(npu_inst_pe_1_2_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_5_n1), .ZN(npu_inst_pe_1_2_5_n76) );
  NOR2_X1 npu_inst_pe_1_2_5_U3 ( .A1(npu_inst_pe_1_2_5_n27), .A2(
        npu_inst_pe_1_2_5_n1), .ZN(npu_inst_pe_1_2_5_n77) );
  FA_X1 npu_inst_pe_1_2_5_sub_77_U2_1 ( .A(npu_inst_int_data_res_2__5__1_), 
        .B(npu_inst_pe_1_2_5_n13), .CI(npu_inst_pe_1_2_5_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_2_5_sub_77_carry_2_), .S(npu_inst_pe_1_2_5_N66) );
  FA_X1 npu_inst_pe_1_2_5_add_79_U1_1 ( .A(npu_inst_int_data_res_2__5__1_), 
        .B(npu_inst_pe_1_2_5_int_data_1_), .CI(
        npu_inst_pe_1_2_5_add_79_carry_1_), .CO(
        npu_inst_pe_1_2_5_add_79_carry_2_), .S(npu_inst_pe_1_2_5_N74) );
  NAND3_X1 npu_inst_pe_1_2_5_U101 ( .A1(npu_inst_pe_1_2_5_n4), .A2(
        npu_inst_pe_1_2_5_n6), .A3(npu_inst_pe_1_2_5_n7), .ZN(
        npu_inst_pe_1_2_5_n44) );
  NAND3_X1 npu_inst_pe_1_2_5_U100 ( .A1(npu_inst_pe_1_2_5_n3), .A2(
        npu_inst_pe_1_2_5_n6), .A3(npu_inst_pe_1_2_5_n7), .ZN(
        npu_inst_pe_1_2_5_n40) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_5_n33), .CK(
        npu_inst_pe_1_2_5_net3995), .RN(npu_inst_pe_1_2_5_n8), .Q(
        npu_inst_int_data_res_2__5__6_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_5_n34), .CK(
        npu_inst_pe_1_2_5_net3995), .RN(npu_inst_pe_1_2_5_n8), .Q(
        npu_inst_int_data_res_2__5__5_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_5_n35), .CK(
        npu_inst_pe_1_2_5_net3995), .RN(npu_inst_pe_1_2_5_n8), .Q(
        npu_inst_int_data_res_2__5__4_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_5_n36), .CK(
        npu_inst_pe_1_2_5_net3995), .RN(npu_inst_pe_1_2_5_n8), .Q(
        npu_inst_int_data_res_2__5__3_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_5_n98), .CK(
        npu_inst_pe_1_2_5_net3995), .RN(npu_inst_pe_1_2_5_n8), .Q(
        npu_inst_int_data_res_2__5__2_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_5_n99), .CK(
        npu_inst_pe_1_2_5_net3995), .RN(npu_inst_pe_1_2_5_n8), .Q(
        npu_inst_int_data_res_2__5__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_5_n32), .CK(
        npu_inst_pe_1_2_5_net3995), .RN(npu_inst_pe_1_2_5_n8), .Q(
        npu_inst_int_data_res_2__5__7_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_5_n100), 
        .CK(npu_inst_pe_1_2_5_net3995), .RN(npu_inst_pe_1_2_5_n8), .Q(
        npu_inst_int_data_res_2__5__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_weight_reg_0_ ( .D(npu_inst_n93), .CK(
        npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n8), .Q(
        npu_inst_pe_1_2_5_int_q_weight_0_), .QN(npu_inst_pe_1_2_5_n27) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_weight_reg_1_ ( .D(npu_inst_n99), .CK(
        npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n8), .Q(
        npu_inst_pe_1_2_5_int_q_weight_1_), .QN(npu_inst_pe_1_2_5_n26) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_5_n112), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n8), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_5_n106), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n8), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_5_n111), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_5_n105), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_5_n110), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_5_n104), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_5_n109), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_5_n103), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_5_n108), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_5_n102), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_5_n107), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_5_n101), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_5_n86), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_5_n87), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n9), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_5_n88), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_5_n89), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_5_n90), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_5_n91), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_5_n92), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_5_n93), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_5_n94), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_5_n95), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_5_n96), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_5_n97), 
        .CK(npu_inst_pe_1_2_5_net4001), .RN(npu_inst_pe_1_2_5_n10), .Q(
        npu_inst_pe_1_2_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_5_net3995) );
  CLKGATETST_X1 npu_inst_pe_1_2_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n46), .SE(1'b0), .GCK(npu_inst_pe_1_2_5_net4001) );
  MUX2_X1 npu_inst_pe_1_2_6_U153 ( .A(npu_inst_pe_1_2_6_n31), .B(
        npu_inst_pe_1_2_6_n28), .S(npu_inst_pe_1_2_6_n7), .Z(
        npu_inst_pe_1_2_6_N93) );
  MUX2_X1 npu_inst_pe_1_2_6_U152 ( .A(npu_inst_pe_1_2_6_n30), .B(
        npu_inst_pe_1_2_6_n29), .S(npu_inst_pe_1_2_6_n5), .Z(
        npu_inst_pe_1_2_6_n31) );
  MUX2_X1 npu_inst_pe_1_2_6_U151 ( .A(npu_inst_pe_1_2_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_6_n3), .Z(
        npu_inst_pe_1_2_6_n30) );
  MUX2_X1 npu_inst_pe_1_2_6_U150 ( .A(npu_inst_pe_1_2_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_6_n3), .Z(
        npu_inst_pe_1_2_6_n29) );
  MUX2_X1 npu_inst_pe_1_2_6_U149 ( .A(npu_inst_pe_1_2_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_6_n3), .Z(
        npu_inst_pe_1_2_6_n28) );
  MUX2_X1 npu_inst_pe_1_2_6_U148 ( .A(npu_inst_pe_1_2_6_n25), .B(
        npu_inst_pe_1_2_6_n22), .S(npu_inst_pe_1_2_6_n7), .Z(
        npu_inst_pe_1_2_6_N94) );
  MUX2_X1 npu_inst_pe_1_2_6_U147 ( .A(npu_inst_pe_1_2_6_n24), .B(
        npu_inst_pe_1_2_6_n23), .S(npu_inst_pe_1_2_6_n5), .Z(
        npu_inst_pe_1_2_6_n25) );
  MUX2_X1 npu_inst_pe_1_2_6_U146 ( .A(npu_inst_pe_1_2_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_6_n3), .Z(
        npu_inst_pe_1_2_6_n24) );
  MUX2_X1 npu_inst_pe_1_2_6_U145 ( .A(npu_inst_pe_1_2_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_6_n3), .Z(
        npu_inst_pe_1_2_6_n23) );
  MUX2_X1 npu_inst_pe_1_2_6_U144 ( .A(npu_inst_pe_1_2_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_6_n3), .Z(
        npu_inst_pe_1_2_6_n22) );
  MUX2_X1 npu_inst_pe_1_2_6_U143 ( .A(npu_inst_pe_1_2_6_n21), .B(
        npu_inst_pe_1_2_6_n18), .S(npu_inst_pe_1_2_6_n7), .Z(
        npu_inst_int_data_x_2__6__1_) );
  MUX2_X1 npu_inst_pe_1_2_6_U142 ( .A(npu_inst_pe_1_2_6_n20), .B(
        npu_inst_pe_1_2_6_n19), .S(npu_inst_pe_1_2_6_n5), .Z(
        npu_inst_pe_1_2_6_n21) );
  MUX2_X1 npu_inst_pe_1_2_6_U141 ( .A(npu_inst_pe_1_2_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_6_n3), .Z(
        npu_inst_pe_1_2_6_n20) );
  MUX2_X1 npu_inst_pe_1_2_6_U140 ( .A(npu_inst_pe_1_2_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_6_n3), .Z(
        npu_inst_pe_1_2_6_n19) );
  MUX2_X1 npu_inst_pe_1_2_6_U139 ( .A(npu_inst_pe_1_2_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_6_n3), .Z(
        npu_inst_pe_1_2_6_n18) );
  MUX2_X1 npu_inst_pe_1_2_6_U138 ( .A(npu_inst_pe_1_2_6_n17), .B(
        npu_inst_pe_1_2_6_n14), .S(npu_inst_pe_1_2_6_n7), .Z(
        npu_inst_int_data_x_2__6__0_) );
  MUX2_X1 npu_inst_pe_1_2_6_U137 ( .A(npu_inst_pe_1_2_6_n16), .B(
        npu_inst_pe_1_2_6_n15), .S(npu_inst_pe_1_2_6_n5), .Z(
        npu_inst_pe_1_2_6_n17) );
  MUX2_X1 npu_inst_pe_1_2_6_U136 ( .A(npu_inst_pe_1_2_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_6_n3), .Z(
        npu_inst_pe_1_2_6_n16) );
  MUX2_X1 npu_inst_pe_1_2_6_U135 ( .A(npu_inst_pe_1_2_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_6_n3), .Z(
        npu_inst_pe_1_2_6_n15) );
  MUX2_X1 npu_inst_pe_1_2_6_U134 ( .A(npu_inst_pe_1_2_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_6_n3), .Z(
        npu_inst_pe_1_2_6_n14) );
  XOR2_X1 npu_inst_pe_1_2_6_U133 ( .A(npu_inst_pe_1_2_6_int_data_0_), .B(
        npu_inst_int_data_res_2__6__0_), .Z(npu_inst_pe_1_2_6_N73) );
  AND2_X1 npu_inst_pe_1_2_6_U132 ( .A1(npu_inst_int_data_res_2__6__0_), .A2(
        npu_inst_pe_1_2_6_int_data_0_), .ZN(npu_inst_pe_1_2_6_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_6_U131 ( .A(npu_inst_int_data_res_2__6__0_), .B(
        npu_inst_pe_1_2_6_n12), .ZN(npu_inst_pe_1_2_6_N65) );
  OR2_X1 npu_inst_pe_1_2_6_U130 ( .A1(npu_inst_pe_1_2_6_n12), .A2(
        npu_inst_int_data_res_2__6__0_), .ZN(npu_inst_pe_1_2_6_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_6_U129 ( .A(npu_inst_int_data_res_2__6__2_), .B(
        npu_inst_pe_1_2_6_add_79_carry_2_), .Z(npu_inst_pe_1_2_6_N75) );
  AND2_X1 npu_inst_pe_1_2_6_U128 ( .A1(npu_inst_pe_1_2_6_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_2__6__2_), .ZN(
        npu_inst_pe_1_2_6_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_6_U127 ( .A(npu_inst_int_data_res_2__6__3_), .B(
        npu_inst_pe_1_2_6_add_79_carry_3_), .Z(npu_inst_pe_1_2_6_N76) );
  AND2_X1 npu_inst_pe_1_2_6_U126 ( .A1(npu_inst_pe_1_2_6_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_2__6__3_), .ZN(
        npu_inst_pe_1_2_6_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_6_U125 ( .A(npu_inst_int_data_res_2__6__4_), .B(
        npu_inst_pe_1_2_6_add_79_carry_4_), .Z(npu_inst_pe_1_2_6_N77) );
  AND2_X1 npu_inst_pe_1_2_6_U124 ( .A1(npu_inst_pe_1_2_6_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_2__6__4_), .ZN(
        npu_inst_pe_1_2_6_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_6_U123 ( .A(npu_inst_int_data_res_2__6__5_), .B(
        npu_inst_pe_1_2_6_add_79_carry_5_), .Z(npu_inst_pe_1_2_6_N78) );
  AND2_X1 npu_inst_pe_1_2_6_U122 ( .A1(npu_inst_pe_1_2_6_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_2__6__5_), .ZN(
        npu_inst_pe_1_2_6_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_6_U121 ( .A(npu_inst_int_data_res_2__6__6_), .B(
        npu_inst_pe_1_2_6_add_79_carry_6_), .Z(npu_inst_pe_1_2_6_N79) );
  AND2_X1 npu_inst_pe_1_2_6_U120 ( .A1(npu_inst_pe_1_2_6_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_2__6__6_), .ZN(
        npu_inst_pe_1_2_6_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_6_U119 ( .A(npu_inst_int_data_res_2__6__7_), .B(
        npu_inst_pe_1_2_6_add_79_carry_7_), .Z(npu_inst_pe_1_2_6_N80) );
  XNOR2_X1 npu_inst_pe_1_2_6_U118 ( .A(npu_inst_pe_1_2_6_sub_77_carry_2_), .B(
        npu_inst_int_data_res_2__6__2_), .ZN(npu_inst_pe_1_2_6_N67) );
  OR2_X1 npu_inst_pe_1_2_6_U117 ( .A1(npu_inst_int_data_res_2__6__2_), .A2(
        npu_inst_pe_1_2_6_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_2_6_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_6_U116 ( .A(npu_inst_pe_1_2_6_sub_77_carry_3_), .B(
        npu_inst_int_data_res_2__6__3_), .ZN(npu_inst_pe_1_2_6_N68) );
  OR2_X1 npu_inst_pe_1_2_6_U115 ( .A1(npu_inst_int_data_res_2__6__3_), .A2(
        npu_inst_pe_1_2_6_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_2_6_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_6_U114 ( .A(npu_inst_pe_1_2_6_sub_77_carry_4_), .B(
        npu_inst_int_data_res_2__6__4_), .ZN(npu_inst_pe_1_2_6_N69) );
  OR2_X1 npu_inst_pe_1_2_6_U113 ( .A1(npu_inst_int_data_res_2__6__4_), .A2(
        npu_inst_pe_1_2_6_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_2_6_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_6_U112 ( .A(npu_inst_pe_1_2_6_sub_77_carry_5_), .B(
        npu_inst_int_data_res_2__6__5_), .ZN(npu_inst_pe_1_2_6_N70) );
  OR2_X1 npu_inst_pe_1_2_6_U111 ( .A1(npu_inst_int_data_res_2__6__5_), .A2(
        npu_inst_pe_1_2_6_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_2_6_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_6_U110 ( .A(npu_inst_pe_1_2_6_sub_77_carry_6_), .B(
        npu_inst_int_data_res_2__6__6_), .ZN(npu_inst_pe_1_2_6_N71) );
  OR2_X1 npu_inst_pe_1_2_6_U109 ( .A1(npu_inst_int_data_res_2__6__6_), .A2(
        npu_inst_pe_1_2_6_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_2_6_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_6_U108 ( .A(npu_inst_int_data_res_2__6__7_), .B(
        npu_inst_pe_1_2_6_sub_77_carry_7_), .ZN(npu_inst_pe_1_2_6_N72) );
  INV_X1 npu_inst_pe_1_2_6_U107 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_2_6_n6)
         );
  INV_X1 npu_inst_pe_1_2_6_U106 ( .A(npu_inst_pe_1_2_6_n6), .ZN(
        npu_inst_pe_1_2_6_n5) );
  INV_X1 npu_inst_pe_1_2_6_U105 ( .A(npu_inst_n39), .ZN(npu_inst_pe_1_2_6_n2)
         );
  AOI22_X1 npu_inst_pe_1_2_6_U104 ( .A1(npu_inst_int_data_y_3__6__0_), .A2(
        npu_inst_pe_1_2_6_n58), .B1(npu_inst_pe_1_2_6_n118), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_6_n57) );
  INV_X1 npu_inst_pe_1_2_6_U103 ( .A(npu_inst_pe_1_2_6_n57), .ZN(
        npu_inst_pe_1_2_6_n107) );
  AOI22_X1 npu_inst_pe_1_2_6_U102 ( .A1(npu_inst_int_data_y_3__6__0_), .A2(
        npu_inst_pe_1_2_6_n54), .B1(npu_inst_pe_1_2_6_n117), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_6_n53) );
  INV_X1 npu_inst_pe_1_2_6_U99 ( .A(npu_inst_pe_1_2_6_n53), .ZN(
        npu_inst_pe_1_2_6_n108) );
  AOI22_X1 npu_inst_pe_1_2_6_U98 ( .A1(npu_inst_int_data_y_3__6__0_), .A2(
        npu_inst_pe_1_2_6_n50), .B1(npu_inst_pe_1_2_6_n116), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_6_n49) );
  INV_X1 npu_inst_pe_1_2_6_U97 ( .A(npu_inst_pe_1_2_6_n49), .ZN(
        npu_inst_pe_1_2_6_n109) );
  AOI22_X1 npu_inst_pe_1_2_6_U96 ( .A1(npu_inst_int_data_y_3__6__0_), .A2(
        npu_inst_pe_1_2_6_n46), .B1(npu_inst_pe_1_2_6_n115), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_6_n45) );
  INV_X1 npu_inst_pe_1_2_6_U95 ( .A(npu_inst_pe_1_2_6_n45), .ZN(
        npu_inst_pe_1_2_6_n110) );
  AOI22_X1 npu_inst_pe_1_2_6_U94 ( .A1(npu_inst_int_data_y_3__6__0_), .A2(
        npu_inst_pe_1_2_6_n42), .B1(npu_inst_pe_1_2_6_n114), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_6_n41) );
  INV_X1 npu_inst_pe_1_2_6_U93 ( .A(npu_inst_pe_1_2_6_n41), .ZN(
        npu_inst_pe_1_2_6_n111) );
  AOI22_X1 npu_inst_pe_1_2_6_U92 ( .A1(npu_inst_int_data_y_3__6__1_), .A2(
        npu_inst_pe_1_2_6_n58), .B1(npu_inst_pe_1_2_6_n118), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_6_n59) );
  INV_X1 npu_inst_pe_1_2_6_U91 ( .A(npu_inst_pe_1_2_6_n59), .ZN(
        npu_inst_pe_1_2_6_n101) );
  AOI22_X1 npu_inst_pe_1_2_6_U90 ( .A1(npu_inst_int_data_y_3__6__1_), .A2(
        npu_inst_pe_1_2_6_n54), .B1(npu_inst_pe_1_2_6_n117), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_6_n55) );
  INV_X1 npu_inst_pe_1_2_6_U89 ( .A(npu_inst_pe_1_2_6_n55), .ZN(
        npu_inst_pe_1_2_6_n102) );
  AOI22_X1 npu_inst_pe_1_2_6_U88 ( .A1(npu_inst_int_data_y_3__6__1_), .A2(
        npu_inst_pe_1_2_6_n50), .B1(npu_inst_pe_1_2_6_n116), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_6_n51) );
  INV_X1 npu_inst_pe_1_2_6_U87 ( .A(npu_inst_pe_1_2_6_n51), .ZN(
        npu_inst_pe_1_2_6_n103) );
  AOI22_X1 npu_inst_pe_1_2_6_U86 ( .A1(npu_inst_int_data_y_3__6__1_), .A2(
        npu_inst_pe_1_2_6_n46), .B1(npu_inst_pe_1_2_6_n115), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_6_n47) );
  INV_X1 npu_inst_pe_1_2_6_U85 ( .A(npu_inst_pe_1_2_6_n47), .ZN(
        npu_inst_pe_1_2_6_n104) );
  AOI22_X1 npu_inst_pe_1_2_6_U84 ( .A1(npu_inst_int_data_y_3__6__1_), .A2(
        npu_inst_pe_1_2_6_n42), .B1(npu_inst_pe_1_2_6_n114), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_6_n43) );
  INV_X1 npu_inst_pe_1_2_6_U83 ( .A(npu_inst_pe_1_2_6_n43), .ZN(
        npu_inst_pe_1_2_6_n105) );
  AOI22_X1 npu_inst_pe_1_2_6_U82 ( .A1(npu_inst_pe_1_2_6_n38), .A2(
        npu_inst_int_data_y_3__6__1_), .B1(npu_inst_pe_1_2_6_n113), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_6_n39) );
  INV_X1 npu_inst_pe_1_2_6_U81 ( .A(npu_inst_pe_1_2_6_n39), .ZN(
        npu_inst_pe_1_2_6_n106) );
  AND2_X1 npu_inst_pe_1_2_6_U80 ( .A1(npu_inst_pe_1_2_6_N93), .A2(npu_inst_n39), .ZN(npu_inst_int_data_y_2__6__0_) );
  NAND2_X1 npu_inst_pe_1_2_6_U79 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_6_n60), .ZN(npu_inst_pe_1_2_6_n74) );
  OAI21_X1 npu_inst_pe_1_2_6_U78 ( .B1(npu_inst_pe_1_2_6_n63), .B2(
        npu_inst_pe_1_2_6_n60), .A(npu_inst_pe_1_2_6_n74), .ZN(
        npu_inst_pe_1_2_6_n97) );
  NAND2_X1 npu_inst_pe_1_2_6_U77 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_6_n60), .ZN(npu_inst_pe_1_2_6_n73) );
  OAI21_X1 npu_inst_pe_1_2_6_U76 ( .B1(npu_inst_pe_1_2_6_n61), .B2(
        npu_inst_pe_1_2_6_n60), .A(npu_inst_pe_1_2_6_n73), .ZN(
        npu_inst_pe_1_2_6_n96) );
  NAND2_X1 npu_inst_pe_1_2_6_U75 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_6_n56), .ZN(npu_inst_pe_1_2_6_n72) );
  OAI21_X1 npu_inst_pe_1_2_6_U74 ( .B1(npu_inst_pe_1_2_6_n63), .B2(
        npu_inst_pe_1_2_6_n56), .A(npu_inst_pe_1_2_6_n72), .ZN(
        npu_inst_pe_1_2_6_n95) );
  NAND2_X1 npu_inst_pe_1_2_6_U73 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_6_n56), .ZN(npu_inst_pe_1_2_6_n71) );
  OAI21_X1 npu_inst_pe_1_2_6_U72 ( .B1(npu_inst_pe_1_2_6_n61), .B2(
        npu_inst_pe_1_2_6_n56), .A(npu_inst_pe_1_2_6_n71), .ZN(
        npu_inst_pe_1_2_6_n94) );
  NAND2_X1 npu_inst_pe_1_2_6_U71 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_6_n52), .ZN(npu_inst_pe_1_2_6_n70) );
  OAI21_X1 npu_inst_pe_1_2_6_U70 ( .B1(npu_inst_pe_1_2_6_n63), .B2(
        npu_inst_pe_1_2_6_n52), .A(npu_inst_pe_1_2_6_n70), .ZN(
        npu_inst_pe_1_2_6_n93) );
  NAND2_X1 npu_inst_pe_1_2_6_U69 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_6_n52), .ZN(npu_inst_pe_1_2_6_n69) );
  OAI21_X1 npu_inst_pe_1_2_6_U68 ( .B1(npu_inst_pe_1_2_6_n61), .B2(
        npu_inst_pe_1_2_6_n52), .A(npu_inst_pe_1_2_6_n69), .ZN(
        npu_inst_pe_1_2_6_n92) );
  NAND2_X1 npu_inst_pe_1_2_6_U67 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_6_n48), .ZN(npu_inst_pe_1_2_6_n68) );
  OAI21_X1 npu_inst_pe_1_2_6_U66 ( .B1(npu_inst_pe_1_2_6_n63), .B2(
        npu_inst_pe_1_2_6_n48), .A(npu_inst_pe_1_2_6_n68), .ZN(
        npu_inst_pe_1_2_6_n91) );
  NAND2_X1 npu_inst_pe_1_2_6_U65 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_6_n48), .ZN(npu_inst_pe_1_2_6_n67) );
  OAI21_X1 npu_inst_pe_1_2_6_U64 ( .B1(npu_inst_pe_1_2_6_n61), .B2(
        npu_inst_pe_1_2_6_n48), .A(npu_inst_pe_1_2_6_n67), .ZN(
        npu_inst_pe_1_2_6_n90) );
  NAND2_X1 npu_inst_pe_1_2_6_U63 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_6_n44), .ZN(npu_inst_pe_1_2_6_n66) );
  OAI21_X1 npu_inst_pe_1_2_6_U62 ( .B1(npu_inst_pe_1_2_6_n63), .B2(
        npu_inst_pe_1_2_6_n44), .A(npu_inst_pe_1_2_6_n66), .ZN(
        npu_inst_pe_1_2_6_n89) );
  NAND2_X1 npu_inst_pe_1_2_6_U61 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_6_n44), .ZN(npu_inst_pe_1_2_6_n65) );
  OAI21_X1 npu_inst_pe_1_2_6_U60 ( .B1(npu_inst_pe_1_2_6_n61), .B2(
        npu_inst_pe_1_2_6_n44), .A(npu_inst_pe_1_2_6_n65), .ZN(
        npu_inst_pe_1_2_6_n88) );
  NAND2_X1 npu_inst_pe_1_2_6_U59 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_6_n40), .ZN(npu_inst_pe_1_2_6_n64) );
  OAI21_X1 npu_inst_pe_1_2_6_U58 ( .B1(npu_inst_pe_1_2_6_n63), .B2(
        npu_inst_pe_1_2_6_n40), .A(npu_inst_pe_1_2_6_n64), .ZN(
        npu_inst_pe_1_2_6_n87) );
  NAND2_X1 npu_inst_pe_1_2_6_U57 ( .A1(npu_inst_pe_1_2_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_6_n40), .ZN(npu_inst_pe_1_2_6_n62) );
  OAI21_X1 npu_inst_pe_1_2_6_U56 ( .B1(npu_inst_pe_1_2_6_n61), .B2(
        npu_inst_pe_1_2_6_n40), .A(npu_inst_pe_1_2_6_n62), .ZN(
        npu_inst_pe_1_2_6_n86) );
  AOI22_X1 npu_inst_pe_1_2_6_U55 ( .A1(npu_inst_pe_1_2_6_n38), .A2(
        npu_inst_int_data_y_3__6__0_), .B1(npu_inst_pe_1_2_6_n113), .B2(
        npu_inst_pe_1_2_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_6_n37) );
  INV_X1 npu_inst_pe_1_2_6_U54 ( .A(npu_inst_pe_1_2_6_n37), .ZN(
        npu_inst_pe_1_2_6_n112) );
  AND2_X1 npu_inst_pe_1_2_6_U53 ( .A1(npu_inst_n39), .A2(npu_inst_pe_1_2_6_N94), .ZN(npu_inst_int_data_y_2__6__1_) );
  AOI222_X1 npu_inst_pe_1_2_6_U52 ( .A1(npu_inst_int_data_res_3__6__0_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N73), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N65), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n84) );
  INV_X1 npu_inst_pe_1_2_6_U51 ( .A(npu_inst_pe_1_2_6_n84), .ZN(
        npu_inst_pe_1_2_6_n100) );
  AOI222_X1 npu_inst_pe_1_2_6_U50 ( .A1(npu_inst_pe_1_2_6_n1), .A2(
        npu_inst_int_data_res_3__6__7_), .B1(npu_inst_pe_1_2_6_N80), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N72), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n75) );
  INV_X1 npu_inst_pe_1_2_6_U49 ( .A(npu_inst_pe_1_2_6_n75), .ZN(
        npu_inst_pe_1_2_6_n32) );
  AOI222_X1 npu_inst_pe_1_2_6_U48 ( .A1(npu_inst_int_data_res_3__6__1_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N74), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N66), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n83) );
  INV_X1 npu_inst_pe_1_2_6_U47 ( .A(npu_inst_pe_1_2_6_n83), .ZN(
        npu_inst_pe_1_2_6_n99) );
  AOI222_X1 npu_inst_pe_1_2_6_U46 ( .A1(npu_inst_int_data_res_3__6__3_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N76), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N68), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n81) );
  INV_X1 npu_inst_pe_1_2_6_U45 ( .A(npu_inst_pe_1_2_6_n81), .ZN(
        npu_inst_pe_1_2_6_n36) );
  AOI222_X1 npu_inst_pe_1_2_6_U44 ( .A1(npu_inst_int_data_res_3__6__4_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N77), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N69), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n80) );
  INV_X1 npu_inst_pe_1_2_6_U43 ( .A(npu_inst_pe_1_2_6_n80), .ZN(
        npu_inst_pe_1_2_6_n35) );
  AOI222_X1 npu_inst_pe_1_2_6_U42 ( .A1(npu_inst_int_data_res_3__6__5_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N78), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N70), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n79) );
  INV_X1 npu_inst_pe_1_2_6_U41 ( .A(npu_inst_pe_1_2_6_n79), .ZN(
        npu_inst_pe_1_2_6_n34) );
  AOI222_X1 npu_inst_pe_1_2_6_U40 ( .A1(npu_inst_int_data_res_3__6__6_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N79), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N71), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n78) );
  INV_X1 npu_inst_pe_1_2_6_U39 ( .A(npu_inst_pe_1_2_6_n78), .ZN(
        npu_inst_pe_1_2_6_n33) );
  AND2_X1 npu_inst_pe_1_2_6_U38 ( .A1(npu_inst_int_data_x_2__6__1_), .A2(
        npu_inst_pe_1_2_6_int_q_weight_1_), .ZN(npu_inst_pe_1_2_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_6_U37 ( .A1(npu_inst_int_data_x_2__6__0_), .A2(
        npu_inst_pe_1_2_6_int_q_weight_1_), .ZN(npu_inst_pe_1_2_6_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_2_6_U36 ( .A(npu_inst_pe_1_2_6_int_data_1_), .ZN(
        npu_inst_pe_1_2_6_n13) );
  NOR3_X1 npu_inst_pe_1_2_6_U35 ( .A1(npu_inst_pe_1_2_6_n26), .A2(npu_inst_n39), .A3(npu_inst_int_ckg[41]), .ZN(npu_inst_pe_1_2_6_n85) );
  OR2_X1 npu_inst_pe_1_2_6_U34 ( .A1(npu_inst_pe_1_2_6_n85), .A2(
        npu_inst_pe_1_2_6_n1), .ZN(npu_inst_pe_1_2_6_N84) );
  AOI222_X1 npu_inst_pe_1_2_6_U33 ( .A1(npu_inst_int_data_res_3__6__2_), .A2(
        npu_inst_pe_1_2_6_n1), .B1(npu_inst_pe_1_2_6_N75), .B2(
        npu_inst_pe_1_2_6_n76), .C1(npu_inst_pe_1_2_6_N67), .C2(
        npu_inst_pe_1_2_6_n77), .ZN(npu_inst_pe_1_2_6_n82) );
  INV_X1 npu_inst_pe_1_2_6_U32 ( .A(npu_inst_pe_1_2_6_n82), .ZN(
        npu_inst_pe_1_2_6_n98) );
  AOI22_X1 npu_inst_pe_1_2_6_U31 ( .A1(npu_inst_n39), .A2(
        npu_inst_int_data_y_3__6__1_), .B1(npu_inst_pe_1_2_6_n2), .B2(
        npu_inst_int_data_x_2__7__1_), .ZN(npu_inst_pe_1_2_6_n63) );
  AOI22_X1 npu_inst_pe_1_2_6_U30 ( .A1(npu_inst_n39), .A2(
        npu_inst_int_data_y_3__6__0_), .B1(npu_inst_pe_1_2_6_n2), .B2(
        npu_inst_int_data_x_2__7__0_), .ZN(npu_inst_pe_1_2_6_n61) );
  INV_X1 npu_inst_pe_1_2_6_U29 ( .A(npu_inst_pe_1_2_6_int_data_0_), .ZN(
        npu_inst_pe_1_2_6_n12) );
  INV_X1 npu_inst_pe_1_2_6_U28 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_2_6_n4)
         );
  OR3_X1 npu_inst_pe_1_2_6_U27 ( .A1(npu_inst_pe_1_2_6_n5), .A2(
        npu_inst_pe_1_2_6_n7), .A3(npu_inst_pe_1_2_6_n4), .ZN(
        npu_inst_pe_1_2_6_n56) );
  OR3_X1 npu_inst_pe_1_2_6_U26 ( .A1(npu_inst_pe_1_2_6_n4), .A2(
        npu_inst_pe_1_2_6_n7), .A3(npu_inst_pe_1_2_6_n6), .ZN(
        npu_inst_pe_1_2_6_n48) );
  INV_X1 npu_inst_pe_1_2_6_U25 ( .A(npu_inst_pe_1_2_6_n4), .ZN(
        npu_inst_pe_1_2_6_n3) );
  OR3_X1 npu_inst_pe_1_2_6_U24 ( .A1(npu_inst_pe_1_2_6_n3), .A2(
        npu_inst_pe_1_2_6_n7), .A3(npu_inst_pe_1_2_6_n6), .ZN(
        npu_inst_pe_1_2_6_n52) );
  OR3_X1 npu_inst_pe_1_2_6_U23 ( .A1(npu_inst_pe_1_2_6_n5), .A2(
        npu_inst_pe_1_2_6_n7), .A3(npu_inst_pe_1_2_6_n3), .ZN(
        npu_inst_pe_1_2_6_n60) );
  BUF_X1 npu_inst_pe_1_2_6_U22 ( .A(npu_inst_n24), .Z(npu_inst_pe_1_2_6_n1) );
  NOR2_X1 npu_inst_pe_1_2_6_U21 ( .A1(npu_inst_pe_1_2_6_n60), .A2(
        npu_inst_pe_1_2_6_n2), .ZN(npu_inst_pe_1_2_6_n58) );
  NOR2_X1 npu_inst_pe_1_2_6_U20 ( .A1(npu_inst_pe_1_2_6_n56), .A2(
        npu_inst_pe_1_2_6_n2), .ZN(npu_inst_pe_1_2_6_n54) );
  NOR2_X1 npu_inst_pe_1_2_6_U19 ( .A1(npu_inst_pe_1_2_6_n52), .A2(
        npu_inst_pe_1_2_6_n2), .ZN(npu_inst_pe_1_2_6_n50) );
  NOR2_X1 npu_inst_pe_1_2_6_U18 ( .A1(npu_inst_pe_1_2_6_n48), .A2(
        npu_inst_pe_1_2_6_n2), .ZN(npu_inst_pe_1_2_6_n46) );
  NOR2_X1 npu_inst_pe_1_2_6_U17 ( .A1(npu_inst_pe_1_2_6_n40), .A2(
        npu_inst_pe_1_2_6_n2), .ZN(npu_inst_pe_1_2_6_n38) );
  NOR2_X1 npu_inst_pe_1_2_6_U16 ( .A1(npu_inst_pe_1_2_6_n44), .A2(
        npu_inst_pe_1_2_6_n2), .ZN(npu_inst_pe_1_2_6_n42) );
  BUF_X1 npu_inst_pe_1_2_6_U15 ( .A(npu_inst_n84), .Z(npu_inst_pe_1_2_6_n7) );
  INV_X1 npu_inst_pe_1_2_6_U14 ( .A(npu_inst_n107), .ZN(npu_inst_pe_1_2_6_n11)
         );
  INV_X1 npu_inst_pe_1_2_6_U13 ( .A(npu_inst_pe_1_2_6_n38), .ZN(
        npu_inst_pe_1_2_6_n113) );
  INV_X1 npu_inst_pe_1_2_6_U12 ( .A(npu_inst_pe_1_2_6_n58), .ZN(
        npu_inst_pe_1_2_6_n118) );
  INV_X1 npu_inst_pe_1_2_6_U11 ( .A(npu_inst_pe_1_2_6_n54), .ZN(
        npu_inst_pe_1_2_6_n117) );
  INV_X1 npu_inst_pe_1_2_6_U10 ( .A(npu_inst_pe_1_2_6_n50), .ZN(
        npu_inst_pe_1_2_6_n116) );
  INV_X1 npu_inst_pe_1_2_6_U9 ( .A(npu_inst_pe_1_2_6_n46), .ZN(
        npu_inst_pe_1_2_6_n115) );
  INV_X1 npu_inst_pe_1_2_6_U8 ( .A(npu_inst_pe_1_2_6_n42), .ZN(
        npu_inst_pe_1_2_6_n114) );
  BUF_X1 npu_inst_pe_1_2_6_U7 ( .A(npu_inst_pe_1_2_6_n11), .Z(
        npu_inst_pe_1_2_6_n10) );
  BUF_X1 npu_inst_pe_1_2_6_U6 ( .A(npu_inst_pe_1_2_6_n11), .Z(
        npu_inst_pe_1_2_6_n9) );
  BUF_X1 npu_inst_pe_1_2_6_U5 ( .A(npu_inst_pe_1_2_6_n11), .Z(
        npu_inst_pe_1_2_6_n8) );
  NOR2_X1 npu_inst_pe_1_2_6_U4 ( .A1(npu_inst_pe_1_2_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_6_n1), .ZN(npu_inst_pe_1_2_6_n76) );
  NOR2_X1 npu_inst_pe_1_2_6_U3 ( .A1(npu_inst_pe_1_2_6_n27), .A2(
        npu_inst_pe_1_2_6_n1), .ZN(npu_inst_pe_1_2_6_n77) );
  FA_X1 npu_inst_pe_1_2_6_sub_77_U2_1 ( .A(npu_inst_int_data_res_2__6__1_), 
        .B(npu_inst_pe_1_2_6_n13), .CI(npu_inst_pe_1_2_6_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_2_6_sub_77_carry_2_), .S(npu_inst_pe_1_2_6_N66) );
  FA_X1 npu_inst_pe_1_2_6_add_79_U1_1 ( .A(npu_inst_int_data_res_2__6__1_), 
        .B(npu_inst_pe_1_2_6_int_data_1_), .CI(
        npu_inst_pe_1_2_6_add_79_carry_1_), .CO(
        npu_inst_pe_1_2_6_add_79_carry_2_), .S(npu_inst_pe_1_2_6_N74) );
  NAND3_X1 npu_inst_pe_1_2_6_U101 ( .A1(npu_inst_pe_1_2_6_n4), .A2(
        npu_inst_pe_1_2_6_n6), .A3(npu_inst_pe_1_2_6_n7), .ZN(
        npu_inst_pe_1_2_6_n44) );
  NAND3_X1 npu_inst_pe_1_2_6_U100 ( .A1(npu_inst_pe_1_2_6_n3), .A2(
        npu_inst_pe_1_2_6_n6), .A3(npu_inst_pe_1_2_6_n7), .ZN(
        npu_inst_pe_1_2_6_n40) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_6_n33), .CK(
        npu_inst_pe_1_2_6_net3972), .RN(npu_inst_pe_1_2_6_n8), .Q(
        npu_inst_int_data_res_2__6__6_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_6_n34), .CK(
        npu_inst_pe_1_2_6_net3972), .RN(npu_inst_pe_1_2_6_n8), .Q(
        npu_inst_int_data_res_2__6__5_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_6_n35), .CK(
        npu_inst_pe_1_2_6_net3972), .RN(npu_inst_pe_1_2_6_n8), .Q(
        npu_inst_int_data_res_2__6__4_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_6_n36), .CK(
        npu_inst_pe_1_2_6_net3972), .RN(npu_inst_pe_1_2_6_n8), .Q(
        npu_inst_int_data_res_2__6__3_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_6_n98), .CK(
        npu_inst_pe_1_2_6_net3972), .RN(npu_inst_pe_1_2_6_n8), .Q(
        npu_inst_int_data_res_2__6__2_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_6_n99), .CK(
        npu_inst_pe_1_2_6_net3972), .RN(npu_inst_pe_1_2_6_n8), .Q(
        npu_inst_int_data_res_2__6__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_6_n32), .CK(
        npu_inst_pe_1_2_6_net3972), .RN(npu_inst_pe_1_2_6_n8), .Q(
        npu_inst_int_data_res_2__6__7_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_6_n100), 
        .CK(npu_inst_pe_1_2_6_net3972), .RN(npu_inst_pe_1_2_6_n8), .Q(
        npu_inst_int_data_res_2__6__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_weight_reg_0_ ( .D(npu_inst_n93), .CK(
        npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n8), .Q(
        npu_inst_pe_1_2_6_int_q_weight_0_), .QN(npu_inst_pe_1_2_6_n27) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_weight_reg_1_ ( .D(npu_inst_n99), .CK(
        npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n8), .Q(
        npu_inst_pe_1_2_6_int_q_weight_1_), .QN(npu_inst_pe_1_2_6_n26) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_6_n112), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n8), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_6_n106), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n8), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_6_n111), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_6_n105), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_6_n110), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_6_n104), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_6_n109), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_6_n103), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_6_n108), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_6_n102), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_6_n107), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_6_n101), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_6_n86), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_6_n87), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n9), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_6_n88), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_6_n89), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_6_n90), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_6_n91), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_6_n92), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_6_n93), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_6_n94), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_6_n95), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_6_n96), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_6_n97), 
        .CK(npu_inst_pe_1_2_6_net3978), .RN(npu_inst_pe_1_2_6_n10), .Q(
        npu_inst_pe_1_2_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_6_net3972) );
  CLKGATETST_X1 npu_inst_pe_1_2_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n46), .SE(1'b0), .GCK(npu_inst_pe_1_2_6_net3978) );
  MUX2_X1 npu_inst_pe_1_2_7_U153 ( .A(npu_inst_pe_1_2_7_n31), .B(
        npu_inst_pe_1_2_7_n28), .S(npu_inst_pe_1_2_7_n7), .Z(
        npu_inst_pe_1_2_7_N93) );
  MUX2_X1 npu_inst_pe_1_2_7_U152 ( .A(npu_inst_pe_1_2_7_n30), .B(
        npu_inst_pe_1_2_7_n29), .S(npu_inst_pe_1_2_7_n5), .Z(
        npu_inst_pe_1_2_7_n31) );
  MUX2_X1 npu_inst_pe_1_2_7_U151 ( .A(npu_inst_pe_1_2_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_2_7_n3), .Z(
        npu_inst_pe_1_2_7_n30) );
  MUX2_X1 npu_inst_pe_1_2_7_U150 ( .A(npu_inst_pe_1_2_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_2_7_n3), .Z(
        npu_inst_pe_1_2_7_n29) );
  MUX2_X1 npu_inst_pe_1_2_7_U149 ( .A(npu_inst_pe_1_2_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_2_7_n3), .Z(
        npu_inst_pe_1_2_7_n28) );
  MUX2_X1 npu_inst_pe_1_2_7_U148 ( .A(npu_inst_pe_1_2_7_n25), .B(
        npu_inst_pe_1_2_7_n22), .S(npu_inst_pe_1_2_7_n7), .Z(
        npu_inst_pe_1_2_7_N94) );
  MUX2_X1 npu_inst_pe_1_2_7_U147 ( .A(npu_inst_pe_1_2_7_n24), .B(
        npu_inst_pe_1_2_7_n23), .S(npu_inst_pe_1_2_7_n5), .Z(
        npu_inst_pe_1_2_7_n25) );
  MUX2_X1 npu_inst_pe_1_2_7_U146 ( .A(npu_inst_pe_1_2_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_2_7_n3), .Z(
        npu_inst_pe_1_2_7_n24) );
  MUX2_X1 npu_inst_pe_1_2_7_U145 ( .A(npu_inst_pe_1_2_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_2_7_n3), .Z(
        npu_inst_pe_1_2_7_n23) );
  MUX2_X1 npu_inst_pe_1_2_7_U144 ( .A(npu_inst_pe_1_2_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_2_7_n3), .Z(
        npu_inst_pe_1_2_7_n22) );
  MUX2_X1 npu_inst_pe_1_2_7_U143 ( .A(npu_inst_pe_1_2_7_n21), .B(
        npu_inst_pe_1_2_7_n18), .S(npu_inst_pe_1_2_7_n7), .Z(
        npu_inst_int_data_x_2__7__1_) );
  MUX2_X1 npu_inst_pe_1_2_7_U142 ( .A(npu_inst_pe_1_2_7_n20), .B(
        npu_inst_pe_1_2_7_n19), .S(npu_inst_pe_1_2_7_n5), .Z(
        npu_inst_pe_1_2_7_n21) );
  MUX2_X1 npu_inst_pe_1_2_7_U141 ( .A(npu_inst_pe_1_2_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_2_7_n3), .Z(
        npu_inst_pe_1_2_7_n20) );
  MUX2_X1 npu_inst_pe_1_2_7_U140 ( .A(npu_inst_pe_1_2_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_2_7_n3), .Z(
        npu_inst_pe_1_2_7_n19) );
  MUX2_X1 npu_inst_pe_1_2_7_U139 ( .A(npu_inst_pe_1_2_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_2_7_n3), .Z(
        npu_inst_pe_1_2_7_n18) );
  MUX2_X1 npu_inst_pe_1_2_7_U138 ( .A(npu_inst_pe_1_2_7_n17), .B(
        npu_inst_pe_1_2_7_n14), .S(npu_inst_pe_1_2_7_n7), .Z(
        npu_inst_int_data_x_2__7__0_) );
  MUX2_X1 npu_inst_pe_1_2_7_U137 ( .A(npu_inst_pe_1_2_7_n16), .B(
        npu_inst_pe_1_2_7_n15), .S(npu_inst_pe_1_2_7_n5), .Z(
        npu_inst_pe_1_2_7_n17) );
  MUX2_X1 npu_inst_pe_1_2_7_U136 ( .A(npu_inst_pe_1_2_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_2_7_n3), .Z(
        npu_inst_pe_1_2_7_n16) );
  MUX2_X1 npu_inst_pe_1_2_7_U135 ( .A(npu_inst_pe_1_2_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_2_7_n3), .Z(
        npu_inst_pe_1_2_7_n15) );
  MUX2_X1 npu_inst_pe_1_2_7_U134 ( .A(npu_inst_pe_1_2_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_2_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_2_7_n3), .Z(
        npu_inst_pe_1_2_7_n14) );
  XOR2_X1 npu_inst_pe_1_2_7_U133 ( .A(npu_inst_pe_1_2_7_int_data_0_), .B(
        npu_inst_int_data_res_2__7__0_), .Z(npu_inst_pe_1_2_7_N73) );
  AND2_X1 npu_inst_pe_1_2_7_U132 ( .A1(npu_inst_int_data_res_2__7__0_), .A2(
        npu_inst_pe_1_2_7_int_data_0_), .ZN(npu_inst_pe_1_2_7_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_2_7_U131 ( .A(npu_inst_int_data_res_2__7__0_), .B(
        npu_inst_pe_1_2_7_n12), .ZN(npu_inst_pe_1_2_7_N65) );
  OR2_X1 npu_inst_pe_1_2_7_U130 ( .A1(npu_inst_pe_1_2_7_n12), .A2(
        npu_inst_int_data_res_2__7__0_), .ZN(npu_inst_pe_1_2_7_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_2_7_U129 ( .A(npu_inst_int_data_res_2__7__2_), .B(
        npu_inst_pe_1_2_7_add_79_carry_2_), .Z(npu_inst_pe_1_2_7_N75) );
  AND2_X1 npu_inst_pe_1_2_7_U128 ( .A1(npu_inst_pe_1_2_7_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_2__7__2_), .ZN(
        npu_inst_pe_1_2_7_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_2_7_U127 ( .A(npu_inst_int_data_res_2__7__3_), .B(
        npu_inst_pe_1_2_7_add_79_carry_3_), .Z(npu_inst_pe_1_2_7_N76) );
  AND2_X1 npu_inst_pe_1_2_7_U126 ( .A1(npu_inst_pe_1_2_7_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_2__7__3_), .ZN(
        npu_inst_pe_1_2_7_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_2_7_U125 ( .A(npu_inst_int_data_res_2__7__4_), .B(
        npu_inst_pe_1_2_7_add_79_carry_4_), .Z(npu_inst_pe_1_2_7_N77) );
  AND2_X1 npu_inst_pe_1_2_7_U124 ( .A1(npu_inst_pe_1_2_7_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_2__7__4_), .ZN(
        npu_inst_pe_1_2_7_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_2_7_U123 ( .A(npu_inst_int_data_res_2__7__5_), .B(
        npu_inst_pe_1_2_7_add_79_carry_5_), .Z(npu_inst_pe_1_2_7_N78) );
  AND2_X1 npu_inst_pe_1_2_7_U122 ( .A1(npu_inst_pe_1_2_7_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_2__7__5_), .ZN(
        npu_inst_pe_1_2_7_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_2_7_U121 ( .A(npu_inst_int_data_res_2__7__6_), .B(
        npu_inst_pe_1_2_7_add_79_carry_6_), .Z(npu_inst_pe_1_2_7_N79) );
  AND2_X1 npu_inst_pe_1_2_7_U120 ( .A1(npu_inst_pe_1_2_7_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_2__7__6_), .ZN(
        npu_inst_pe_1_2_7_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_2_7_U119 ( .A(npu_inst_int_data_res_2__7__7_), .B(
        npu_inst_pe_1_2_7_add_79_carry_7_), .Z(npu_inst_pe_1_2_7_N80) );
  XNOR2_X1 npu_inst_pe_1_2_7_U118 ( .A(npu_inst_pe_1_2_7_sub_77_carry_2_), .B(
        npu_inst_int_data_res_2__7__2_), .ZN(npu_inst_pe_1_2_7_N67) );
  OR2_X1 npu_inst_pe_1_2_7_U117 ( .A1(npu_inst_int_data_res_2__7__2_), .A2(
        npu_inst_pe_1_2_7_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_2_7_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_2_7_U116 ( .A(npu_inst_pe_1_2_7_sub_77_carry_3_), .B(
        npu_inst_int_data_res_2__7__3_), .ZN(npu_inst_pe_1_2_7_N68) );
  OR2_X1 npu_inst_pe_1_2_7_U115 ( .A1(npu_inst_int_data_res_2__7__3_), .A2(
        npu_inst_pe_1_2_7_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_2_7_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_2_7_U114 ( .A(npu_inst_pe_1_2_7_sub_77_carry_4_), .B(
        npu_inst_int_data_res_2__7__4_), .ZN(npu_inst_pe_1_2_7_N69) );
  OR2_X1 npu_inst_pe_1_2_7_U113 ( .A1(npu_inst_int_data_res_2__7__4_), .A2(
        npu_inst_pe_1_2_7_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_2_7_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_2_7_U112 ( .A(npu_inst_pe_1_2_7_sub_77_carry_5_), .B(
        npu_inst_int_data_res_2__7__5_), .ZN(npu_inst_pe_1_2_7_N70) );
  OR2_X1 npu_inst_pe_1_2_7_U111 ( .A1(npu_inst_int_data_res_2__7__5_), .A2(
        npu_inst_pe_1_2_7_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_2_7_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_2_7_U110 ( .A(npu_inst_pe_1_2_7_sub_77_carry_6_), .B(
        npu_inst_int_data_res_2__7__6_), .ZN(npu_inst_pe_1_2_7_N71) );
  OR2_X1 npu_inst_pe_1_2_7_U109 ( .A1(npu_inst_int_data_res_2__7__6_), .A2(
        npu_inst_pe_1_2_7_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_2_7_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_2_7_U108 ( .A(npu_inst_int_data_res_2__7__7_), .B(
        npu_inst_pe_1_2_7_sub_77_carry_7_), .ZN(npu_inst_pe_1_2_7_N72) );
  INV_X1 npu_inst_pe_1_2_7_U107 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_2_7_n6)
         );
  INV_X1 npu_inst_pe_1_2_7_U106 ( .A(npu_inst_pe_1_2_7_n6), .ZN(
        npu_inst_pe_1_2_7_n5) );
  INV_X1 npu_inst_pe_1_2_7_U105 ( .A(npu_inst_n39), .ZN(npu_inst_pe_1_2_7_n2)
         );
  AOI22_X1 npu_inst_pe_1_2_7_U104 ( .A1(npu_inst_int_data_y_3__7__0_), .A2(
        npu_inst_pe_1_2_7_n58), .B1(npu_inst_pe_1_2_7_n118), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_2_7_n57) );
  INV_X1 npu_inst_pe_1_2_7_U103 ( .A(npu_inst_pe_1_2_7_n57), .ZN(
        npu_inst_pe_1_2_7_n107) );
  AOI22_X1 npu_inst_pe_1_2_7_U102 ( .A1(npu_inst_int_data_y_3__7__0_), .A2(
        npu_inst_pe_1_2_7_n54), .B1(npu_inst_pe_1_2_7_n117), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_2_7_n53) );
  INV_X1 npu_inst_pe_1_2_7_U99 ( .A(npu_inst_pe_1_2_7_n53), .ZN(
        npu_inst_pe_1_2_7_n108) );
  AOI22_X1 npu_inst_pe_1_2_7_U98 ( .A1(npu_inst_int_data_y_3__7__0_), .A2(
        npu_inst_pe_1_2_7_n50), .B1(npu_inst_pe_1_2_7_n116), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_2_7_n49) );
  INV_X1 npu_inst_pe_1_2_7_U97 ( .A(npu_inst_pe_1_2_7_n49), .ZN(
        npu_inst_pe_1_2_7_n109) );
  AOI22_X1 npu_inst_pe_1_2_7_U96 ( .A1(npu_inst_int_data_y_3__7__0_), .A2(
        npu_inst_pe_1_2_7_n46), .B1(npu_inst_pe_1_2_7_n115), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_2_7_n45) );
  INV_X1 npu_inst_pe_1_2_7_U95 ( .A(npu_inst_pe_1_2_7_n45), .ZN(
        npu_inst_pe_1_2_7_n110) );
  AOI22_X1 npu_inst_pe_1_2_7_U94 ( .A1(npu_inst_int_data_y_3__7__0_), .A2(
        npu_inst_pe_1_2_7_n42), .B1(npu_inst_pe_1_2_7_n114), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_2_7_n41) );
  INV_X1 npu_inst_pe_1_2_7_U93 ( .A(npu_inst_pe_1_2_7_n41), .ZN(
        npu_inst_pe_1_2_7_n111) );
  AOI22_X1 npu_inst_pe_1_2_7_U92 ( .A1(npu_inst_int_data_y_3__7__1_), .A2(
        npu_inst_pe_1_2_7_n58), .B1(npu_inst_pe_1_2_7_n118), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_2_7_n59) );
  INV_X1 npu_inst_pe_1_2_7_U91 ( .A(npu_inst_pe_1_2_7_n59), .ZN(
        npu_inst_pe_1_2_7_n101) );
  AOI22_X1 npu_inst_pe_1_2_7_U90 ( .A1(npu_inst_int_data_y_3__7__1_), .A2(
        npu_inst_pe_1_2_7_n54), .B1(npu_inst_pe_1_2_7_n117), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_2_7_n55) );
  INV_X1 npu_inst_pe_1_2_7_U89 ( .A(npu_inst_pe_1_2_7_n55), .ZN(
        npu_inst_pe_1_2_7_n102) );
  AOI22_X1 npu_inst_pe_1_2_7_U88 ( .A1(npu_inst_int_data_y_3__7__1_), .A2(
        npu_inst_pe_1_2_7_n50), .B1(npu_inst_pe_1_2_7_n116), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_2_7_n51) );
  INV_X1 npu_inst_pe_1_2_7_U87 ( .A(npu_inst_pe_1_2_7_n51), .ZN(
        npu_inst_pe_1_2_7_n103) );
  AOI22_X1 npu_inst_pe_1_2_7_U86 ( .A1(npu_inst_int_data_y_3__7__1_), .A2(
        npu_inst_pe_1_2_7_n46), .B1(npu_inst_pe_1_2_7_n115), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_2_7_n47) );
  INV_X1 npu_inst_pe_1_2_7_U85 ( .A(npu_inst_pe_1_2_7_n47), .ZN(
        npu_inst_pe_1_2_7_n104) );
  AOI22_X1 npu_inst_pe_1_2_7_U84 ( .A1(npu_inst_int_data_y_3__7__1_), .A2(
        npu_inst_pe_1_2_7_n42), .B1(npu_inst_pe_1_2_7_n114), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_2_7_n43) );
  INV_X1 npu_inst_pe_1_2_7_U83 ( .A(npu_inst_pe_1_2_7_n43), .ZN(
        npu_inst_pe_1_2_7_n105) );
  AOI22_X1 npu_inst_pe_1_2_7_U82 ( .A1(npu_inst_pe_1_2_7_n38), .A2(
        npu_inst_int_data_y_3__7__1_), .B1(npu_inst_pe_1_2_7_n113), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_2_7_n39) );
  INV_X1 npu_inst_pe_1_2_7_U81 ( .A(npu_inst_pe_1_2_7_n39), .ZN(
        npu_inst_pe_1_2_7_n106) );
  AND2_X1 npu_inst_pe_1_2_7_U80 ( .A1(npu_inst_pe_1_2_7_N93), .A2(npu_inst_n39), .ZN(npu_inst_int_data_y_2__7__0_) );
  AOI22_X1 npu_inst_pe_1_2_7_U79 ( .A1(npu_inst_pe_1_2_7_n38), .A2(
        npu_inst_int_data_y_3__7__0_), .B1(npu_inst_pe_1_2_7_n113), .B2(
        npu_inst_pe_1_2_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_2_7_n37) );
  INV_X1 npu_inst_pe_1_2_7_U78 ( .A(npu_inst_pe_1_2_7_n37), .ZN(
        npu_inst_pe_1_2_7_n112) );
  AND2_X1 npu_inst_pe_1_2_7_U77 ( .A1(npu_inst_n39), .A2(npu_inst_pe_1_2_7_N94), .ZN(npu_inst_int_data_y_2__7__1_) );
  AOI222_X1 npu_inst_pe_1_2_7_U76 ( .A1(npu_inst_int_data_res_3__7__0_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N73), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N65), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n84) );
  INV_X1 npu_inst_pe_1_2_7_U75 ( .A(npu_inst_pe_1_2_7_n84), .ZN(
        npu_inst_pe_1_2_7_n100) );
  AOI222_X1 npu_inst_pe_1_2_7_U74 ( .A1(npu_inst_pe_1_2_7_n1), .A2(
        npu_inst_int_data_res_3__7__7_), .B1(npu_inst_pe_1_2_7_N80), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N72), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n75) );
  INV_X1 npu_inst_pe_1_2_7_U73 ( .A(npu_inst_pe_1_2_7_n75), .ZN(
        npu_inst_pe_1_2_7_n32) );
  AOI222_X1 npu_inst_pe_1_2_7_U72 ( .A1(npu_inst_int_data_res_3__7__1_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N74), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N66), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n83) );
  INV_X1 npu_inst_pe_1_2_7_U71 ( .A(npu_inst_pe_1_2_7_n83), .ZN(
        npu_inst_pe_1_2_7_n99) );
  AOI222_X1 npu_inst_pe_1_2_7_U70 ( .A1(npu_inst_int_data_res_3__7__3_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N76), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N68), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n81) );
  INV_X1 npu_inst_pe_1_2_7_U69 ( .A(npu_inst_pe_1_2_7_n81), .ZN(
        npu_inst_pe_1_2_7_n36) );
  AOI222_X1 npu_inst_pe_1_2_7_U68 ( .A1(npu_inst_int_data_res_3__7__4_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N77), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N69), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n80) );
  INV_X1 npu_inst_pe_1_2_7_U67 ( .A(npu_inst_pe_1_2_7_n80), .ZN(
        npu_inst_pe_1_2_7_n35) );
  AOI222_X1 npu_inst_pe_1_2_7_U66 ( .A1(npu_inst_int_data_res_3__7__5_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N78), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N70), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n79) );
  INV_X1 npu_inst_pe_1_2_7_U65 ( .A(npu_inst_pe_1_2_7_n79), .ZN(
        npu_inst_pe_1_2_7_n34) );
  AOI222_X1 npu_inst_pe_1_2_7_U64 ( .A1(npu_inst_int_data_res_3__7__6_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N79), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N71), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n78) );
  INV_X1 npu_inst_pe_1_2_7_U63 ( .A(npu_inst_pe_1_2_7_n78), .ZN(
        npu_inst_pe_1_2_7_n33) );
  AND2_X1 npu_inst_pe_1_2_7_U62 ( .A1(npu_inst_int_data_x_2__7__1_), .A2(
        npu_inst_pe_1_2_7_int_q_weight_1_), .ZN(npu_inst_pe_1_2_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_2_7_U61 ( .A1(npu_inst_int_data_x_2__7__0_), .A2(
        npu_inst_pe_1_2_7_int_q_weight_1_), .ZN(npu_inst_pe_1_2_7_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_2_7_U60 ( .A(npu_inst_pe_1_2_7_int_data_1_), .ZN(
        npu_inst_pe_1_2_7_n13) );
  NAND2_X1 npu_inst_pe_1_2_7_U59 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_2_7_n60), .ZN(npu_inst_pe_1_2_7_n74) );
  OAI21_X1 npu_inst_pe_1_2_7_U58 ( .B1(npu_inst_pe_1_2_7_n63), .B2(
        npu_inst_pe_1_2_7_n60), .A(npu_inst_pe_1_2_7_n74), .ZN(
        npu_inst_pe_1_2_7_n97) );
  NAND2_X1 npu_inst_pe_1_2_7_U57 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_2_7_n60), .ZN(npu_inst_pe_1_2_7_n73) );
  OAI21_X1 npu_inst_pe_1_2_7_U56 ( .B1(npu_inst_pe_1_2_7_n61), .B2(
        npu_inst_pe_1_2_7_n60), .A(npu_inst_pe_1_2_7_n73), .ZN(
        npu_inst_pe_1_2_7_n96) );
  NAND2_X1 npu_inst_pe_1_2_7_U55 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_2_7_n56), .ZN(npu_inst_pe_1_2_7_n72) );
  OAI21_X1 npu_inst_pe_1_2_7_U54 ( .B1(npu_inst_pe_1_2_7_n63), .B2(
        npu_inst_pe_1_2_7_n56), .A(npu_inst_pe_1_2_7_n72), .ZN(
        npu_inst_pe_1_2_7_n95) );
  NAND2_X1 npu_inst_pe_1_2_7_U53 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_2_7_n56), .ZN(npu_inst_pe_1_2_7_n71) );
  OAI21_X1 npu_inst_pe_1_2_7_U52 ( .B1(npu_inst_pe_1_2_7_n61), .B2(
        npu_inst_pe_1_2_7_n56), .A(npu_inst_pe_1_2_7_n71), .ZN(
        npu_inst_pe_1_2_7_n94) );
  NAND2_X1 npu_inst_pe_1_2_7_U51 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_2_7_n52), .ZN(npu_inst_pe_1_2_7_n70) );
  OAI21_X1 npu_inst_pe_1_2_7_U50 ( .B1(npu_inst_pe_1_2_7_n63), .B2(
        npu_inst_pe_1_2_7_n52), .A(npu_inst_pe_1_2_7_n70), .ZN(
        npu_inst_pe_1_2_7_n93) );
  NAND2_X1 npu_inst_pe_1_2_7_U49 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_2_7_n52), .ZN(npu_inst_pe_1_2_7_n69) );
  OAI21_X1 npu_inst_pe_1_2_7_U48 ( .B1(npu_inst_pe_1_2_7_n61), .B2(
        npu_inst_pe_1_2_7_n52), .A(npu_inst_pe_1_2_7_n69), .ZN(
        npu_inst_pe_1_2_7_n92) );
  NAND2_X1 npu_inst_pe_1_2_7_U47 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_2_7_n48), .ZN(npu_inst_pe_1_2_7_n68) );
  OAI21_X1 npu_inst_pe_1_2_7_U46 ( .B1(npu_inst_pe_1_2_7_n63), .B2(
        npu_inst_pe_1_2_7_n48), .A(npu_inst_pe_1_2_7_n68), .ZN(
        npu_inst_pe_1_2_7_n91) );
  NAND2_X1 npu_inst_pe_1_2_7_U45 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_2_7_n48), .ZN(npu_inst_pe_1_2_7_n67) );
  OAI21_X1 npu_inst_pe_1_2_7_U44 ( .B1(npu_inst_pe_1_2_7_n61), .B2(
        npu_inst_pe_1_2_7_n48), .A(npu_inst_pe_1_2_7_n67), .ZN(
        npu_inst_pe_1_2_7_n90) );
  NAND2_X1 npu_inst_pe_1_2_7_U43 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_2_7_n44), .ZN(npu_inst_pe_1_2_7_n66) );
  OAI21_X1 npu_inst_pe_1_2_7_U42 ( .B1(npu_inst_pe_1_2_7_n63), .B2(
        npu_inst_pe_1_2_7_n44), .A(npu_inst_pe_1_2_7_n66), .ZN(
        npu_inst_pe_1_2_7_n89) );
  NAND2_X1 npu_inst_pe_1_2_7_U41 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_2_7_n44), .ZN(npu_inst_pe_1_2_7_n65) );
  OAI21_X1 npu_inst_pe_1_2_7_U40 ( .B1(npu_inst_pe_1_2_7_n61), .B2(
        npu_inst_pe_1_2_7_n44), .A(npu_inst_pe_1_2_7_n65), .ZN(
        npu_inst_pe_1_2_7_n88) );
  NAND2_X1 npu_inst_pe_1_2_7_U39 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_2_7_n40), .ZN(npu_inst_pe_1_2_7_n64) );
  OAI21_X1 npu_inst_pe_1_2_7_U38 ( .B1(npu_inst_pe_1_2_7_n63), .B2(
        npu_inst_pe_1_2_7_n40), .A(npu_inst_pe_1_2_7_n64), .ZN(
        npu_inst_pe_1_2_7_n87) );
  NAND2_X1 npu_inst_pe_1_2_7_U37 ( .A1(npu_inst_pe_1_2_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_2_7_n40), .ZN(npu_inst_pe_1_2_7_n62) );
  OAI21_X1 npu_inst_pe_1_2_7_U36 ( .B1(npu_inst_pe_1_2_7_n61), .B2(
        npu_inst_pe_1_2_7_n40), .A(npu_inst_pe_1_2_7_n62), .ZN(
        npu_inst_pe_1_2_7_n86) );
  NOR3_X1 npu_inst_pe_1_2_7_U35 ( .A1(npu_inst_pe_1_2_7_n26), .A2(npu_inst_n39), .A3(npu_inst_int_ckg[40]), .ZN(npu_inst_pe_1_2_7_n85) );
  OR2_X1 npu_inst_pe_1_2_7_U34 ( .A1(npu_inst_pe_1_2_7_n85), .A2(
        npu_inst_pe_1_2_7_n1), .ZN(npu_inst_pe_1_2_7_N84) );
  AOI222_X1 npu_inst_pe_1_2_7_U33 ( .A1(npu_inst_int_data_res_3__7__2_), .A2(
        npu_inst_pe_1_2_7_n1), .B1(npu_inst_pe_1_2_7_N75), .B2(
        npu_inst_pe_1_2_7_n76), .C1(npu_inst_pe_1_2_7_N67), .C2(
        npu_inst_pe_1_2_7_n77), .ZN(npu_inst_pe_1_2_7_n82) );
  INV_X1 npu_inst_pe_1_2_7_U32 ( .A(npu_inst_pe_1_2_7_n82), .ZN(
        npu_inst_pe_1_2_7_n98) );
  INV_X1 npu_inst_pe_1_2_7_U31 ( .A(npu_inst_pe_1_2_7_int_data_0_), .ZN(
        npu_inst_pe_1_2_7_n12) );
  INV_X1 npu_inst_pe_1_2_7_U30 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_2_7_n4)
         );
  AOI22_X1 npu_inst_pe_1_2_7_U29 ( .A1(npu_inst_n39), .A2(
        npu_inst_int_data_y_3__7__1_), .B1(npu_inst_pe_1_2_7_n2), .B2(
        int_i_data_h_npu[11]), .ZN(npu_inst_pe_1_2_7_n63) );
  AOI22_X1 npu_inst_pe_1_2_7_U28 ( .A1(npu_inst_n39), .A2(
        npu_inst_int_data_y_3__7__0_), .B1(npu_inst_pe_1_2_7_n2), .B2(
        int_i_data_h_npu[10]), .ZN(npu_inst_pe_1_2_7_n61) );
  OR3_X1 npu_inst_pe_1_2_7_U27 ( .A1(npu_inst_pe_1_2_7_n5), .A2(
        npu_inst_pe_1_2_7_n7), .A3(npu_inst_pe_1_2_7_n4), .ZN(
        npu_inst_pe_1_2_7_n56) );
  OR3_X1 npu_inst_pe_1_2_7_U26 ( .A1(npu_inst_pe_1_2_7_n4), .A2(
        npu_inst_pe_1_2_7_n7), .A3(npu_inst_pe_1_2_7_n6), .ZN(
        npu_inst_pe_1_2_7_n48) );
  INV_X1 npu_inst_pe_1_2_7_U25 ( .A(npu_inst_pe_1_2_7_n4), .ZN(
        npu_inst_pe_1_2_7_n3) );
  OR3_X1 npu_inst_pe_1_2_7_U24 ( .A1(npu_inst_pe_1_2_7_n3), .A2(
        npu_inst_pe_1_2_7_n7), .A3(npu_inst_pe_1_2_7_n6), .ZN(
        npu_inst_pe_1_2_7_n52) );
  OR3_X1 npu_inst_pe_1_2_7_U23 ( .A1(npu_inst_pe_1_2_7_n5), .A2(
        npu_inst_pe_1_2_7_n7), .A3(npu_inst_pe_1_2_7_n3), .ZN(
        npu_inst_pe_1_2_7_n60) );
  BUF_X1 npu_inst_pe_1_2_7_U22 ( .A(npu_inst_n24), .Z(npu_inst_pe_1_2_7_n1) );
  NOR2_X1 npu_inst_pe_1_2_7_U21 ( .A1(npu_inst_pe_1_2_7_n60), .A2(
        npu_inst_pe_1_2_7_n2), .ZN(npu_inst_pe_1_2_7_n58) );
  NOR2_X1 npu_inst_pe_1_2_7_U20 ( .A1(npu_inst_pe_1_2_7_n56), .A2(
        npu_inst_pe_1_2_7_n2), .ZN(npu_inst_pe_1_2_7_n54) );
  NOR2_X1 npu_inst_pe_1_2_7_U19 ( .A1(npu_inst_pe_1_2_7_n52), .A2(
        npu_inst_pe_1_2_7_n2), .ZN(npu_inst_pe_1_2_7_n50) );
  NOR2_X1 npu_inst_pe_1_2_7_U18 ( .A1(npu_inst_pe_1_2_7_n48), .A2(
        npu_inst_pe_1_2_7_n2), .ZN(npu_inst_pe_1_2_7_n46) );
  NOR2_X1 npu_inst_pe_1_2_7_U17 ( .A1(npu_inst_pe_1_2_7_n40), .A2(
        npu_inst_pe_1_2_7_n2), .ZN(npu_inst_pe_1_2_7_n38) );
  NOR2_X1 npu_inst_pe_1_2_7_U16 ( .A1(npu_inst_pe_1_2_7_n44), .A2(
        npu_inst_pe_1_2_7_n2), .ZN(npu_inst_pe_1_2_7_n42) );
  BUF_X1 npu_inst_pe_1_2_7_U15 ( .A(npu_inst_n84), .Z(npu_inst_pe_1_2_7_n7) );
  INV_X1 npu_inst_pe_1_2_7_U14 ( .A(npu_inst_n107), .ZN(npu_inst_pe_1_2_7_n11)
         );
  INV_X1 npu_inst_pe_1_2_7_U13 ( .A(npu_inst_pe_1_2_7_n38), .ZN(
        npu_inst_pe_1_2_7_n113) );
  INV_X1 npu_inst_pe_1_2_7_U12 ( .A(npu_inst_pe_1_2_7_n58), .ZN(
        npu_inst_pe_1_2_7_n118) );
  INV_X1 npu_inst_pe_1_2_7_U11 ( .A(npu_inst_pe_1_2_7_n54), .ZN(
        npu_inst_pe_1_2_7_n117) );
  INV_X1 npu_inst_pe_1_2_7_U10 ( .A(npu_inst_pe_1_2_7_n50), .ZN(
        npu_inst_pe_1_2_7_n116) );
  INV_X1 npu_inst_pe_1_2_7_U9 ( .A(npu_inst_pe_1_2_7_n46), .ZN(
        npu_inst_pe_1_2_7_n115) );
  INV_X1 npu_inst_pe_1_2_7_U8 ( .A(npu_inst_pe_1_2_7_n42), .ZN(
        npu_inst_pe_1_2_7_n114) );
  BUF_X1 npu_inst_pe_1_2_7_U7 ( .A(npu_inst_pe_1_2_7_n11), .Z(
        npu_inst_pe_1_2_7_n10) );
  BUF_X1 npu_inst_pe_1_2_7_U6 ( .A(npu_inst_pe_1_2_7_n11), .Z(
        npu_inst_pe_1_2_7_n9) );
  BUF_X1 npu_inst_pe_1_2_7_U5 ( .A(npu_inst_pe_1_2_7_n11), .Z(
        npu_inst_pe_1_2_7_n8) );
  NOR2_X1 npu_inst_pe_1_2_7_U4 ( .A1(npu_inst_pe_1_2_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_2_7_n1), .ZN(npu_inst_pe_1_2_7_n76) );
  NOR2_X1 npu_inst_pe_1_2_7_U3 ( .A1(npu_inst_pe_1_2_7_n27), .A2(
        npu_inst_pe_1_2_7_n1), .ZN(npu_inst_pe_1_2_7_n77) );
  FA_X1 npu_inst_pe_1_2_7_sub_77_U2_1 ( .A(npu_inst_int_data_res_2__7__1_), 
        .B(npu_inst_pe_1_2_7_n13), .CI(npu_inst_pe_1_2_7_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_2_7_sub_77_carry_2_), .S(npu_inst_pe_1_2_7_N66) );
  FA_X1 npu_inst_pe_1_2_7_add_79_U1_1 ( .A(npu_inst_int_data_res_2__7__1_), 
        .B(npu_inst_pe_1_2_7_int_data_1_), .CI(
        npu_inst_pe_1_2_7_add_79_carry_1_), .CO(
        npu_inst_pe_1_2_7_add_79_carry_2_), .S(npu_inst_pe_1_2_7_N74) );
  NAND3_X1 npu_inst_pe_1_2_7_U101 ( .A1(npu_inst_pe_1_2_7_n4), .A2(
        npu_inst_pe_1_2_7_n6), .A3(npu_inst_pe_1_2_7_n7), .ZN(
        npu_inst_pe_1_2_7_n44) );
  NAND3_X1 npu_inst_pe_1_2_7_U100 ( .A1(npu_inst_pe_1_2_7_n3), .A2(
        npu_inst_pe_1_2_7_n6), .A3(npu_inst_pe_1_2_7_n7), .ZN(
        npu_inst_pe_1_2_7_n40) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_2_7_n33), .CK(
        npu_inst_pe_1_2_7_net3949), .RN(npu_inst_pe_1_2_7_n8), .Q(
        npu_inst_int_data_res_2__7__6_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_2_7_n34), .CK(
        npu_inst_pe_1_2_7_net3949), .RN(npu_inst_pe_1_2_7_n8), .Q(
        npu_inst_int_data_res_2__7__5_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_2_7_n35), .CK(
        npu_inst_pe_1_2_7_net3949), .RN(npu_inst_pe_1_2_7_n8), .Q(
        npu_inst_int_data_res_2__7__4_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_2_7_n36), .CK(
        npu_inst_pe_1_2_7_net3949), .RN(npu_inst_pe_1_2_7_n8), .Q(
        npu_inst_int_data_res_2__7__3_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_2_7_n98), .CK(
        npu_inst_pe_1_2_7_net3949), .RN(npu_inst_pe_1_2_7_n8), .Q(
        npu_inst_int_data_res_2__7__2_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_2_7_n99), .CK(
        npu_inst_pe_1_2_7_net3949), .RN(npu_inst_pe_1_2_7_n8), .Q(
        npu_inst_int_data_res_2__7__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_2_7_n32), .CK(
        npu_inst_pe_1_2_7_net3949), .RN(npu_inst_pe_1_2_7_n8), .Q(
        npu_inst_int_data_res_2__7__7_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_2_7_n100), 
        .CK(npu_inst_pe_1_2_7_net3949), .RN(npu_inst_pe_1_2_7_n8), .Q(
        npu_inst_int_data_res_2__7__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_weight_reg_0_ ( .D(npu_inst_n93), .CK(
        npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n8), .Q(
        npu_inst_pe_1_2_7_int_q_weight_0_), .QN(npu_inst_pe_1_2_7_n27) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_weight_reg_1_ ( .D(npu_inst_n99), .CK(
        npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n8), .Q(
        npu_inst_pe_1_2_7_int_q_weight_1_), .QN(npu_inst_pe_1_2_7_n26) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_2_7_n112), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n8), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_2_7_n106), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n8), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_2_7_n111), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_2_7_n105), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_2_7_n110), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_2_7_n104), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_2_7_n109), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_2_7_n103), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_2_7_n108), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_2_7_n102), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_2_7_n107), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_2_7_n101), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_2_7_n86), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_2_7_n87), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n9), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_2_7_n88), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_2_7_n89), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_2_7_n90), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_2_7_n91), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_2_7_n92), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_2_7_n93), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_2_7_n94), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_2_7_n95), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_2_7_n96), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_2_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_2_7_n97), 
        .CK(npu_inst_pe_1_2_7_net3955), .RN(npu_inst_pe_1_2_7_n10), .Q(
        npu_inst_pe_1_2_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_2_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_2_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_2_7_net3949) );
  CLKGATETST_X1 npu_inst_pe_1_2_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n46), .SE(1'b0), .GCK(npu_inst_pe_1_2_7_net3955) );
  MUX2_X1 npu_inst_pe_1_3_0_U153 ( .A(npu_inst_pe_1_3_0_n31), .B(
        npu_inst_pe_1_3_0_n28), .S(npu_inst_pe_1_3_0_n7), .Z(
        npu_inst_pe_1_3_0_N93) );
  MUX2_X1 npu_inst_pe_1_3_0_U152 ( .A(npu_inst_pe_1_3_0_n30), .B(
        npu_inst_pe_1_3_0_n29), .S(npu_inst_pe_1_3_0_n5), .Z(
        npu_inst_pe_1_3_0_n31) );
  MUX2_X1 npu_inst_pe_1_3_0_U151 ( .A(npu_inst_pe_1_3_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_0_n3), .Z(
        npu_inst_pe_1_3_0_n30) );
  MUX2_X1 npu_inst_pe_1_3_0_U150 ( .A(npu_inst_pe_1_3_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_0_n3), .Z(
        npu_inst_pe_1_3_0_n29) );
  MUX2_X1 npu_inst_pe_1_3_0_U149 ( .A(npu_inst_pe_1_3_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_0_n3), .Z(
        npu_inst_pe_1_3_0_n28) );
  MUX2_X1 npu_inst_pe_1_3_0_U148 ( .A(npu_inst_pe_1_3_0_n25), .B(
        npu_inst_pe_1_3_0_n22), .S(npu_inst_pe_1_3_0_n7), .Z(
        npu_inst_pe_1_3_0_N94) );
  MUX2_X1 npu_inst_pe_1_3_0_U147 ( .A(npu_inst_pe_1_3_0_n24), .B(
        npu_inst_pe_1_3_0_n23), .S(npu_inst_pe_1_3_0_n5), .Z(
        npu_inst_pe_1_3_0_n25) );
  MUX2_X1 npu_inst_pe_1_3_0_U146 ( .A(npu_inst_pe_1_3_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_0_n3), .Z(
        npu_inst_pe_1_3_0_n24) );
  MUX2_X1 npu_inst_pe_1_3_0_U145 ( .A(npu_inst_pe_1_3_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_0_n3), .Z(
        npu_inst_pe_1_3_0_n23) );
  MUX2_X1 npu_inst_pe_1_3_0_U144 ( .A(npu_inst_pe_1_3_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_0_n3), .Z(
        npu_inst_pe_1_3_0_n22) );
  MUX2_X1 npu_inst_pe_1_3_0_U143 ( .A(npu_inst_pe_1_3_0_n21), .B(
        npu_inst_pe_1_3_0_n18), .S(npu_inst_pe_1_3_0_n7), .Z(
        npu_inst_pe_1_3_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_3_0_U142 ( .A(npu_inst_pe_1_3_0_n20), .B(
        npu_inst_pe_1_3_0_n19), .S(npu_inst_pe_1_3_0_n5), .Z(
        npu_inst_pe_1_3_0_n21) );
  MUX2_X1 npu_inst_pe_1_3_0_U141 ( .A(npu_inst_pe_1_3_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_0_n3), .Z(
        npu_inst_pe_1_3_0_n20) );
  MUX2_X1 npu_inst_pe_1_3_0_U140 ( .A(npu_inst_pe_1_3_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_0_n3), .Z(
        npu_inst_pe_1_3_0_n19) );
  MUX2_X1 npu_inst_pe_1_3_0_U139 ( .A(npu_inst_pe_1_3_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_0_n3), .Z(
        npu_inst_pe_1_3_0_n18) );
  MUX2_X1 npu_inst_pe_1_3_0_U138 ( .A(npu_inst_pe_1_3_0_n17), .B(
        npu_inst_pe_1_3_0_n14), .S(npu_inst_pe_1_3_0_n7), .Z(
        npu_inst_pe_1_3_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_3_0_U137 ( .A(npu_inst_pe_1_3_0_n16), .B(
        npu_inst_pe_1_3_0_n15), .S(npu_inst_pe_1_3_0_n5), .Z(
        npu_inst_pe_1_3_0_n17) );
  MUX2_X1 npu_inst_pe_1_3_0_U136 ( .A(npu_inst_pe_1_3_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_0_n3), .Z(
        npu_inst_pe_1_3_0_n16) );
  MUX2_X1 npu_inst_pe_1_3_0_U135 ( .A(npu_inst_pe_1_3_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_0_n3), .Z(
        npu_inst_pe_1_3_0_n15) );
  MUX2_X1 npu_inst_pe_1_3_0_U134 ( .A(npu_inst_pe_1_3_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_0_n3), .Z(
        npu_inst_pe_1_3_0_n14) );
  XOR2_X1 npu_inst_pe_1_3_0_U133 ( .A(npu_inst_pe_1_3_0_int_data_0_), .B(
        npu_inst_int_data_res_3__0__0_), .Z(npu_inst_pe_1_3_0_N73) );
  AND2_X1 npu_inst_pe_1_3_0_U132 ( .A1(npu_inst_int_data_res_3__0__0_), .A2(
        npu_inst_pe_1_3_0_int_data_0_), .ZN(npu_inst_pe_1_3_0_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_0_U131 ( .A(npu_inst_int_data_res_3__0__0_), .B(
        npu_inst_pe_1_3_0_n12), .ZN(npu_inst_pe_1_3_0_N65) );
  OR2_X1 npu_inst_pe_1_3_0_U130 ( .A1(npu_inst_pe_1_3_0_n12), .A2(
        npu_inst_int_data_res_3__0__0_), .ZN(npu_inst_pe_1_3_0_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_0_U129 ( .A(npu_inst_int_data_res_3__0__2_), .B(
        npu_inst_pe_1_3_0_add_79_carry_2_), .Z(npu_inst_pe_1_3_0_N75) );
  AND2_X1 npu_inst_pe_1_3_0_U128 ( .A1(npu_inst_pe_1_3_0_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_3__0__2_), .ZN(
        npu_inst_pe_1_3_0_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_0_U127 ( .A(npu_inst_int_data_res_3__0__3_), .B(
        npu_inst_pe_1_3_0_add_79_carry_3_), .Z(npu_inst_pe_1_3_0_N76) );
  AND2_X1 npu_inst_pe_1_3_0_U126 ( .A1(npu_inst_pe_1_3_0_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_3__0__3_), .ZN(
        npu_inst_pe_1_3_0_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_0_U125 ( .A(npu_inst_int_data_res_3__0__4_), .B(
        npu_inst_pe_1_3_0_add_79_carry_4_), .Z(npu_inst_pe_1_3_0_N77) );
  AND2_X1 npu_inst_pe_1_3_0_U124 ( .A1(npu_inst_pe_1_3_0_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_3__0__4_), .ZN(
        npu_inst_pe_1_3_0_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_0_U123 ( .A(npu_inst_int_data_res_3__0__5_), .B(
        npu_inst_pe_1_3_0_add_79_carry_5_), .Z(npu_inst_pe_1_3_0_N78) );
  AND2_X1 npu_inst_pe_1_3_0_U122 ( .A1(npu_inst_pe_1_3_0_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_3__0__5_), .ZN(
        npu_inst_pe_1_3_0_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_0_U121 ( .A(npu_inst_int_data_res_3__0__6_), .B(
        npu_inst_pe_1_3_0_add_79_carry_6_), .Z(npu_inst_pe_1_3_0_N79) );
  AND2_X1 npu_inst_pe_1_3_0_U120 ( .A1(npu_inst_pe_1_3_0_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_3__0__6_), .ZN(
        npu_inst_pe_1_3_0_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_0_U119 ( .A(npu_inst_int_data_res_3__0__7_), .B(
        npu_inst_pe_1_3_0_add_79_carry_7_), .Z(npu_inst_pe_1_3_0_N80) );
  XNOR2_X1 npu_inst_pe_1_3_0_U118 ( .A(npu_inst_pe_1_3_0_sub_77_carry_2_), .B(
        npu_inst_int_data_res_3__0__2_), .ZN(npu_inst_pe_1_3_0_N67) );
  OR2_X1 npu_inst_pe_1_3_0_U117 ( .A1(npu_inst_int_data_res_3__0__2_), .A2(
        npu_inst_pe_1_3_0_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_3_0_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_0_U116 ( .A(npu_inst_pe_1_3_0_sub_77_carry_3_), .B(
        npu_inst_int_data_res_3__0__3_), .ZN(npu_inst_pe_1_3_0_N68) );
  OR2_X1 npu_inst_pe_1_3_0_U115 ( .A1(npu_inst_int_data_res_3__0__3_), .A2(
        npu_inst_pe_1_3_0_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_3_0_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_0_U114 ( .A(npu_inst_pe_1_3_0_sub_77_carry_4_), .B(
        npu_inst_int_data_res_3__0__4_), .ZN(npu_inst_pe_1_3_0_N69) );
  OR2_X1 npu_inst_pe_1_3_0_U113 ( .A1(npu_inst_int_data_res_3__0__4_), .A2(
        npu_inst_pe_1_3_0_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_3_0_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_0_U112 ( .A(npu_inst_pe_1_3_0_sub_77_carry_5_), .B(
        npu_inst_int_data_res_3__0__5_), .ZN(npu_inst_pe_1_3_0_N70) );
  OR2_X1 npu_inst_pe_1_3_0_U111 ( .A1(npu_inst_int_data_res_3__0__5_), .A2(
        npu_inst_pe_1_3_0_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_3_0_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_0_U110 ( .A(npu_inst_pe_1_3_0_sub_77_carry_6_), .B(
        npu_inst_int_data_res_3__0__6_), .ZN(npu_inst_pe_1_3_0_N71) );
  OR2_X1 npu_inst_pe_1_3_0_U109 ( .A1(npu_inst_int_data_res_3__0__6_), .A2(
        npu_inst_pe_1_3_0_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_3_0_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_0_U108 ( .A(npu_inst_int_data_res_3__0__7_), .B(
        npu_inst_pe_1_3_0_sub_77_carry_7_), .ZN(npu_inst_pe_1_3_0_N72) );
  INV_X1 npu_inst_pe_1_3_0_U107 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_3_0_n6)
         );
  INV_X1 npu_inst_pe_1_3_0_U106 ( .A(npu_inst_pe_1_3_0_n6), .ZN(
        npu_inst_pe_1_3_0_n5) );
  INV_X1 npu_inst_pe_1_3_0_U105 ( .A(npu_inst_n39), .ZN(npu_inst_pe_1_3_0_n2)
         );
  AOI22_X1 npu_inst_pe_1_3_0_U104 ( .A1(npu_inst_int_data_y_4__0__0_), .A2(
        npu_inst_pe_1_3_0_n58), .B1(npu_inst_pe_1_3_0_n118), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_0_n57) );
  INV_X1 npu_inst_pe_1_3_0_U103 ( .A(npu_inst_pe_1_3_0_n57), .ZN(
        npu_inst_pe_1_3_0_n107) );
  AOI22_X1 npu_inst_pe_1_3_0_U102 ( .A1(npu_inst_int_data_y_4__0__0_), .A2(
        npu_inst_pe_1_3_0_n54), .B1(npu_inst_pe_1_3_0_n117), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_0_n53) );
  INV_X1 npu_inst_pe_1_3_0_U99 ( .A(npu_inst_pe_1_3_0_n53), .ZN(
        npu_inst_pe_1_3_0_n108) );
  AOI22_X1 npu_inst_pe_1_3_0_U98 ( .A1(npu_inst_int_data_y_4__0__0_), .A2(
        npu_inst_pe_1_3_0_n50), .B1(npu_inst_pe_1_3_0_n116), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_0_n49) );
  INV_X1 npu_inst_pe_1_3_0_U97 ( .A(npu_inst_pe_1_3_0_n49), .ZN(
        npu_inst_pe_1_3_0_n109) );
  AOI22_X1 npu_inst_pe_1_3_0_U96 ( .A1(npu_inst_int_data_y_4__0__0_), .A2(
        npu_inst_pe_1_3_0_n46), .B1(npu_inst_pe_1_3_0_n115), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_0_n45) );
  INV_X1 npu_inst_pe_1_3_0_U95 ( .A(npu_inst_pe_1_3_0_n45), .ZN(
        npu_inst_pe_1_3_0_n110) );
  AOI22_X1 npu_inst_pe_1_3_0_U94 ( .A1(npu_inst_int_data_y_4__0__0_), .A2(
        npu_inst_pe_1_3_0_n42), .B1(npu_inst_pe_1_3_0_n114), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_0_n41) );
  INV_X1 npu_inst_pe_1_3_0_U93 ( .A(npu_inst_pe_1_3_0_n41), .ZN(
        npu_inst_pe_1_3_0_n111) );
  AOI22_X1 npu_inst_pe_1_3_0_U92 ( .A1(npu_inst_int_data_y_4__0__1_), .A2(
        npu_inst_pe_1_3_0_n58), .B1(npu_inst_pe_1_3_0_n118), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_0_n59) );
  INV_X1 npu_inst_pe_1_3_0_U91 ( .A(npu_inst_pe_1_3_0_n59), .ZN(
        npu_inst_pe_1_3_0_n101) );
  AOI22_X1 npu_inst_pe_1_3_0_U90 ( .A1(npu_inst_int_data_y_4__0__1_), .A2(
        npu_inst_pe_1_3_0_n54), .B1(npu_inst_pe_1_3_0_n117), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_0_n55) );
  INV_X1 npu_inst_pe_1_3_0_U89 ( .A(npu_inst_pe_1_3_0_n55), .ZN(
        npu_inst_pe_1_3_0_n102) );
  AOI22_X1 npu_inst_pe_1_3_0_U88 ( .A1(npu_inst_int_data_y_4__0__1_), .A2(
        npu_inst_pe_1_3_0_n50), .B1(npu_inst_pe_1_3_0_n116), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_0_n51) );
  INV_X1 npu_inst_pe_1_3_0_U87 ( .A(npu_inst_pe_1_3_0_n51), .ZN(
        npu_inst_pe_1_3_0_n103) );
  AOI22_X1 npu_inst_pe_1_3_0_U86 ( .A1(npu_inst_int_data_y_4__0__1_), .A2(
        npu_inst_pe_1_3_0_n46), .B1(npu_inst_pe_1_3_0_n115), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_0_n47) );
  INV_X1 npu_inst_pe_1_3_0_U85 ( .A(npu_inst_pe_1_3_0_n47), .ZN(
        npu_inst_pe_1_3_0_n104) );
  AOI22_X1 npu_inst_pe_1_3_0_U84 ( .A1(npu_inst_int_data_y_4__0__1_), .A2(
        npu_inst_pe_1_3_0_n42), .B1(npu_inst_pe_1_3_0_n114), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_0_n43) );
  INV_X1 npu_inst_pe_1_3_0_U83 ( .A(npu_inst_pe_1_3_0_n43), .ZN(
        npu_inst_pe_1_3_0_n105) );
  AOI22_X1 npu_inst_pe_1_3_0_U82 ( .A1(npu_inst_pe_1_3_0_n38), .A2(
        npu_inst_int_data_y_4__0__1_), .B1(npu_inst_pe_1_3_0_n113), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_0_n39) );
  INV_X1 npu_inst_pe_1_3_0_U81 ( .A(npu_inst_pe_1_3_0_n39), .ZN(
        npu_inst_pe_1_3_0_n106) );
  AND2_X1 npu_inst_pe_1_3_0_U80 ( .A1(npu_inst_pe_1_3_0_N93), .A2(npu_inst_n39), .ZN(npu_inst_int_data_y_3__0__0_) );
  NAND2_X1 npu_inst_pe_1_3_0_U79 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_0_n60), .ZN(npu_inst_pe_1_3_0_n74) );
  OAI21_X1 npu_inst_pe_1_3_0_U78 ( .B1(npu_inst_pe_1_3_0_n63), .B2(
        npu_inst_pe_1_3_0_n60), .A(npu_inst_pe_1_3_0_n74), .ZN(
        npu_inst_pe_1_3_0_n97) );
  NAND2_X1 npu_inst_pe_1_3_0_U77 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_0_n60), .ZN(npu_inst_pe_1_3_0_n73) );
  OAI21_X1 npu_inst_pe_1_3_0_U76 ( .B1(npu_inst_pe_1_3_0_n61), .B2(
        npu_inst_pe_1_3_0_n60), .A(npu_inst_pe_1_3_0_n73), .ZN(
        npu_inst_pe_1_3_0_n96) );
  NAND2_X1 npu_inst_pe_1_3_0_U75 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_0_n56), .ZN(npu_inst_pe_1_3_0_n72) );
  OAI21_X1 npu_inst_pe_1_3_0_U74 ( .B1(npu_inst_pe_1_3_0_n63), .B2(
        npu_inst_pe_1_3_0_n56), .A(npu_inst_pe_1_3_0_n72), .ZN(
        npu_inst_pe_1_3_0_n95) );
  NAND2_X1 npu_inst_pe_1_3_0_U73 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_0_n56), .ZN(npu_inst_pe_1_3_0_n71) );
  OAI21_X1 npu_inst_pe_1_3_0_U72 ( .B1(npu_inst_pe_1_3_0_n61), .B2(
        npu_inst_pe_1_3_0_n56), .A(npu_inst_pe_1_3_0_n71), .ZN(
        npu_inst_pe_1_3_0_n94) );
  NAND2_X1 npu_inst_pe_1_3_0_U71 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_0_n52), .ZN(npu_inst_pe_1_3_0_n70) );
  OAI21_X1 npu_inst_pe_1_3_0_U70 ( .B1(npu_inst_pe_1_3_0_n63), .B2(
        npu_inst_pe_1_3_0_n52), .A(npu_inst_pe_1_3_0_n70), .ZN(
        npu_inst_pe_1_3_0_n93) );
  NAND2_X1 npu_inst_pe_1_3_0_U69 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_0_n52), .ZN(npu_inst_pe_1_3_0_n69) );
  OAI21_X1 npu_inst_pe_1_3_0_U68 ( .B1(npu_inst_pe_1_3_0_n61), .B2(
        npu_inst_pe_1_3_0_n52), .A(npu_inst_pe_1_3_0_n69), .ZN(
        npu_inst_pe_1_3_0_n92) );
  NAND2_X1 npu_inst_pe_1_3_0_U67 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_0_n48), .ZN(npu_inst_pe_1_3_0_n68) );
  OAI21_X1 npu_inst_pe_1_3_0_U66 ( .B1(npu_inst_pe_1_3_0_n63), .B2(
        npu_inst_pe_1_3_0_n48), .A(npu_inst_pe_1_3_0_n68), .ZN(
        npu_inst_pe_1_3_0_n91) );
  NAND2_X1 npu_inst_pe_1_3_0_U65 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_0_n48), .ZN(npu_inst_pe_1_3_0_n67) );
  OAI21_X1 npu_inst_pe_1_3_0_U64 ( .B1(npu_inst_pe_1_3_0_n61), .B2(
        npu_inst_pe_1_3_0_n48), .A(npu_inst_pe_1_3_0_n67), .ZN(
        npu_inst_pe_1_3_0_n90) );
  NAND2_X1 npu_inst_pe_1_3_0_U63 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_0_n44), .ZN(npu_inst_pe_1_3_0_n66) );
  OAI21_X1 npu_inst_pe_1_3_0_U62 ( .B1(npu_inst_pe_1_3_0_n63), .B2(
        npu_inst_pe_1_3_0_n44), .A(npu_inst_pe_1_3_0_n66), .ZN(
        npu_inst_pe_1_3_0_n89) );
  NAND2_X1 npu_inst_pe_1_3_0_U61 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_0_n44), .ZN(npu_inst_pe_1_3_0_n65) );
  OAI21_X1 npu_inst_pe_1_3_0_U60 ( .B1(npu_inst_pe_1_3_0_n61), .B2(
        npu_inst_pe_1_3_0_n44), .A(npu_inst_pe_1_3_0_n65), .ZN(
        npu_inst_pe_1_3_0_n88) );
  NAND2_X1 npu_inst_pe_1_3_0_U59 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_0_n40), .ZN(npu_inst_pe_1_3_0_n64) );
  OAI21_X1 npu_inst_pe_1_3_0_U58 ( .B1(npu_inst_pe_1_3_0_n63), .B2(
        npu_inst_pe_1_3_0_n40), .A(npu_inst_pe_1_3_0_n64), .ZN(
        npu_inst_pe_1_3_0_n87) );
  NAND2_X1 npu_inst_pe_1_3_0_U57 ( .A1(npu_inst_pe_1_3_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_0_n40), .ZN(npu_inst_pe_1_3_0_n62) );
  OAI21_X1 npu_inst_pe_1_3_0_U56 ( .B1(npu_inst_pe_1_3_0_n61), .B2(
        npu_inst_pe_1_3_0_n40), .A(npu_inst_pe_1_3_0_n62), .ZN(
        npu_inst_pe_1_3_0_n86) );
  AOI22_X1 npu_inst_pe_1_3_0_U55 ( .A1(npu_inst_pe_1_3_0_n38), .A2(
        npu_inst_int_data_y_4__0__0_), .B1(npu_inst_pe_1_3_0_n113), .B2(
        npu_inst_pe_1_3_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_0_n37) );
  INV_X1 npu_inst_pe_1_3_0_U54 ( .A(npu_inst_pe_1_3_0_n37), .ZN(
        npu_inst_pe_1_3_0_n112) );
  AND2_X1 npu_inst_pe_1_3_0_U53 ( .A1(npu_inst_n39), .A2(npu_inst_pe_1_3_0_N94), .ZN(npu_inst_int_data_y_3__0__1_) );
  AOI222_X1 npu_inst_pe_1_3_0_U52 ( .A1(npu_inst_int_data_res_4__0__0_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N73), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N65), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n84) );
  INV_X1 npu_inst_pe_1_3_0_U51 ( .A(npu_inst_pe_1_3_0_n84), .ZN(
        npu_inst_pe_1_3_0_n100) );
  AOI222_X1 npu_inst_pe_1_3_0_U50 ( .A1(npu_inst_pe_1_3_0_n1), .A2(
        npu_inst_int_data_res_4__0__7_), .B1(npu_inst_pe_1_3_0_N80), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N72), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n75) );
  INV_X1 npu_inst_pe_1_3_0_U49 ( .A(npu_inst_pe_1_3_0_n75), .ZN(
        npu_inst_pe_1_3_0_n32) );
  AOI222_X1 npu_inst_pe_1_3_0_U48 ( .A1(npu_inst_int_data_res_4__0__1_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N74), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N66), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n83) );
  INV_X1 npu_inst_pe_1_3_0_U47 ( .A(npu_inst_pe_1_3_0_n83), .ZN(
        npu_inst_pe_1_3_0_n99) );
  AOI222_X1 npu_inst_pe_1_3_0_U46 ( .A1(npu_inst_int_data_res_4__0__3_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N76), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N68), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n81) );
  INV_X1 npu_inst_pe_1_3_0_U45 ( .A(npu_inst_pe_1_3_0_n81), .ZN(
        npu_inst_pe_1_3_0_n36) );
  AOI222_X1 npu_inst_pe_1_3_0_U44 ( .A1(npu_inst_int_data_res_4__0__4_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N77), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N69), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n80) );
  INV_X1 npu_inst_pe_1_3_0_U43 ( .A(npu_inst_pe_1_3_0_n80), .ZN(
        npu_inst_pe_1_3_0_n35) );
  AOI222_X1 npu_inst_pe_1_3_0_U42 ( .A1(npu_inst_int_data_res_4__0__5_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N78), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N70), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n79) );
  INV_X1 npu_inst_pe_1_3_0_U41 ( .A(npu_inst_pe_1_3_0_n79), .ZN(
        npu_inst_pe_1_3_0_n34) );
  AOI222_X1 npu_inst_pe_1_3_0_U40 ( .A1(npu_inst_int_data_res_4__0__6_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N79), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N71), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n78) );
  INV_X1 npu_inst_pe_1_3_0_U39 ( .A(npu_inst_pe_1_3_0_n78), .ZN(
        npu_inst_pe_1_3_0_n33) );
  AND2_X1 npu_inst_pe_1_3_0_U38 ( .A1(npu_inst_pe_1_3_0_o_data_h_1_), .A2(
        npu_inst_pe_1_3_0_int_q_weight_1_), .ZN(npu_inst_pe_1_3_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_0_U37 ( .A1(npu_inst_pe_1_3_0_o_data_h_0_), .A2(
        npu_inst_pe_1_3_0_int_q_weight_1_), .ZN(npu_inst_pe_1_3_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_3_0_U36 ( .A(npu_inst_pe_1_3_0_int_data_1_), .ZN(
        npu_inst_pe_1_3_0_n13) );
  NOR3_X1 npu_inst_pe_1_3_0_U35 ( .A1(npu_inst_pe_1_3_0_n26), .A2(npu_inst_n39), .A3(npu_inst_int_ckg[39]), .ZN(npu_inst_pe_1_3_0_n85) );
  OR2_X1 npu_inst_pe_1_3_0_U34 ( .A1(npu_inst_pe_1_3_0_n85), .A2(
        npu_inst_pe_1_3_0_n1), .ZN(npu_inst_pe_1_3_0_N84) );
  AOI222_X1 npu_inst_pe_1_3_0_U33 ( .A1(npu_inst_int_data_res_4__0__2_), .A2(
        npu_inst_pe_1_3_0_n1), .B1(npu_inst_pe_1_3_0_N75), .B2(
        npu_inst_pe_1_3_0_n76), .C1(npu_inst_pe_1_3_0_N67), .C2(
        npu_inst_pe_1_3_0_n77), .ZN(npu_inst_pe_1_3_0_n82) );
  INV_X1 npu_inst_pe_1_3_0_U32 ( .A(npu_inst_pe_1_3_0_n82), .ZN(
        npu_inst_pe_1_3_0_n98) );
  AOI22_X1 npu_inst_pe_1_3_0_U31 ( .A1(npu_inst_n39), .A2(
        npu_inst_int_data_y_4__0__1_), .B1(npu_inst_pe_1_3_0_n2), .B2(
        npu_inst_int_data_x_3__1__1_), .ZN(npu_inst_pe_1_3_0_n63) );
  AOI22_X1 npu_inst_pe_1_3_0_U30 ( .A1(npu_inst_n39), .A2(
        npu_inst_int_data_y_4__0__0_), .B1(npu_inst_pe_1_3_0_n2), .B2(
        npu_inst_int_data_x_3__1__0_), .ZN(npu_inst_pe_1_3_0_n61) );
  INV_X1 npu_inst_pe_1_3_0_U29 ( .A(npu_inst_pe_1_3_0_int_data_0_), .ZN(
        npu_inst_pe_1_3_0_n12) );
  INV_X1 npu_inst_pe_1_3_0_U28 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_3_0_n4)
         );
  OR3_X1 npu_inst_pe_1_3_0_U27 ( .A1(npu_inst_pe_1_3_0_n5), .A2(
        npu_inst_pe_1_3_0_n7), .A3(npu_inst_pe_1_3_0_n4), .ZN(
        npu_inst_pe_1_3_0_n56) );
  OR3_X1 npu_inst_pe_1_3_0_U26 ( .A1(npu_inst_pe_1_3_0_n4), .A2(
        npu_inst_pe_1_3_0_n7), .A3(npu_inst_pe_1_3_0_n6), .ZN(
        npu_inst_pe_1_3_0_n48) );
  INV_X1 npu_inst_pe_1_3_0_U25 ( .A(npu_inst_pe_1_3_0_n4), .ZN(
        npu_inst_pe_1_3_0_n3) );
  OR3_X1 npu_inst_pe_1_3_0_U24 ( .A1(npu_inst_pe_1_3_0_n3), .A2(
        npu_inst_pe_1_3_0_n7), .A3(npu_inst_pe_1_3_0_n6), .ZN(
        npu_inst_pe_1_3_0_n52) );
  OR3_X1 npu_inst_pe_1_3_0_U23 ( .A1(npu_inst_pe_1_3_0_n5), .A2(
        npu_inst_pe_1_3_0_n7), .A3(npu_inst_pe_1_3_0_n3), .ZN(
        npu_inst_pe_1_3_0_n60) );
  BUF_X1 npu_inst_pe_1_3_0_U22 ( .A(npu_inst_n24), .Z(npu_inst_pe_1_3_0_n1) );
  NOR2_X1 npu_inst_pe_1_3_0_U21 ( .A1(npu_inst_pe_1_3_0_n60), .A2(
        npu_inst_pe_1_3_0_n2), .ZN(npu_inst_pe_1_3_0_n58) );
  NOR2_X1 npu_inst_pe_1_3_0_U20 ( .A1(npu_inst_pe_1_3_0_n56), .A2(
        npu_inst_pe_1_3_0_n2), .ZN(npu_inst_pe_1_3_0_n54) );
  NOR2_X1 npu_inst_pe_1_3_0_U19 ( .A1(npu_inst_pe_1_3_0_n52), .A2(
        npu_inst_pe_1_3_0_n2), .ZN(npu_inst_pe_1_3_0_n50) );
  NOR2_X1 npu_inst_pe_1_3_0_U18 ( .A1(npu_inst_pe_1_3_0_n48), .A2(
        npu_inst_pe_1_3_0_n2), .ZN(npu_inst_pe_1_3_0_n46) );
  NOR2_X1 npu_inst_pe_1_3_0_U17 ( .A1(npu_inst_pe_1_3_0_n40), .A2(
        npu_inst_pe_1_3_0_n2), .ZN(npu_inst_pe_1_3_0_n38) );
  NOR2_X1 npu_inst_pe_1_3_0_U16 ( .A1(npu_inst_pe_1_3_0_n44), .A2(
        npu_inst_pe_1_3_0_n2), .ZN(npu_inst_pe_1_3_0_n42) );
  BUF_X1 npu_inst_pe_1_3_0_U15 ( .A(npu_inst_n83), .Z(npu_inst_pe_1_3_0_n7) );
  INV_X1 npu_inst_pe_1_3_0_U14 ( .A(npu_inst_n107), .ZN(npu_inst_pe_1_3_0_n11)
         );
  INV_X1 npu_inst_pe_1_3_0_U13 ( .A(npu_inst_pe_1_3_0_n38), .ZN(
        npu_inst_pe_1_3_0_n113) );
  INV_X1 npu_inst_pe_1_3_0_U12 ( .A(npu_inst_pe_1_3_0_n58), .ZN(
        npu_inst_pe_1_3_0_n118) );
  INV_X1 npu_inst_pe_1_3_0_U11 ( .A(npu_inst_pe_1_3_0_n54), .ZN(
        npu_inst_pe_1_3_0_n117) );
  INV_X1 npu_inst_pe_1_3_0_U10 ( .A(npu_inst_pe_1_3_0_n50), .ZN(
        npu_inst_pe_1_3_0_n116) );
  INV_X1 npu_inst_pe_1_3_0_U9 ( .A(npu_inst_pe_1_3_0_n46), .ZN(
        npu_inst_pe_1_3_0_n115) );
  INV_X1 npu_inst_pe_1_3_0_U8 ( .A(npu_inst_pe_1_3_0_n42), .ZN(
        npu_inst_pe_1_3_0_n114) );
  BUF_X1 npu_inst_pe_1_3_0_U7 ( .A(npu_inst_pe_1_3_0_n11), .Z(
        npu_inst_pe_1_3_0_n10) );
  BUF_X1 npu_inst_pe_1_3_0_U6 ( .A(npu_inst_pe_1_3_0_n11), .Z(
        npu_inst_pe_1_3_0_n9) );
  BUF_X1 npu_inst_pe_1_3_0_U5 ( .A(npu_inst_pe_1_3_0_n11), .Z(
        npu_inst_pe_1_3_0_n8) );
  NOR2_X1 npu_inst_pe_1_3_0_U4 ( .A1(npu_inst_pe_1_3_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_0_n1), .ZN(npu_inst_pe_1_3_0_n76) );
  NOR2_X1 npu_inst_pe_1_3_0_U3 ( .A1(npu_inst_pe_1_3_0_n27), .A2(
        npu_inst_pe_1_3_0_n1), .ZN(npu_inst_pe_1_3_0_n77) );
  FA_X1 npu_inst_pe_1_3_0_sub_77_U2_1 ( .A(npu_inst_int_data_res_3__0__1_), 
        .B(npu_inst_pe_1_3_0_n13), .CI(npu_inst_pe_1_3_0_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_3_0_sub_77_carry_2_), .S(npu_inst_pe_1_3_0_N66) );
  FA_X1 npu_inst_pe_1_3_0_add_79_U1_1 ( .A(npu_inst_int_data_res_3__0__1_), 
        .B(npu_inst_pe_1_3_0_int_data_1_), .CI(
        npu_inst_pe_1_3_0_add_79_carry_1_), .CO(
        npu_inst_pe_1_3_0_add_79_carry_2_), .S(npu_inst_pe_1_3_0_N74) );
  NAND3_X1 npu_inst_pe_1_3_0_U101 ( .A1(npu_inst_pe_1_3_0_n4), .A2(
        npu_inst_pe_1_3_0_n6), .A3(npu_inst_pe_1_3_0_n7), .ZN(
        npu_inst_pe_1_3_0_n44) );
  NAND3_X1 npu_inst_pe_1_3_0_U100 ( .A1(npu_inst_pe_1_3_0_n3), .A2(
        npu_inst_pe_1_3_0_n6), .A3(npu_inst_pe_1_3_0_n7), .ZN(
        npu_inst_pe_1_3_0_n40) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_0_n33), .CK(
        npu_inst_pe_1_3_0_net3926), .RN(npu_inst_pe_1_3_0_n8), .Q(
        npu_inst_int_data_res_3__0__6_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_0_n34), .CK(
        npu_inst_pe_1_3_0_net3926), .RN(npu_inst_pe_1_3_0_n8), .Q(
        npu_inst_int_data_res_3__0__5_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_0_n35), .CK(
        npu_inst_pe_1_3_0_net3926), .RN(npu_inst_pe_1_3_0_n8), .Q(
        npu_inst_int_data_res_3__0__4_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_0_n36), .CK(
        npu_inst_pe_1_3_0_net3926), .RN(npu_inst_pe_1_3_0_n8), .Q(
        npu_inst_int_data_res_3__0__3_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_0_n98), .CK(
        npu_inst_pe_1_3_0_net3926), .RN(npu_inst_pe_1_3_0_n8), .Q(
        npu_inst_int_data_res_3__0__2_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_0_n99), .CK(
        npu_inst_pe_1_3_0_net3926), .RN(npu_inst_pe_1_3_0_n8), .Q(
        npu_inst_int_data_res_3__0__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_0_n32), .CK(
        npu_inst_pe_1_3_0_net3926), .RN(npu_inst_pe_1_3_0_n8), .Q(
        npu_inst_int_data_res_3__0__7_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_0_n100), 
        .CK(npu_inst_pe_1_3_0_net3926), .RN(npu_inst_pe_1_3_0_n8), .Q(
        npu_inst_int_data_res_3__0__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_weight_reg_0_ ( .D(npu_inst_n93), .CK(
        npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n8), .Q(
        npu_inst_pe_1_3_0_int_q_weight_0_), .QN(npu_inst_pe_1_3_0_n27) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_weight_reg_1_ ( .D(npu_inst_n99), .CK(
        npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n8), .Q(
        npu_inst_pe_1_3_0_int_q_weight_1_), .QN(npu_inst_pe_1_3_0_n26) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_0_n112), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n8), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_0_n106), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n8), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_0_n111), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_0_n105), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_0_n110), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_0_n104), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_0_n109), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_0_n103), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_0_n108), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_0_n102), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_0_n107), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_0_n101), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_0_n86), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_0_n87), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n9), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_0_n88), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_0_n89), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_0_n90), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_0_n91), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_0_n92), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_0_n93), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_0_n94), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_0_n95), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_0_n96), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_0_n97), 
        .CK(npu_inst_pe_1_3_0_net3932), .RN(npu_inst_pe_1_3_0_n10), .Q(
        npu_inst_pe_1_3_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_0_net3926) );
  CLKGATETST_X1 npu_inst_pe_1_3_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n46), .SE(1'b0), .GCK(npu_inst_pe_1_3_0_net3932) );
  MUX2_X1 npu_inst_pe_1_3_1_U153 ( .A(npu_inst_pe_1_3_1_n31), .B(
        npu_inst_pe_1_3_1_n28), .S(npu_inst_pe_1_3_1_n7), .Z(
        npu_inst_pe_1_3_1_N93) );
  MUX2_X1 npu_inst_pe_1_3_1_U152 ( .A(npu_inst_pe_1_3_1_n30), .B(
        npu_inst_pe_1_3_1_n29), .S(npu_inst_pe_1_3_1_n5), .Z(
        npu_inst_pe_1_3_1_n31) );
  MUX2_X1 npu_inst_pe_1_3_1_U151 ( .A(npu_inst_pe_1_3_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_1_n3), .Z(
        npu_inst_pe_1_3_1_n30) );
  MUX2_X1 npu_inst_pe_1_3_1_U150 ( .A(npu_inst_pe_1_3_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_1_n3), .Z(
        npu_inst_pe_1_3_1_n29) );
  MUX2_X1 npu_inst_pe_1_3_1_U149 ( .A(npu_inst_pe_1_3_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_1_n3), .Z(
        npu_inst_pe_1_3_1_n28) );
  MUX2_X1 npu_inst_pe_1_3_1_U148 ( .A(npu_inst_pe_1_3_1_n25), .B(
        npu_inst_pe_1_3_1_n22), .S(npu_inst_pe_1_3_1_n7), .Z(
        npu_inst_pe_1_3_1_N94) );
  MUX2_X1 npu_inst_pe_1_3_1_U147 ( .A(npu_inst_pe_1_3_1_n24), .B(
        npu_inst_pe_1_3_1_n23), .S(npu_inst_pe_1_3_1_n5), .Z(
        npu_inst_pe_1_3_1_n25) );
  MUX2_X1 npu_inst_pe_1_3_1_U146 ( .A(npu_inst_pe_1_3_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_1_n3), .Z(
        npu_inst_pe_1_3_1_n24) );
  MUX2_X1 npu_inst_pe_1_3_1_U145 ( .A(npu_inst_pe_1_3_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_1_n3), .Z(
        npu_inst_pe_1_3_1_n23) );
  MUX2_X1 npu_inst_pe_1_3_1_U144 ( .A(npu_inst_pe_1_3_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_1_n3), .Z(
        npu_inst_pe_1_3_1_n22) );
  MUX2_X1 npu_inst_pe_1_3_1_U143 ( .A(npu_inst_pe_1_3_1_n21), .B(
        npu_inst_pe_1_3_1_n18), .S(npu_inst_pe_1_3_1_n7), .Z(
        npu_inst_int_data_x_3__1__1_) );
  MUX2_X1 npu_inst_pe_1_3_1_U142 ( .A(npu_inst_pe_1_3_1_n20), .B(
        npu_inst_pe_1_3_1_n19), .S(npu_inst_pe_1_3_1_n5), .Z(
        npu_inst_pe_1_3_1_n21) );
  MUX2_X1 npu_inst_pe_1_3_1_U141 ( .A(npu_inst_pe_1_3_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_1_n3), .Z(
        npu_inst_pe_1_3_1_n20) );
  MUX2_X1 npu_inst_pe_1_3_1_U140 ( .A(npu_inst_pe_1_3_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_1_n3), .Z(
        npu_inst_pe_1_3_1_n19) );
  MUX2_X1 npu_inst_pe_1_3_1_U139 ( .A(npu_inst_pe_1_3_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_1_n3), .Z(
        npu_inst_pe_1_3_1_n18) );
  MUX2_X1 npu_inst_pe_1_3_1_U138 ( .A(npu_inst_pe_1_3_1_n17), .B(
        npu_inst_pe_1_3_1_n14), .S(npu_inst_pe_1_3_1_n7), .Z(
        npu_inst_int_data_x_3__1__0_) );
  MUX2_X1 npu_inst_pe_1_3_1_U137 ( .A(npu_inst_pe_1_3_1_n16), .B(
        npu_inst_pe_1_3_1_n15), .S(npu_inst_pe_1_3_1_n5), .Z(
        npu_inst_pe_1_3_1_n17) );
  MUX2_X1 npu_inst_pe_1_3_1_U136 ( .A(npu_inst_pe_1_3_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_1_n3), .Z(
        npu_inst_pe_1_3_1_n16) );
  MUX2_X1 npu_inst_pe_1_3_1_U135 ( .A(npu_inst_pe_1_3_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_1_n3), .Z(
        npu_inst_pe_1_3_1_n15) );
  MUX2_X1 npu_inst_pe_1_3_1_U134 ( .A(npu_inst_pe_1_3_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_1_n3), .Z(
        npu_inst_pe_1_3_1_n14) );
  XOR2_X1 npu_inst_pe_1_3_1_U133 ( .A(npu_inst_pe_1_3_1_int_data_0_), .B(
        npu_inst_int_data_res_3__1__0_), .Z(npu_inst_pe_1_3_1_N73) );
  AND2_X1 npu_inst_pe_1_3_1_U132 ( .A1(npu_inst_int_data_res_3__1__0_), .A2(
        npu_inst_pe_1_3_1_int_data_0_), .ZN(npu_inst_pe_1_3_1_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_1_U131 ( .A(npu_inst_int_data_res_3__1__0_), .B(
        npu_inst_pe_1_3_1_n12), .ZN(npu_inst_pe_1_3_1_N65) );
  OR2_X1 npu_inst_pe_1_3_1_U130 ( .A1(npu_inst_pe_1_3_1_n12), .A2(
        npu_inst_int_data_res_3__1__0_), .ZN(npu_inst_pe_1_3_1_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_1_U129 ( .A(npu_inst_int_data_res_3__1__2_), .B(
        npu_inst_pe_1_3_1_add_79_carry_2_), .Z(npu_inst_pe_1_3_1_N75) );
  AND2_X1 npu_inst_pe_1_3_1_U128 ( .A1(npu_inst_pe_1_3_1_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_3__1__2_), .ZN(
        npu_inst_pe_1_3_1_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_1_U127 ( .A(npu_inst_int_data_res_3__1__3_), .B(
        npu_inst_pe_1_3_1_add_79_carry_3_), .Z(npu_inst_pe_1_3_1_N76) );
  AND2_X1 npu_inst_pe_1_3_1_U126 ( .A1(npu_inst_pe_1_3_1_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_3__1__3_), .ZN(
        npu_inst_pe_1_3_1_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_1_U125 ( .A(npu_inst_int_data_res_3__1__4_), .B(
        npu_inst_pe_1_3_1_add_79_carry_4_), .Z(npu_inst_pe_1_3_1_N77) );
  AND2_X1 npu_inst_pe_1_3_1_U124 ( .A1(npu_inst_pe_1_3_1_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_3__1__4_), .ZN(
        npu_inst_pe_1_3_1_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_1_U123 ( .A(npu_inst_int_data_res_3__1__5_), .B(
        npu_inst_pe_1_3_1_add_79_carry_5_), .Z(npu_inst_pe_1_3_1_N78) );
  AND2_X1 npu_inst_pe_1_3_1_U122 ( .A1(npu_inst_pe_1_3_1_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_3__1__5_), .ZN(
        npu_inst_pe_1_3_1_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_1_U121 ( .A(npu_inst_int_data_res_3__1__6_), .B(
        npu_inst_pe_1_3_1_add_79_carry_6_), .Z(npu_inst_pe_1_3_1_N79) );
  AND2_X1 npu_inst_pe_1_3_1_U120 ( .A1(npu_inst_pe_1_3_1_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_3__1__6_), .ZN(
        npu_inst_pe_1_3_1_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_1_U119 ( .A(npu_inst_int_data_res_3__1__7_), .B(
        npu_inst_pe_1_3_1_add_79_carry_7_), .Z(npu_inst_pe_1_3_1_N80) );
  XNOR2_X1 npu_inst_pe_1_3_1_U118 ( .A(npu_inst_pe_1_3_1_sub_77_carry_2_), .B(
        npu_inst_int_data_res_3__1__2_), .ZN(npu_inst_pe_1_3_1_N67) );
  OR2_X1 npu_inst_pe_1_3_1_U117 ( .A1(npu_inst_int_data_res_3__1__2_), .A2(
        npu_inst_pe_1_3_1_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_3_1_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_1_U116 ( .A(npu_inst_pe_1_3_1_sub_77_carry_3_), .B(
        npu_inst_int_data_res_3__1__3_), .ZN(npu_inst_pe_1_3_1_N68) );
  OR2_X1 npu_inst_pe_1_3_1_U115 ( .A1(npu_inst_int_data_res_3__1__3_), .A2(
        npu_inst_pe_1_3_1_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_3_1_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_1_U114 ( .A(npu_inst_pe_1_3_1_sub_77_carry_4_), .B(
        npu_inst_int_data_res_3__1__4_), .ZN(npu_inst_pe_1_3_1_N69) );
  OR2_X1 npu_inst_pe_1_3_1_U113 ( .A1(npu_inst_int_data_res_3__1__4_), .A2(
        npu_inst_pe_1_3_1_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_3_1_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_1_U112 ( .A(npu_inst_pe_1_3_1_sub_77_carry_5_), .B(
        npu_inst_int_data_res_3__1__5_), .ZN(npu_inst_pe_1_3_1_N70) );
  OR2_X1 npu_inst_pe_1_3_1_U111 ( .A1(npu_inst_int_data_res_3__1__5_), .A2(
        npu_inst_pe_1_3_1_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_3_1_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_1_U110 ( .A(npu_inst_pe_1_3_1_sub_77_carry_6_), .B(
        npu_inst_int_data_res_3__1__6_), .ZN(npu_inst_pe_1_3_1_N71) );
  OR2_X1 npu_inst_pe_1_3_1_U109 ( .A1(npu_inst_int_data_res_3__1__6_), .A2(
        npu_inst_pe_1_3_1_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_3_1_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_1_U108 ( .A(npu_inst_int_data_res_3__1__7_), .B(
        npu_inst_pe_1_3_1_sub_77_carry_7_), .ZN(npu_inst_pe_1_3_1_N72) );
  INV_X1 npu_inst_pe_1_3_1_U107 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_3_1_n6)
         );
  INV_X1 npu_inst_pe_1_3_1_U106 ( .A(npu_inst_pe_1_3_1_n6), .ZN(
        npu_inst_pe_1_3_1_n5) );
  INV_X1 npu_inst_pe_1_3_1_U105 ( .A(npu_inst_n39), .ZN(npu_inst_pe_1_3_1_n2)
         );
  AOI22_X1 npu_inst_pe_1_3_1_U104 ( .A1(npu_inst_int_data_y_4__1__0_), .A2(
        npu_inst_pe_1_3_1_n58), .B1(npu_inst_pe_1_3_1_n118), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_1_n57) );
  INV_X1 npu_inst_pe_1_3_1_U103 ( .A(npu_inst_pe_1_3_1_n57), .ZN(
        npu_inst_pe_1_3_1_n107) );
  AOI22_X1 npu_inst_pe_1_3_1_U102 ( .A1(npu_inst_int_data_y_4__1__0_), .A2(
        npu_inst_pe_1_3_1_n54), .B1(npu_inst_pe_1_3_1_n117), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_1_n53) );
  INV_X1 npu_inst_pe_1_3_1_U99 ( .A(npu_inst_pe_1_3_1_n53), .ZN(
        npu_inst_pe_1_3_1_n108) );
  AOI22_X1 npu_inst_pe_1_3_1_U98 ( .A1(npu_inst_int_data_y_4__1__0_), .A2(
        npu_inst_pe_1_3_1_n50), .B1(npu_inst_pe_1_3_1_n116), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_1_n49) );
  INV_X1 npu_inst_pe_1_3_1_U97 ( .A(npu_inst_pe_1_3_1_n49), .ZN(
        npu_inst_pe_1_3_1_n109) );
  AOI22_X1 npu_inst_pe_1_3_1_U96 ( .A1(npu_inst_int_data_y_4__1__0_), .A2(
        npu_inst_pe_1_3_1_n46), .B1(npu_inst_pe_1_3_1_n115), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_1_n45) );
  INV_X1 npu_inst_pe_1_3_1_U95 ( .A(npu_inst_pe_1_3_1_n45), .ZN(
        npu_inst_pe_1_3_1_n110) );
  AOI22_X1 npu_inst_pe_1_3_1_U94 ( .A1(npu_inst_int_data_y_4__1__0_), .A2(
        npu_inst_pe_1_3_1_n42), .B1(npu_inst_pe_1_3_1_n114), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_1_n41) );
  INV_X1 npu_inst_pe_1_3_1_U93 ( .A(npu_inst_pe_1_3_1_n41), .ZN(
        npu_inst_pe_1_3_1_n111) );
  AOI22_X1 npu_inst_pe_1_3_1_U92 ( .A1(npu_inst_int_data_y_4__1__1_), .A2(
        npu_inst_pe_1_3_1_n58), .B1(npu_inst_pe_1_3_1_n118), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_1_n59) );
  INV_X1 npu_inst_pe_1_3_1_U91 ( .A(npu_inst_pe_1_3_1_n59), .ZN(
        npu_inst_pe_1_3_1_n101) );
  AOI22_X1 npu_inst_pe_1_3_1_U90 ( .A1(npu_inst_int_data_y_4__1__1_), .A2(
        npu_inst_pe_1_3_1_n54), .B1(npu_inst_pe_1_3_1_n117), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_1_n55) );
  INV_X1 npu_inst_pe_1_3_1_U89 ( .A(npu_inst_pe_1_3_1_n55), .ZN(
        npu_inst_pe_1_3_1_n102) );
  AOI22_X1 npu_inst_pe_1_3_1_U88 ( .A1(npu_inst_int_data_y_4__1__1_), .A2(
        npu_inst_pe_1_3_1_n50), .B1(npu_inst_pe_1_3_1_n116), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_1_n51) );
  INV_X1 npu_inst_pe_1_3_1_U87 ( .A(npu_inst_pe_1_3_1_n51), .ZN(
        npu_inst_pe_1_3_1_n103) );
  AOI22_X1 npu_inst_pe_1_3_1_U86 ( .A1(npu_inst_int_data_y_4__1__1_), .A2(
        npu_inst_pe_1_3_1_n46), .B1(npu_inst_pe_1_3_1_n115), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_1_n47) );
  INV_X1 npu_inst_pe_1_3_1_U85 ( .A(npu_inst_pe_1_3_1_n47), .ZN(
        npu_inst_pe_1_3_1_n104) );
  AOI22_X1 npu_inst_pe_1_3_1_U84 ( .A1(npu_inst_int_data_y_4__1__1_), .A2(
        npu_inst_pe_1_3_1_n42), .B1(npu_inst_pe_1_3_1_n114), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_1_n43) );
  INV_X1 npu_inst_pe_1_3_1_U83 ( .A(npu_inst_pe_1_3_1_n43), .ZN(
        npu_inst_pe_1_3_1_n105) );
  AOI22_X1 npu_inst_pe_1_3_1_U82 ( .A1(npu_inst_pe_1_3_1_n38), .A2(
        npu_inst_int_data_y_4__1__1_), .B1(npu_inst_pe_1_3_1_n113), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_1_n39) );
  INV_X1 npu_inst_pe_1_3_1_U81 ( .A(npu_inst_pe_1_3_1_n39), .ZN(
        npu_inst_pe_1_3_1_n106) );
  AND2_X1 npu_inst_pe_1_3_1_U80 ( .A1(npu_inst_pe_1_3_1_N93), .A2(npu_inst_n39), .ZN(npu_inst_int_data_y_3__1__0_) );
  NAND2_X1 npu_inst_pe_1_3_1_U79 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_1_n60), .ZN(npu_inst_pe_1_3_1_n74) );
  OAI21_X1 npu_inst_pe_1_3_1_U78 ( .B1(npu_inst_pe_1_3_1_n63), .B2(
        npu_inst_pe_1_3_1_n60), .A(npu_inst_pe_1_3_1_n74), .ZN(
        npu_inst_pe_1_3_1_n97) );
  NAND2_X1 npu_inst_pe_1_3_1_U77 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_1_n60), .ZN(npu_inst_pe_1_3_1_n73) );
  OAI21_X1 npu_inst_pe_1_3_1_U76 ( .B1(npu_inst_pe_1_3_1_n61), .B2(
        npu_inst_pe_1_3_1_n60), .A(npu_inst_pe_1_3_1_n73), .ZN(
        npu_inst_pe_1_3_1_n96) );
  NAND2_X1 npu_inst_pe_1_3_1_U75 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_1_n56), .ZN(npu_inst_pe_1_3_1_n72) );
  OAI21_X1 npu_inst_pe_1_3_1_U74 ( .B1(npu_inst_pe_1_3_1_n63), .B2(
        npu_inst_pe_1_3_1_n56), .A(npu_inst_pe_1_3_1_n72), .ZN(
        npu_inst_pe_1_3_1_n95) );
  NAND2_X1 npu_inst_pe_1_3_1_U73 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_1_n56), .ZN(npu_inst_pe_1_3_1_n71) );
  OAI21_X1 npu_inst_pe_1_3_1_U72 ( .B1(npu_inst_pe_1_3_1_n61), .B2(
        npu_inst_pe_1_3_1_n56), .A(npu_inst_pe_1_3_1_n71), .ZN(
        npu_inst_pe_1_3_1_n94) );
  NAND2_X1 npu_inst_pe_1_3_1_U71 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_1_n52), .ZN(npu_inst_pe_1_3_1_n70) );
  OAI21_X1 npu_inst_pe_1_3_1_U70 ( .B1(npu_inst_pe_1_3_1_n63), .B2(
        npu_inst_pe_1_3_1_n52), .A(npu_inst_pe_1_3_1_n70), .ZN(
        npu_inst_pe_1_3_1_n93) );
  NAND2_X1 npu_inst_pe_1_3_1_U69 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_1_n52), .ZN(npu_inst_pe_1_3_1_n69) );
  OAI21_X1 npu_inst_pe_1_3_1_U68 ( .B1(npu_inst_pe_1_3_1_n61), .B2(
        npu_inst_pe_1_3_1_n52), .A(npu_inst_pe_1_3_1_n69), .ZN(
        npu_inst_pe_1_3_1_n92) );
  NAND2_X1 npu_inst_pe_1_3_1_U67 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_1_n48), .ZN(npu_inst_pe_1_3_1_n68) );
  OAI21_X1 npu_inst_pe_1_3_1_U66 ( .B1(npu_inst_pe_1_3_1_n63), .B2(
        npu_inst_pe_1_3_1_n48), .A(npu_inst_pe_1_3_1_n68), .ZN(
        npu_inst_pe_1_3_1_n91) );
  NAND2_X1 npu_inst_pe_1_3_1_U65 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_1_n48), .ZN(npu_inst_pe_1_3_1_n67) );
  OAI21_X1 npu_inst_pe_1_3_1_U64 ( .B1(npu_inst_pe_1_3_1_n61), .B2(
        npu_inst_pe_1_3_1_n48), .A(npu_inst_pe_1_3_1_n67), .ZN(
        npu_inst_pe_1_3_1_n90) );
  NAND2_X1 npu_inst_pe_1_3_1_U63 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_1_n44), .ZN(npu_inst_pe_1_3_1_n66) );
  OAI21_X1 npu_inst_pe_1_3_1_U62 ( .B1(npu_inst_pe_1_3_1_n63), .B2(
        npu_inst_pe_1_3_1_n44), .A(npu_inst_pe_1_3_1_n66), .ZN(
        npu_inst_pe_1_3_1_n89) );
  NAND2_X1 npu_inst_pe_1_3_1_U61 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_1_n44), .ZN(npu_inst_pe_1_3_1_n65) );
  OAI21_X1 npu_inst_pe_1_3_1_U60 ( .B1(npu_inst_pe_1_3_1_n61), .B2(
        npu_inst_pe_1_3_1_n44), .A(npu_inst_pe_1_3_1_n65), .ZN(
        npu_inst_pe_1_3_1_n88) );
  NAND2_X1 npu_inst_pe_1_3_1_U59 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_1_n40), .ZN(npu_inst_pe_1_3_1_n64) );
  OAI21_X1 npu_inst_pe_1_3_1_U58 ( .B1(npu_inst_pe_1_3_1_n63), .B2(
        npu_inst_pe_1_3_1_n40), .A(npu_inst_pe_1_3_1_n64), .ZN(
        npu_inst_pe_1_3_1_n87) );
  NAND2_X1 npu_inst_pe_1_3_1_U57 ( .A1(npu_inst_pe_1_3_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_1_n40), .ZN(npu_inst_pe_1_3_1_n62) );
  OAI21_X1 npu_inst_pe_1_3_1_U56 ( .B1(npu_inst_pe_1_3_1_n61), .B2(
        npu_inst_pe_1_3_1_n40), .A(npu_inst_pe_1_3_1_n62), .ZN(
        npu_inst_pe_1_3_1_n86) );
  AOI22_X1 npu_inst_pe_1_3_1_U55 ( .A1(npu_inst_pe_1_3_1_n38), .A2(
        npu_inst_int_data_y_4__1__0_), .B1(npu_inst_pe_1_3_1_n113), .B2(
        npu_inst_pe_1_3_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_1_n37) );
  INV_X1 npu_inst_pe_1_3_1_U54 ( .A(npu_inst_pe_1_3_1_n37), .ZN(
        npu_inst_pe_1_3_1_n112) );
  AND2_X1 npu_inst_pe_1_3_1_U53 ( .A1(npu_inst_n39), .A2(npu_inst_pe_1_3_1_N94), .ZN(npu_inst_int_data_y_3__1__1_) );
  AOI222_X1 npu_inst_pe_1_3_1_U52 ( .A1(npu_inst_int_data_res_4__1__0_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N73), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N65), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n84) );
  INV_X1 npu_inst_pe_1_3_1_U51 ( .A(npu_inst_pe_1_3_1_n84), .ZN(
        npu_inst_pe_1_3_1_n100) );
  AOI222_X1 npu_inst_pe_1_3_1_U50 ( .A1(npu_inst_pe_1_3_1_n1), .A2(
        npu_inst_int_data_res_4__1__7_), .B1(npu_inst_pe_1_3_1_N80), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N72), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n75) );
  INV_X1 npu_inst_pe_1_3_1_U49 ( .A(npu_inst_pe_1_3_1_n75), .ZN(
        npu_inst_pe_1_3_1_n32) );
  AOI222_X1 npu_inst_pe_1_3_1_U48 ( .A1(npu_inst_int_data_res_4__1__1_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N74), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N66), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n83) );
  INV_X1 npu_inst_pe_1_3_1_U47 ( .A(npu_inst_pe_1_3_1_n83), .ZN(
        npu_inst_pe_1_3_1_n99) );
  AOI222_X1 npu_inst_pe_1_3_1_U46 ( .A1(npu_inst_int_data_res_4__1__3_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N76), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N68), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n81) );
  INV_X1 npu_inst_pe_1_3_1_U45 ( .A(npu_inst_pe_1_3_1_n81), .ZN(
        npu_inst_pe_1_3_1_n36) );
  AOI222_X1 npu_inst_pe_1_3_1_U44 ( .A1(npu_inst_int_data_res_4__1__4_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N77), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N69), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n80) );
  INV_X1 npu_inst_pe_1_3_1_U43 ( .A(npu_inst_pe_1_3_1_n80), .ZN(
        npu_inst_pe_1_3_1_n35) );
  AOI222_X1 npu_inst_pe_1_3_1_U42 ( .A1(npu_inst_int_data_res_4__1__5_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N78), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N70), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n79) );
  INV_X1 npu_inst_pe_1_3_1_U41 ( .A(npu_inst_pe_1_3_1_n79), .ZN(
        npu_inst_pe_1_3_1_n34) );
  AOI222_X1 npu_inst_pe_1_3_1_U40 ( .A1(npu_inst_int_data_res_4__1__6_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N79), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N71), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n78) );
  INV_X1 npu_inst_pe_1_3_1_U39 ( .A(npu_inst_pe_1_3_1_n78), .ZN(
        npu_inst_pe_1_3_1_n33) );
  AND2_X1 npu_inst_pe_1_3_1_U38 ( .A1(npu_inst_int_data_x_3__1__1_), .A2(
        npu_inst_pe_1_3_1_int_q_weight_1_), .ZN(npu_inst_pe_1_3_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_1_U37 ( .A1(npu_inst_int_data_x_3__1__0_), .A2(
        npu_inst_pe_1_3_1_int_q_weight_1_), .ZN(npu_inst_pe_1_3_1_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_3_1_U36 ( .A(npu_inst_pe_1_3_1_int_data_1_), .ZN(
        npu_inst_pe_1_3_1_n13) );
  NOR3_X1 npu_inst_pe_1_3_1_U35 ( .A1(npu_inst_pe_1_3_1_n26), .A2(npu_inst_n39), .A3(npu_inst_int_ckg[38]), .ZN(npu_inst_pe_1_3_1_n85) );
  OR2_X1 npu_inst_pe_1_3_1_U34 ( .A1(npu_inst_pe_1_3_1_n85), .A2(
        npu_inst_pe_1_3_1_n1), .ZN(npu_inst_pe_1_3_1_N84) );
  AOI222_X1 npu_inst_pe_1_3_1_U33 ( .A1(npu_inst_int_data_res_4__1__2_), .A2(
        npu_inst_pe_1_3_1_n1), .B1(npu_inst_pe_1_3_1_N75), .B2(
        npu_inst_pe_1_3_1_n76), .C1(npu_inst_pe_1_3_1_N67), .C2(
        npu_inst_pe_1_3_1_n77), .ZN(npu_inst_pe_1_3_1_n82) );
  INV_X1 npu_inst_pe_1_3_1_U32 ( .A(npu_inst_pe_1_3_1_n82), .ZN(
        npu_inst_pe_1_3_1_n98) );
  AOI22_X1 npu_inst_pe_1_3_1_U31 ( .A1(npu_inst_n39), .A2(
        npu_inst_int_data_y_4__1__1_), .B1(npu_inst_pe_1_3_1_n2), .B2(
        npu_inst_int_data_x_3__2__1_), .ZN(npu_inst_pe_1_3_1_n63) );
  AOI22_X1 npu_inst_pe_1_3_1_U30 ( .A1(npu_inst_n39), .A2(
        npu_inst_int_data_y_4__1__0_), .B1(npu_inst_pe_1_3_1_n2), .B2(
        npu_inst_int_data_x_3__2__0_), .ZN(npu_inst_pe_1_3_1_n61) );
  INV_X1 npu_inst_pe_1_3_1_U29 ( .A(npu_inst_pe_1_3_1_int_data_0_), .ZN(
        npu_inst_pe_1_3_1_n12) );
  INV_X1 npu_inst_pe_1_3_1_U28 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_3_1_n4)
         );
  OR3_X1 npu_inst_pe_1_3_1_U27 ( .A1(npu_inst_pe_1_3_1_n5), .A2(
        npu_inst_pe_1_3_1_n7), .A3(npu_inst_pe_1_3_1_n4), .ZN(
        npu_inst_pe_1_3_1_n56) );
  OR3_X1 npu_inst_pe_1_3_1_U26 ( .A1(npu_inst_pe_1_3_1_n4), .A2(
        npu_inst_pe_1_3_1_n7), .A3(npu_inst_pe_1_3_1_n6), .ZN(
        npu_inst_pe_1_3_1_n48) );
  INV_X1 npu_inst_pe_1_3_1_U25 ( .A(npu_inst_pe_1_3_1_n4), .ZN(
        npu_inst_pe_1_3_1_n3) );
  OR3_X1 npu_inst_pe_1_3_1_U24 ( .A1(npu_inst_pe_1_3_1_n3), .A2(
        npu_inst_pe_1_3_1_n7), .A3(npu_inst_pe_1_3_1_n6), .ZN(
        npu_inst_pe_1_3_1_n52) );
  OR3_X1 npu_inst_pe_1_3_1_U23 ( .A1(npu_inst_pe_1_3_1_n5), .A2(
        npu_inst_pe_1_3_1_n7), .A3(npu_inst_pe_1_3_1_n3), .ZN(
        npu_inst_pe_1_3_1_n60) );
  BUF_X1 npu_inst_pe_1_3_1_U22 ( .A(npu_inst_n23), .Z(npu_inst_pe_1_3_1_n1) );
  NOR2_X1 npu_inst_pe_1_3_1_U21 ( .A1(npu_inst_pe_1_3_1_n60), .A2(
        npu_inst_pe_1_3_1_n2), .ZN(npu_inst_pe_1_3_1_n58) );
  NOR2_X1 npu_inst_pe_1_3_1_U20 ( .A1(npu_inst_pe_1_3_1_n56), .A2(
        npu_inst_pe_1_3_1_n2), .ZN(npu_inst_pe_1_3_1_n54) );
  NOR2_X1 npu_inst_pe_1_3_1_U19 ( .A1(npu_inst_pe_1_3_1_n52), .A2(
        npu_inst_pe_1_3_1_n2), .ZN(npu_inst_pe_1_3_1_n50) );
  NOR2_X1 npu_inst_pe_1_3_1_U18 ( .A1(npu_inst_pe_1_3_1_n48), .A2(
        npu_inst_pe_1_3_1_n2), .ZN(npu_inst_pe_1_3_1_n46) );
  NOR2_X1 npu_inst_pe_1_3_1_U17 ( .A1(npu_inst_pe_1_3_1_n40), .A2(
        npu_inst_pe_1_3_1_n2), .ZN(npu_inst_pe_1_3_1_n38) );
  NOR2_X1 npu_inst_pe_1_3_1_U16 ( .A1(npu_inst_pe_1_3_1_n44), .A2(
        npu_inst_pe_1_3_1_n2), .ZN(npu_inst_pe_1_3_1_n42) );
  BUF_X1 npu_inst_pe_1_3_1_U15 ( .A(npu_inst_n83), .Z(npu_inst_pe_1_3_1_n7) );
  INV_X1 npu_inst_pe_1_3_1_U14 ( .A(npu_inst_n107), .ZN(npu_inst_pe_1_3_1_n11)
         );
  INV_X1 npu_inst_pe_1_3_1_U13 ( .A(npu_inst_pe_1_3_1_n38), .ZN(
        npu_inst_pe_1_3_1_n113) );
  INV_X1 npu_inst_pe_1_3_1_U12 ( .A(npu_inst_pe_1_3_1_n58), .ZN(
        npu_inst_pe_1_3_1_n118) );
  INV_X1 npu_inst_pe_1_3_1_U11 ( .A(npu_inst_pe_1_3_1_n54), .ZN(
        npu_inst_pe_1_3_1_n117) );
  INV_X1 npu_inst_pe_1_3_1_U10 ( .A(npu_inst_pe_1_3_1_n50), .ZN(
        npu_inst_pe_1_3_1_n116) );
  INV_X1 npu_inst_pe_1_3_1_U9 ( .A(npu_inst_pe_1_3_1_n46), .ZN(
        npu_inst_pe_1_3_1_n115) );
  INV_X1 npu_inst_pe_1_3_1_U8 ( .A(npu_inst_pe_1_3_1_n42), .ZN(
        npu_inst_pe_1_3_1_n114) );
  BUF_X1 npu_inst_pe_1_3_1_U7 ( .A(npu_inst_pe_1_3_1_n11), .Z(
        npu_inst_pe_1_3_1_n10) );
  BUF_X1 npu_inst_pe_1_3_1_U6 ( .A(npu_inst_pe_1_3_1_n11), .Z(
        npu_inst_pe_1_3_1_n9) );
  BUF_X1 npu_inst_pe_1_3_1_U5 ( .A(npu_inst_pe_1_3_1_n11), .Z(
        npu_inst_pe_1_3_1_n8) );
  NOR2_X1 npu_inst_pe_1_3_1_U4 ( .A1(npu_inst_pe_1_3_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_1_n1), .ZN(npu_inst_pe_1_3_1_n76) );
  NOR2_X1 npu_inst_pe_1_3_1_U3 ( .A1(npu_inst_pe_1_3_1_n27), .A2(
        npu_inst_pe_1_3_1_n1), .ZN(npu_inst_pe_1_3_1_n77) );
  FA_X1 npu_inst_pe_1_3_1_sub_77_U2_1 ( .A(npu_inst_int_data_res_3__1__1_), 
        .B(npu_inst_pe_1_3_1_n13), .CI(npu_inst_pe_1_3_1_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_3_1_sub_77_carry_2_), .S(npu_inst_pe_1_3_1_N66) );
  FA_X1 npu_inst_pe_1_3_1_add_79_U1_1 ( .A(npu_inst_int_data_res_3__1__1_), 
        .B(npu_inst_pe_1_3_1_int_data_1_), .CI(
        npu_inst_pe_1_3_1_add_79_carry_1_), .CO(
        npu_inst_pe_1_3_1_add_79_carry_2_), .S(npu_inst_pe_1_3_1_N74) );
  NAND3_X1 npu_inst_pe_1_3_1_U101 ( .A1(npu_inst_pe_1_3_1_n4), .A2(
        npu_inst_pe_1_3_1_n6), .A3(npu_inst_pe_1_3_1_n7), .ZN(
        npu_inst_pe_1_3_1_n44) );
  NAND3_X1 npu_inst_pe_1_3_1_U100 ( .A1(npu_inst_pe_1_3_1_n3), .A2(
        npu_inst_pe_1_3_1_n6), .A3(npu_inst_pe_1_3_1_n7), .ZN(
        npu_inst_pe_1_3_1_n40) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_1_n33), .CK(
        npu_inst_pe_1_3_1_net3903), .RN(npu_inst_pe_1_3_1_n8), .Q(
        npu_inst_int_data_res_3__1__6_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_1_n34), .CK(
        npu_inst_pe_1_3_1_net3903), .RN(npu_inst_pe_1_3_1_n8), .Q(
        npu_inst_int_data_res_3__1__5_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_1_n35), .CK(
        npu_inst_pe_1_3_1_net3903), .RN(npu_inst_pe_1_3_1_n8), .Q(
        npu_inst_int_data_res_3__1__4_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_1_n36), .CK(
        npu_inst_pe_1_3_1_net3903), .RN(npu_inst_pe_1_3_1_n8), .Q(
        npu_inst_int_data_res_3__1__3_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_1_n98), .CK(
        npu_inst_pe_1_3_1_net3903), .RN(npu_inst_pe_1_3_1_n8), .Q(
        npu_inst_int_data_res_3__1__2_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_1_n99), .CK(
        npu_inst_pe_1_3_1_net3903), .RN(npu_inst_pe_1_3_1_n8), .Q(
        npu_inst_int_data_res_3__1__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_1_n32), .CK(
        npu_inst_pe_1_3_1_net3903), .RN(npu_inst_pe_1_3_1_n8), .Q(
        npu_inst_int_data_res_3__1__7_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_1_n100), 
        .CK(npu_inst_pe_1_3_1_net3903), .RN(npu_inst_pe_1_3_1_n8), .Q(
        npu_inst_int_data_res_3__1__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_weight_reg_0_ ( .D(npu_inst_n93), .CK(
        npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n8), .Q(
        npu_inst_pe_1_3_1_int_q_weight_0_), .QN(npu_inst_pe_1_3_1_n27) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_weight_reg_1_ ( .D(npu_inst_n99), .CK(
        npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n8), .Q(
        npu_inst_pe_1_3_1_int_q_weight_1_), .QN(npu_inst_pe_1_3_1_n26) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_1_n112), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n8), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_1_n106), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n8), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_1_n111), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_1_n105), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_1_n110), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_1_n104), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_1_n109), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_1_n103), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_1_n108), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_1_n102), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_1_n107), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_1_n101), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_1_n86), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_1_n87), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n9), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_1_n88), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_1_n89), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_1_n90), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_1_n91), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_1_n92), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_1_n93), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_1_n94), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_1_n95), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_1_n96), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_1_n97), 
        .CK(npu_inst_pe_1_3_1_net3909), .RN(npu_inst_pe_1_3_1_n10), .Q(
        npu_inst_pe_1_3_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_1_net3903) );
  CLKGATETST_X1 npu_inst_pe_1_3_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n46), .SE(1'b0), .GCK(npu_inst_pe_1_3_1_net3909) );
  MUX2_X1 npu_inst_pe_1_3_2_U153 ( .A(npu_inst_pe_1_3_2_n31), .B(
        npu_inst_pe_1_3_2_n28), .S(npu_inst_pe_1_3_2_n7), .Z(
        npu_inst_pe_1_3_2_N93) );
  MUX2_X1 npu_inst_pe_1_3_2_U152 ( .A(npu_inst_pe_1_3_2_n30), .B(
        npu_inst_pe_1_3_2_n29), .S(npu_inst_pe_1_3_2_n5), .Z(
        npu_inst_pe_1_3_2_n31) );
  MUX2_X1 npu_inst_pe_1_3_2_U151 ( .A(npu_inst_pe_1_3_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_2_n3), .Z(
        npu_inst_pe_1_3_2_n30) );
  MUX2_X1 npu_inst_pe_1_3_2_U150 ( .A(npu_inst_pe_1_3_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_2_n3), .Z(
        npu_inst_pe_1_3_2_n29) );
  MUX2_X1 npu_inst_pe_1_3_2_U149 ( .A(npu_inst_pe_1_3_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_2_n3), .Z(
        npu_inst_pe_1_3_2_n28) );
  MUX2_X1 npu_inst_pe_1_3_2_U148 ( .A(npu_inst_pe_1_3_2_n25), .B(
        npu_inst_pe_1_3_2_n22), .S(npu_inst_pe_1_3_2_n7), .Z(
        npu_inst_pe_1_3_2_N94) );
  MUX2_X1 npu_inst_pe_1_3_2_U147 ( .A(npu_inst_pe_1_3_2_n24), .B(
        npu_inst_pe_1_3_2_n23), .S(npu_inst_pe_1_3_2_n5), .Z(
        npu_inst_pe_1_3_2_n25) );
  MUX2_X1 npu_inst_pe_1_3_2_U146 ( .A(npu_inst_pe_1_3_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_2_n3), .Z(
        npu_inst_pe_1_3_2_n24) );
  MUX2_X1 npu_inst_pe_1_3_2_U145 ( .A(npu_inst_pe_1_3_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_2_n3), .Z(
        npu_inst_pe_1_3_2_n23) );
  MUX2_X1 npu_inst_pe_1_3_2_U144 ( .A(npu_inst_pe_1_3_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_2_n3), .Z(
        npu_inst_pe_1_3_2_n22) );
  MUX2_X1 npu_inst_pe_1_3_2_U143 ( .A(npu_inst_pe_1_3_2_n21), .B(
        npu_inst_pe_1_3_2_n18), .S(npu_inst_pe_1_3_2_n7), .Z(
        npu_inst_int_data_x_3__2__1_) );
  MUX2_X1 npu_inst_pe_1_3_2_U142 ( .A(npu_inst_pe_1_3_2_n20), .B(
        npu_inst_pe_1_3_2_n19), .S(npu_inst_pe_1_3_2_n5), .Z(
        npu_inst_pe_1_3_2_n21) );
  MUX2_X1 npu_inst_pe_1_3_2_U141 ( .A(npu_inst_pe_1_3_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_2_n3), .Z(
        npu_inst_pe_1_3_2_n20) );
  MUX2_X1 npu_inst_pe_1_3_2_U140 ( .A(npu_inst_pe_1_3_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_2_n3), .Z(
        npu_inst_pe_1_3_2_n19) );
  MUX2_X1 npu_inst_pe_1_3_2_U139 ( .A(npu_inst_pe_1_3_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_2_n3), .Z(
        npu_inst_pe_1_3_2_n18) );
  MUX2_X1 npu_inst_pe_1_3_2_U138 ( .A(npu_inst_pe_1_3_2_n17), .B(
        npu_inst_pe_1_3_2_n14), .S(npu_inst_pe_1_3_2_n7), .Z(
        npu_inst_int_data_x_3__2__0_) );
  MUX2_X1 npu_inst_pe_1_3_2_U137 ( .A(npu_inst_pe_1_3_2_n16), .B(
        npu_inst_pe_1_3_2_n15), .S(npu_inst_pe_1_3_2_n5), .Z(
        npu_inst_pe_1_3_2_n17) );
  MUX2_X1 npu_inst_pe_1_3_2_U136 ( .A(npu_inst_pe_1_3_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_2_n3), .Z(
        npu_inst_pe_1_3_2_n16) );
  MUX2_X1 npu_inst_pe_1_3_2_U135 ( .A(npu_inst_pe_1_3_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_2_n3), .Z(
        npu_inst_pe_1_3_2_n15) );
  MUX2_X1 npu_inst_pe_1_3_2_U134 ( .A(npu_inst_pe_1_3_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_2_n3), .Z(
        npu_inst_pe_1_3_2_n14) );
  XOR2_X1 npu_inst_pe_1_3_2_U133 ( .A(npu_inst_pe_1_3_2_int_data_0_), .B(
        npu_inst_int_data_res_3__2__0_), .Z(npu_inst_pe_1_3_2_N73) );
  AND2_X1 npu_inst_pe_1_3_2_U132 ( .A1(npu_inst_int_data_res_3__2__0_), .A2(
        npu_inst_pe_1_3_2_int_data_0_), .ZN(npu_inst_pe_1_3_2_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_2_U131 ( .A(npu_inst_int_data_res_3__2__0_), .B(
        npu_inst_pe_1_3_2_n12), .ZN(npu_inst_pe_1_3_2_N65) );
  OR2_X1 npu_inst_pe_1_3_2_U130 ( .A1(npu_inst_pe_1_3_2_n12), .A2(
        npu_inst_int_data_res_3__2__0_), .ZN(npu_inst_pe_1_3_2_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_2_U129 ( .A(npu_inst_int_data_res_3__2__2_), .B(
        npu_inst_pe_1_3_2_add_79_carry_2_), .Z(npu_inst_pe_1_3_2_N75) );
  AND2_X1 npu_inst_pe_1_3_2_U128 ( .A1(npu_inst_pe_1_3_2_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_3__2__2_), .ZN(
        npu_inst_pe_1_3_2_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_2_U127 ( .A(npu_inst_int_data_res_3__2__3_), .B(
        npu_inst_pe_1_3_2_add_79_carry_3_), .Z(npu_inst_pe_1_3_2_N76) );
  AND2_X1 npu_inst_pe_1_3_2_U126 ( .A1(npu_inst_pe_1_3_2_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_3__2__3_), .ZN(
        npu_inst_pe_1_3_2_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_2_U125 ( .A(npu_inst_int_data_res_3__2__4_), .B(
        npu_inst_pe_1_3_2_add_79_carry_4_), .Z(npu_inst_pe_1_3_2_N77) );
  AND2_X1 npu_inst_pe_1_3_2_U124 ( .A1(npu_inst_pe_1_3_2_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_3__2__4_), .ZN(
        npu_inst_pe_1_3_2_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_2_U123 ( .A(npu_inst_int_data_res_3__2__5_), .B(
        npu_inst_pe_1_3_2_add_79_carry_5_), .Z(npu_inst_pe_1_3_2_N78) );
  AND2_X1 npu_inst_pe_1_3_2_U122 ( .A1(npu_inst_pe_1_3_2_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_3__2__5_), .ZN(
        npu_inst_pe_1_3_2_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_2_U121 ( .A(npu_inst_int_data_res_3__2__6_), .B(
        npu_inst_pe_1_3_2_add_79_carry_6_), .Z(npu_inst_pe_1_3_2_N79) );
  AND2_X1 npu_inst_pe_1_3_2_U120 ( .A1(npu_inst_pe_1_3_2_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_3__2__6_), .ZN(
        npu_inst_pe_1_3_2_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_2_U119 ( .A(npu_inst_int_data_res_3__2__7_), .B(
        npu_inst_pe_1_3_2_add_79_carry_7_), .Z(npu_inst_pe_1_3_2_N80) );
  XNOR2_X1 npu_inst_pe_1_3_2_U118 ( .A(npu_inst_pe_1_3_2_sub_77_carry_2_), .B(
        npu_inst_int_data_res_3__2__2_), .ZN(npu_inst_pe_1_3_2_N67) );
  OR2_X1 npu_inst_pe_1_3_2_U117 ( .A1(npu_inst_int_data_res_3__2__2_), .A2(
        npu_inst_pe_1_3_2_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_3_2_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_2_U116 ( .A(npu_inst_pe_1_3_2_sub_77_carry_3_), .B(
        npu_inst_int_data_res_3__2__3_), .ZN(npu_inst_pe_1_3_2_N68) );
  OR2_X1 npu_inst_pe_1_3_2_U115 ( .A1(npu_inst_int_data_res_3__2__3_), .A2(
        npu_inst_pe_1_3_2_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_3_2_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_2_U114 ( .A(npu_inst_pe_1_3_2_sub_77_carry_4_), .B(
        npu_inst_int_data_res_3__2__4_), .ZN(npu_inst_pe_1_3_2_N69) );
  OR2_X1 npu_inst_pe_1_3_2_U113 ( .A1(npu_inst_int_data_res_3__2__4_), .A2(
        npu_inst_pe_1_3_2_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_3_2_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_2_U112 ( .A(npu_inst_pe_1_3_2_sub_77_carry_5_), .B(
        npu_inst_int_data_res_3__2__5_), .ZN(npu_inst_pe_1_3_2_N70) );
  OR2_X1 npu_inst_pe_1_3_2_U111 ( .A1(npu_inst_int_data_res_3__2__5_), .A2(
        npu_inst_pe_1_3_2_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_3_2_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_2_U110 ( .A(npu_inst_pe_1_3_2_sub_77_carry_6_), .B(
        npu_inst_int_data_res_3__2__6_), .ZN(npu_inst_pe_1_3_2_N71) );
  OR2_X1 npu_inst_pe_1_3_2_U109 ( .A1(npu_inst_int_data_res_3__2__6_), .A2(
        npu_inst_pe_1_3_2_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_3_2_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_2_U108 ( .A(npu_inst_int_data_res_3__2__7_), .B(
        npu_inst_pe_1_3_2_sub_77_carry_7_), .ZN(npu_inst_pe_1_3_2_N72) );
  INV_X1 npu_inst_pe_1_3_2_U107 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_3_2_n6)
         );
  INV_X1 npu_inst_pe_1_3_2_U106 ( .A(npu_inst_pe_1_3_2_n6), .ZN(
        npu_inst_pe_1_3_2_n5) );
  INV_X1 npu_inst_pe_1_3_2_U105 ( .A(npu_inst_n39), .ZN(npu_inst_pe_1_3_2_n2)
         );
  AOI22_X1 npu_inst_pe_1_3_2_U104 ( .A1(npu_inst_int_data_y_4__2__0_), .A2(
        npu_inst_pe_1_3_2_n58), .B1(npu_inst_pe_1_3_2_n118), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_2_n57) );
  INV_X1 npu_inst_pe_1_3_2_U103 ( .A(npu_inst_pe_1_3_2_n57), .ZN(
        npu_inst_pe_1_3_2_n107) );
  AOI22_X1 npu_inst_pe_1_3_2_U102 ( .A1(npu_inst_int_data_y_4__2__0_), .A2(
        npu_inst_pe_1_3_2_n54), .B1(npu_inst_pe_1_3_2_n117), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_2_n53) );
  INV_X1 npu_inst_pe_1_3_2_U99 ( .A(npu_inst_pe_1_3_2_n53), .ZN(
        npu_inst_pe_1_3_2_n108) );
  AOI22_X1 npu_inst_pe_1_3_2_U98 ( .A1(npu_inst_int_data_y_4__2__0_), .A2(
        npu_inst_pe_1_3_2_n50), .B1(npu_inst_pe_1_3_2_n116), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_2_n49) );
  INV_X1 npu_inst_pe_1_3_2_U97 ( .A(npu_inst_pe_1_3_2_n49), .ZN(
        npu_inst_pe_1_3_2_n109) );
  AOI22_X1 npu_inst_pe_1_3_2_U96 ( .A1(npu_inst_int_data_y_4__2__0_), .A2(
        npu_inst_pe_1_3_2_n46), .B1(npu_inst_pe_1_3_2_n115), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_2_n45) );
  INV_X1 npu_inst_pe_1_3_2_U95 ( .A(npu_inst_pe_1_3_2_n45), .ZN(
        npu_inst_pe_1_3_2_n110) );
  AOI22_X1 npu_inst_pe_1_3_2_U94 ( .A1(npu_inst_int_data_y_4__2__0_), .A2(
        npu_inst_pe_1_3_2_n42), .B1(npu_inst_pe_1_3_2_n114), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_2_n41) );
  INV_X1 npu_inst_pe_1_3_2_U93 ( .A(npu_inst_pe_1_3_2_n41), .ZN(
        npu_inst_pe_1_3_2_n111) );
  AOI22_X1 npu_inst_pe_1_3_2_U92 ( .A1(npu_inst_int_data_y_4__2__1_), .A2(
        npu_inst_pe_1_3_2_n58), .B1(npu_inst_pe_1_3_2_n118), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_2_n59) );
  INV_X1 npu_inst_pe_1_3_2_U91 ( .A(npu_inst_pe_1_3_2_n59), .ZN(
        npu_inst_pe_1_3_2_n101) );
  AOI22_X1 npu_inst_pe_1_3_2_U90 ( .A1(npu_inst_int_data_y_4__2__1_), .A2(
        npu_inst_pe_1_3_2_n54), .B1(npu_inst_pe_1_3_2_n117), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_2_n55) );
  INV_X1 npu_inst_pe_1_3_2_U89 ( .A(npu_inst_pe_1_3_2_n55), .ZN(
        npu_inst_pe_1_3_2_n102) );
  AOI22_X1 npu_inst_pe_1_3_2_U88 ( .A1(npu_inst_int_data_y_4__2__1_), .A2(
        npu_inst_pe_1_3_2_n50), .B1(npu_inst_pe_1_3_2_n116), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_2_n51) );
  INV_X1 npu_inst_pe_1_3_2_U87 ( .A(npu_inst_pe_1_3_2_n51), .ZN(
        npu_inst_pe_1_3_2_n103) );
  AOI22_X1 npu_inst_pe_1_3_2_U86 ( .A1(npu_inst_int_data_y_4__2__1_), .A2(
        npu_inst_pe_1_3_2_n46), .B1(npu_inst_pe_1_3_2_n115), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_2_n47) );
  INV_X1 npu_inst_pe_1_3_2_U85 ( .A(npu_inst_pe_1_3_2_n47), .ZN(
        npu_inst_pe_1_3_2_n104) );
  AOI22_X1 npu_inst_pe_1_3_2_U84 ( .A1(npu_inst_int_data_y_4__2__1_), .A2(
        npu_inst_pe_1_3_2_n42), .B1(npu_inst_pe_1_3_2_n114), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_2_n43) );
  INV_X1 npu_inst_pe_1_3_2_U83 ( .A(npu_inst_pe_1_3_2_n43), .ZN(
        npu_inst_pe_1_3_2_n105) );
  AOI22_X1 npu_inst_pe_1_3_2_U82 ( .A1(npu_inst_pe_1_3_2_n38), .A2(
        npu_inst_int_data_y_4__2__1_), .B1(npu_inst_pe_1_3_2_n113), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_2_n39) );
  INV_X1 npu_inst_pe_1_3_2_U81 ( .A(npu_inst_pe_1_3_2_n39), .ZN(
        npu_inst_pe_1_3_2_n106) );
  AND2_X1 npu_inst_pe_1_3_2_U80 ( .A1(npu_inst_pe_1_3_2_N93), .A2(npu_inst_n39), .ZN(npu_inst_int_data_y_3__2__0_) );
  NAND2_X1 npu_inst_pe_1_3_2_U79 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_2_n60), .ZN(npu_inst_pe_1_3_2_n74) );
  OAI21_X1 npu_inst_pe_1_3_2_U78 ( .B1(npu_inst_pe_1_3_2_n63), .B2(
        npu_inst_pe_1_3_2_n60), .A(npu_inst_pe_1_3_2_n74), .ZN(
        npu_inst_pe_1_3_2_n97) );
  NAND2_X1 npu_inst_pe_1_3_2_U77 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_2_n60), .ZN(npu_inst_pe_1_3_2_n73) );
  OAI21_X1 npu_inst_pe_1_3_2_U76 ( .B1(npu_inst_pe_1_3_2_n61), .B2(
        npu_inst_pe_1_3_2_n60), .A(npu_inst_pe_1_3_2_n73), .ZN(
        npu_inst_pe_1_3_2_n96) );
  NAND2_X1 npu_inst_pe_1_3_2_U75 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_2_n56), .ZN(npu_inst_pe_1_3_2_n72) );
  OAI21_X1 npu_inst_pe_1_3_2_U74 ( .B1(npu_inst_pe_1_3_2_n63), .B2(
        npu_inst_pe_1_3_2_n56), .A(npu_inst_pe_1_3_2_n72), .ZN(
        npu_inst_pe_1_3_2_n95) );
  NAND2_X1 npu_inst_pe_1_3_2_U73 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_2_n56), .ZN(npu_inst_pe_1_3_2_n71) );
  OAI21_X1 npu_inst_pe_1_3_2_U72 ( .B1(npu_inst_pe_1_3_2_n61), .B2(
        npu_inst_pe_1_3_2_n56), .A(npu_inst_pe_1_3_2_n71), .ZN(
        npu_inst_pe_1_3_2_n94) );
  NAND2_X1 npu_inst_pe_1_3_2_U71 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_2_n52), .ZN(npu_inst_pe_1_3_2_n70) );
  OAI21_X1 npu_inst_pe_1_3_2_U70 ( .B1(npu_inst_pe_1_3_2_n63), .B2(
        npu_inst_pe_1_3_2_n52), .A(npu_inst_pe_1_3_2_n70), .ZN(
        npu_inst_pe_1_3_2_n93) );
  NAND2_X1 npu_inst_pe_1_3_2_U69 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_2_n52), .ZN(npu_inst_pe_1_3_2_n69) );
  OAI21_X1 npu_inst_pe_1_3_2_U68 ( .B1(npu_inst_pe_1_3_2_n61), .B2(
        npu_inst_pe_1_3_2_n52), .A(npu_inst_pe_1_3_2_n69), .ZN(
        npu_inst_pe_1_3_2_n92) );
  NAND2_X1 npu_inst_pe_1_3_2_U67 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_2_n48), .ZN(npu_inst_pe_1_3_2_n68) );
  OAI21_X1 npu_inst_pe_1_3_2_U66 ( .B1(npu_inst_pe_1_3_2_n63), .B2(
        npu_inst_pe_1_3_2_n48), .A(npu_inst_pe_1_3_2_n68), .ZN(
        npu_inst_pe_1_3_2_n91) );
  NAND2_X1 npu_inst_pe_1_3_2_U65 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_2_n48), .ZN(npu_inst_pe_1_3_2_n67) );
  OAI21_X1 npu_inst_pe_1_3_2_U64 ( .B1(npu_inst_pe_1_3_2_n61), .B2(
        npu_inst_pe_1_3_2_n48), .A(npu_inst_pe_1_3_2_n67), .ZN(
        npu_inst_pe_1_3_2_n90) );
  NAND2_X1 npu_inst_pe_1_3_2_U63 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_2_n44), .ZN(npu_inst_pe_1_3_2_n66) );
  OAI21_X1 npu_inst_pe_1_3_2_U62 ( .B1(npu_inst_pe_1_3_2_n63), .B2(
        npu_inst_pe_1_3_2_n44), .A(npu_inst_pe_1_3_2_n66), .ZN(
        npu_inst_pe_1_3_2_n89) );
  NAND2_X1 npu_inst_pe_1_3_2_U61 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_2_n44), .ZN(npu_inst_pe_1_3_2_n65) );
  OAI21_X1 npu_inst_pe_1_3_2_U60 ( .B1(npu_inst_pe_1_3_2_n61), .B2(
        npu_inst_pe_1_3_2_n44), .A(npu_inst_pe_1_3_2_n65), .ZN(
        npu_inst_pe_1_3_2_n88) );
  NAND2_X1 npu_inst_pe_1_3_2_U59 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_2_n40), .ZN(npu_inst_pe_1_3_2_n64) );
  OAI21_X1 npu_inst_pe_1_3_2_U58 ( .B1(npu_inst_pe_1_3_2_n63), .B2(
        npu_inst_pe_1_3_2_n40), .A(npu_inst_pe_1_3_2_n64), .ZN(
        npu_inst_pe_1_3_2_n87) );
  NAND2_X1 npu_inst_pe_1_3_2_U57 ( .A1(npu_inst_pe_1_3_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_2_n40), .ZN(npu_inst_pe_1_3_2_n62) );
  OAI21_X1 npu_inst_pe_1_3_2_U56 ( .B1(npu_inst_pe_1_3_2_n61), .B2(
        npu_inst_pe_1_3_2_n40), .A(npu_inst_pe_1_3_2_n62), .ZN(
        npu_inst_pe_1_3_2_n86) );
  AOI22_X1 npu_inst_pe_1_3_2_U55 ( .A1(npu_inst_pe_1_3_2_n38), .A2(
        npu_inst_int_data_y_4__2__0_), .B1(npu_inst_pe_1_3_2_n113), .B2(
        npu_inst_pe_1_3_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_2_n37) );
  INV_X1 npu_inst_pe_1_3_2_U54 ( .A(npu_inst_pe_1_3_2_n37), .ZN(
        npu_inst_pe_1_3_2_n112) );
  AND2_X1 npu_inst_pe_1_3_2_U53 ( .A1(npu_inst_n39), .A2(npu_inst_pe_1_3_2_N94), .ZN(npu_inst_int_data_y_3__2__1_) );
  AOI222_X1 npu_inst_pe_1_3_2_U52 ( .A1(npu_inst_int_data_res_4__2__0_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N73), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N65), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n84) );
  INV_X1 npu_inst_pe_1_3_2_U51 ( .A(npu_inst_pe_1_3_2_n84), .ZN(
        npu_inst_pe_1_3_2_n100) );
  AOI222_X1 npu_inst_pe_1_3_2_U50 ( .A1(npu_inst_pe_1_3_2_n1), .A2(
        npu_inst_int_data_res_4__2__7_), .B1(npu_inst_pe_1_3_2_N80), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N72), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n75) );
  INV_X1 npu_inst_pe_1_3_2_U49 ( .A(npu_inst_pe_1_3_2_n75), .ZN(
        npu_inst_pe_1_3_2_n32) );
  AOI222_X1 npu_inst_pe_1_3_2_U48 ( .A1(npu_inst_int_data_res_4__2__1_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N74), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N66), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n83) );
  INV_X1 npu_inst_pe_1_3_2_U47 ( .A(npu_inst_pe_1_3_2_n83), .ZN(
        npu_inst_pe_1_3_2_n99) );
  AOI222_X1 npu_inst_pe_1_3_2_U46 ( .A1(npu_inst_int_data_res_4__2__3_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N76), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N68), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n81) );
  INV_X1 npu_inst_pe_1_3_2_U45 ( .A(npu_inst_pe_1_3_2_n81), .ZN(
        npu_inst_pe_1_3_2_n36) );
  AOI222_X1 npu_inst_pe_1_3_2_U44 ( .A1(npu_inst_int_data_res_4__2__4_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N77), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N69), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n80) );
  INV_X1 npu_inst_pe_1_3_2_U43 ( .A(npu_inst_pe_1_3_2_n80), .ZN(
        npu_inst_pe_1_3_2_n35) );
  AOI222_X1 npu_inst_pe_1_3_2_U42 ( .A1(npu_inst_int_data_res_4__2__5_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N78), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N70), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n79) );
  INV_X1 npu_inst_pe_1_3_2_U41 ( .A(npu_inst_pe_1_3_2_n79), .ZN(
        npu_inst_pe_1_3_2_n34) );
  AOI222_X1 npu_inst_pe_1_3_2_U40 ( .A1(npu_inst_int_data_res_4__2__6_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N79), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N71), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n78) );
  INV_X1 npu_inst_pe_1_3_2_U39 ( .A(npu_inst_pe_1_3_2_n78), .ZN(
        npu_inst_pe_1_3_2_n33) );
  AND2_X1 npu_inst_pe_1_3_2_U38 ( .A1(npu_inst_int_data_x_3__2__1_), .A2(
        npu_inst_pe_1_3_2_int_q_weight_1_), .ZN(npu_inst_pe_1_3_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_2_U37 ( .A1(npu_inst_int_data_x_3__2__0_), .A2(
        npu_inst_pe_1_3_2_int_q_weight_1_), .ZN(npu_inst_pe_1_3_2_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_3_2_U36 ( .A(npu_inst_pe_1_3_2_int_data_1_), .ZN(
        npu_inst_pe_1_3_2_n13) );
  NOR3_X1 npu_inst_pe_1_3_2_U35 ( .A1(npu_inst_pe_1_3_2_n26), .A2(npu_inst_n39), .A3(npu_inst_int_ckg[37]), .ZN(npu_inst_pe_1_3_2_n85) );
  OR2_X1 npu_inst_pe_1_3_2_U34 ( .A1(npu_inst_pe_1_3_2_n85), .A2(
        npu_inst_pe_1_3_2_n1), .ZN(npu_inst_pe_1_3_2_N84) );
  AOI222_X1 npu_inst_pe_1_3_2_U33 ( .A1(npu_inst_int_data_res_4__2__2_), .A2(
        npu_inst_pe_1_3_2_n1), .B1(npu_inst_pe_1_3_2_N75), .B2(
        npu_inst_pe_1_3_2_n76), .C1(npu_inst_pe_1_3_2_N67), .C2(
        npu_inst_pe_1_3_2_n77), .ZN(npu_inst_pe_1_3_2_n82) );
  INV_X1 npu_inst_pe_1_3_2_U32 ( .A(npu_inst_pe_1_3_2_n82), .ZN(
        npu_inst_pe_1_3_2_n98) );
  AOI22_X1 npu_inst_pe_1_3_2_U31 ( .A1(npu_inst_n39), .A2(
        npu_inst_int_data_y_4__2__1_), .B1(npu_inst_pe_1_3_2_n2), .B2(
        npu_inst_int_data_x_3__3__1_), .ZN(npu_inst_pe_1_3_2_n63) );
  AOI22_X1 npu_inst_pe_1_3_2_U30 ( .A1(npu_inst_n39), .A2(
        npu_inst_int_data_y_4__2__0_), .B1(npu_inst_pe_1_3_2_n2), .B2(
        npu_inst_int_data_x_3__3__0_), .ZN(npu_inst_pe_1_3_2_n61) );
  INV_X1 npu_inst_pe_1_3_2_U29 ( .A(npu_inst_pe_1_3_2_int_data_0_), .ZN(
        npu_inst_pe_1_3_2_n12) );
  INV_X1 npu_inst_pe_1_3_2_U28 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_3_2_n4)
         );
  OR3_X1 npu_inst_pe_1_3_2_U27 ( .A1(npu_inst_pe_1_3_2_n5), .A2(
        npu_inst_pe_1_3_2_n7), .A3(npu_inst_pe_1_3_2_n4), .ZN(
        npu_inst_pe_1_3_2_n56) );
  OR3_X1 npu_inst_pe_1_3_2_U26 ( .A1(npu_inst_pe_1_3_2_n4), .A2(
        npu_inst_pe_1_3_2_n7), .A3(npu_inst_pe_1_3_2_n6), .ZN(
        npu_inst_pe_1_3_2_n48) );
  INV_X1 npu_inst_pe_1_3_2_U25 ( .A(npu_inst_pe_1_3_2_n4), .ZN(
        npu_inst_pe_1_3_2_n3) );
  OR3_X1 npu_inst_pe_1_3_2_U24 ( .A1(npu_inst_pe_1_3_2_n3), .A2(
        npu_inst_pe_1_3_2_n7), .A3(npu_inst_pe_1_3_2_n6), .ZN(
        npu_inst_pe_1_3_2_n52) );
  OR3_X1 npu_inst_pe_1_3_2_U23 ( .A1(npu_inst_pe_1_3_2_n5), .A2(
        npu_inst_pe_1_3_2_n7), .A3(npu_inst_pe_1_3_2_n3), .ZN(
        npu_inst_pe_1_3_2_n60) );
  BUF_X1 npu_inst_pe_1_3_2_U22 ( .A(npu_inst_n23), .Z(npu_inst_pe_1_3_2_n1) );
  NOR2_X1 npu_inst_pe_1_3_2_U21 ( .A1(npu_inst_pe_1_3_2_n60), .A2(
        npu_inst_pe_1_3_2_n2), .ZN(npu_inst_pe_1_3_2_n58) );
  NOR2_X1 npu_inst_pe_1_3_2_U20 ( .A1(npu_inst_pe_1_3_2_n56), .A2(
        npu_inst_pe_1_3_2_n2), .ZN(npu_inst_pe_1_3_2_n54) );
  NOR2_X1 npu_inst_pe_1_3_2_U19 ( .A1(npu_inst_pe_1_3_2_n52), .A2(
        npu_inst_pe_1_3_2_n2), .ZN(npu_inst_pe_1_3_2_n50) );
  NOR2_X1 npu_inst_pe_1_3_2_U18 ( .A1(npu_inst_pe_1_3_2_n48), .A2(
        npu_inst_pe_1_3_2_n2), .ZN(npu_inst_pe_1_3_2_n46) );
  NOR2_X1 npu_inst_pe_1_3_2_U17 ( .A1(npu_inst_pe_1_3_2_n40), .A2(
        npu_inst_pe_1_3_2_n2), .ZN(npu_inst_pe_1_3_2_n38) );
  NOR2_X1 npu_inst_pe_1_3_2_U16 ( .A1(npu_inst_pe_1_3_2_n44), .A2(
        npu_inst_pe_1_3_2_n2), .ZN(npu_inst_pe_1_3_2_n42) );
  BUF_X1 npu_inst_pe_1_3_2_U15 ( .A(npu_inst_n83), .Z(npu_inst_pe_1_3_2_n7) );
  INV_X1 npu_inst_pe_1_3_2_U14 ( .A(npu_inst_n107), .ZN(npu_inst_pe_1_3_2_n11)
         );
  INV_X1 npu_inst_pe_1_3_2_U13 ( .A(npu_inst_pe_1_3_2_n38), .ZN(
        npu_inst_pe_1_3_2_n113) );
  INV_X1 npu_inst_pe_1_3_2_U12 ( .A(npu_inst_pe_1_3_2_n58), .ZN(
        npu_inst_pe_1_3_2_n118) );
  INV_X1 npu_inst_pe_1_3_2_U11 ( .A(npu_inst_pe_1_3_2_n54), .ZN(
        npu_inst_pe_1_3_2_n117) );
  INV_X1 npu_inst_pe_1_3_2_U10 ( .A(npu_inst_pe_1_3_2_n50), .ZN(
        npu_inst_pe_1_3_2_n116) );
  INV_X1 npu_inst_pe_1_3_2_U9 ( .A(npu_inst_pe_1_3_2_n46), .ZN(
        npu_inst_pe_1_3_2_n115) );
  INV_X1 npu_inst_pe_1_3_2_U8 ( .A(npu_inst_pe_1_3_2_n42), .ZN(
        npu_inst_pe_1_3_2_n114) );
  BUF_X1 npu_inst_pe_1_3_2_U7 ( .A(npu_inst_pe_1_3_2_n11), .Z(
        npu_inst_pe_1_3_2_n10) );
  BUF_X1 npu_inst_pe_1_3_2_U6 ( .A(npu_inst_pe_1_3_2_n11), .Z(
        npu_inst_pe_1_3_2_n9) );
  BUF_X1 npu_inst_pe_1_3_2_U5 ( .A(npu_inst_pe_1_3_2_n11), .Z(
        npu_inst_pe_1_3_2_n8) );
  NOR2_X1 npu_inst_pe_1_3_2_U4 ( .A1(npu_inst_pe_1_3_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_2_n1), .ZN(npu_inst_pe_1_3_2_n76) );
  NOR2_X1 npu_inst_pe_1_3_2_U3 ( .A1(npu_inst_pe_1_3_2_n27), .A2(
        npu_inst_pe_1_3_2_n1), .ZN(npu_inst_pe_1_3_2_n77) );
  FA_X1 npu_inst_pe_1_3_2_sub_77_U2_1 ( .A(npu_inst_int_data_res_3__2__1_), 
        .B(npu_inst_pe_1_3_2_n13), .CI(npu_inst_pe_1_3_2_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_3_2_sub_77_carry_2_), .S(npu_inst_pe_1_3_2_N66) );
  FA_X1 npu_inst_pe_1_3_2_add_79_U1_1 ( .A(npu_inst_int_data_res_3__2__1_), 
        .B(npu_inst_pe_1_3_2_int_data_1_), .CI(
        npu_inst_pe_1_3_2_add_79_carry_1_), .CO(
        npu_inst_pe_1_3_2_add_79_carry_2_), .S(npu_inst_pe_1_3_2_N74) );
  NAND3_X1 npu_inst_pe_1_3_2_U101 ( .A1(npu_inst_pe_1_3_2_n4), .A2(
        npu_inst_pe_1_3_2_n6), .A3(npu_inst_pe_1_3_2_n7), .ZN(
        npu_inst_pe_1_3_2_n44) );
  NAND3_X1 npu_inst_pe_1_3_2_U100 ( .A1(npu_inst_pe_1_3_2_n3), .A2(
        npu_inst_pe_1_3_2_n6), .A3(npu_inst_pe_1_3_2_n7), .ZN(
        npu_inst_pe_1_3_2_n40) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_2_n33), .CK(
        npu_inst_pe_1_3_2_net3880), .RN(npu_inst_pe_1_3_2_n8), .Q(
        npu_inst_int_data_res_3__2__6_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_2_n34), .CK(
        npu_inst_pe_1_3_2_net3880), .RN(npu_inst_pe_1_3_2_n8), .Q(
        npu_inst_int_data_res_3__2__5_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_2_n35), .CK(
        npu_inst_pe_1_3_2_net3880), .RN(npu_inst_pe_1_3_2_n8), .Q(
        npu_inst_int_data_res_3__2__4_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_2_n36), .CK(
        npu_inst_pe_1_3_2_net3880), .RN(npu_inst_pe_1_3_2_n8), .Q(
        npu_inst_int_data_res_3__2__3_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_2_n98), .CK(
        npu_inst_pe_1_3_2_net3880), .RN(npu_inst_pe_1_3_2_n8), .Q(
        npu_inst_int_data_res_3__2__2_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_2_n99), .CK(
        npu_inst_pe_1_3_2_net3880), .RN(npu_inst_pe_1_3_2_n8), .Q(
        npu_inst_int_data_res_3__2__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_2_n32), .CK(
        npu_inst_pe_1_3_2_net3880), .RN(npu_inst_pe_1_3_2_n8), .Q(
        npu_inst_int_data_res_3__2__7_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_2_n100), 
        .CK(npu_inst_pe_1_3_2_net3880), .RN(npu_inst_pe_1_3_2_n8), .Q(
        npu_inst_int_data_res_3__2__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_weight_reg_0_ ( .D(npu_inst_n93), .CK(
        npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n8), .Q(
        npu_inst_pe_1_3_2_int_q_weight_0_), .QN(npu_inst_pe_1_3_2_n27) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_weight_reg_1_ ( .D(npu_inst_n99), .CK(
        npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n8), .Q(
        npu_inst_pe_1_3_2_int_q_weight_1_), .QN(npu_inst_pe_1_3_2_n26) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_2_n112), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n8), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_2_n106), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n8), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_2_n111), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_2_n105), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_2_n110), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_2_n104), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_2_n109), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_2_n103), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_2_n108), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_2_n102), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_2_n107), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_2_n101), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_2_n86), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_2_n87), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n9), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_2_n88), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_2_n89), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_2_n90), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_2_n91), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_2_n92), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_2_n93), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_2_n94), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_2_n95), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_2_n96), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_2_n97), 
        .CK(npu_inst_pe_1_3_2_net3886), .RN(npu_inst_pe_1_3_2_n10), .Q(
        npu_inst_pe_1_3_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_2_net3880) );
  CLKGATETST_X1 npu_inst_pe_1_3_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n46), .SE(1'b0), .GCK(npu_inst_pe_1_3_2_net3886) );
  MUX2_X1 npu_inst_pe_1_3_3_U153 ( .A(npu_inst_pe_1_3_3_n31), .B(
        npu_inst_pe_1_3_3_n28), .S(npu_inst_pe_1_3_3_n7), .Z(
        npu_inst_pe_1_3_3_N93) );
  MUX2_X1 npu_inst_pe_1_3_3_U152 ( .A(npu_inst_pe_1_3_3_n30), .B(
        npu_inst_pe_1_3_3_n29), .S(npu_inst_pe_1_3_3_n5), .Z(
        npu_inst_pe_1_3_3_n31) );
  MUX2_X1 npu_inst_pe_1_3_3_U151 ( .A(npu_inst_pe_1_3_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_3_n3), .Z(
        npu_inst_pe_1_3_3_n30) );
  MUX2_X1 npu_inst_pe_1_3_3_U150 ( .A(npu_inst_pe_1_3_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_3_n3), .Z(
        npu_inst_pe_1_3_3_n29) );
  MUX2_X1 npu_inst_pe_1_3_3_U149 ( .A(npu_inst_pe_1_3_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_3_n3), .Z(
        npu_inst_pe_1_3_3_n28) );
  MUX2_X1 npu_inst_pe_1_3_3_U148 ( .A(npu_inst_pe_1_3_3_n25), .B(
        npu_inst_pe_1_3_3_n22), .S(npu_inst_pe_1_3_3_n7), .Z(
        npu_inst_pe_1_3_3_N94) );
  MUX2_X1 npu_inst_pe_1_3_3_U147 ( .A(npu_inst_pe_1_3_3_n24), .B(
        npu_inst_pe_1_3_3_n23), .S(npu_inst_pe_1_3_3_n5), .Z(
        npu_inst_pe_1_3_3_n25) );
  MUX2_X1 npu_inst_pe_1_3_3_U146 ( .A(npu_inst_pe_1_3_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_3_n3), .Z(
        npu_inst_pe_1_3_3_n24) );
  MUX2_X1 npu_inst_pe_1_3_3_U145 ( .A(npu_inst_pe_1_3_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_3_n3), .Z(
        npu_inst_pe_1_3_3_n23) );
  MUX2_X1 npu_inst_pe_1_3_3_U144 ( .A(npu_inst_pe_1_3_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_3_n3), .Z(
        npu_inst_pe_1_3_3_n22) );
  MUX2_X1 npu_inst_pe_1_3_3_U143 ( .A(npu_inst_pe_1_3_3_n21), .B(
        npu_inst_pe_1_3_3_n18), .S(npu_inst_pe_1_3_3_n7), .Z(
        npu_inst_int_data_x_3__3__1_) );
  MUX2_X1 npu_inst_pe_1_3_3_U142 ( .A(npu_inst_pe_1_3_3_n20), .B(
        npu_inst_pe_1_3_3_n19), .S(npu_inst_pe_1_3_3_n5), .Z(
        npu_inst_pe_1_3_3_n21) );
  MUX2_X1 npu_inst_pe_1_3_3_U141 ( .A(npu_inst_pe_1_3_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_3_n3), .Z(
        npu_inst_pe_1_3_3_n20) );
  MUX2_X1 npu_inst_pe_1_3_3_U140 ( .A(npu_inst_pe_1_3_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_3_n3), .Z(
        npu_inst_pe_1_3_3_n19) );
  MUX2_X1 npu_inst_pe_1_3_3_U139 ( .A(npu_inst_pe_1_3_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_3_n3), .Z(
        npu_inst_pe_1_3_3_n18) );
  MUX2_X1 npu_inst_pe_1_3_3_U138 ( .A(npu_inst_pe_1_3_3_n17), .B(
        npu_inst_pe_1_3_3_n14), .S(npu_inst_pe_1_3_3_n7), .Z(
        npu_inst_int_data_x_3__3__0_) );
  MUX2_X1 npu_inst_pe_1_3_3_U137 ( .A(npu_inst_pe_1_3_3_n16), .B(
        npu_inst_pe_1_3_3_n15), .S(npu_inst_pe_1_3_3_n5), .Z(
        npu_inst_pe_1_3_3_n17) );
  MUX2_X1 npu_inst_pe_1_3_3_U136 ( .A(npu_inst_pe_1_3_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_3_n3), .Z(
        npu_inst_pe_1_3_3_n16) );
  MUX2_X1 npu_inst_pe_1_3_3_U135 ( .A(npu_inst_pe_1_3_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_3_n3), .Z(
        npu_inst_pe_1_3_3_n15) );
  MUX2_X1 npu_inst_pe_1_3_3_U134 ( .A(npu_inst_pe_1_3_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_3_n3), .Z(
        npu_inst_pe_1_3_3_n14) );
  XOR2_X1 npu_inst_pe_1_3_3_U133 ( .A(npu_inst_pe_1_3_3_int_data_0_), .B(
        npu_inst_int_data_res_3__3__0_), .Z(npu_inst_pe_1_3_3_N73) );
  AND2_X1 npu_inst_pe_1_3_3_U132 ( .A1(npu_inst_int_data_res_3__3__0_), .A2(
        npu_inst_pe_1_3_3_int_data_0_), .ZN(npu_inst_pe_1_3_3_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_3_U131 ( .A(npu_inst_int_data_res_3__3__0_), .B(
        npu_inst_pe_1_3_3_n12), .ZN(npu_inst_pe_1_3_3_N65) );
  OR2_X1 npu_inst_pe_1_3_3_U130 ( .A1(npu_inst_pe_1_3_3_n12), .A2(
        npu_inst_int_data_res_3__3__0_), .ZN(npu_inst_pe_1_3_3_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_3_U129 ( .A(npu_inst_int_data_res_3__3__2_), .B(
        npu_inst_pe_1_3_3_add_79_carry_2_), .Z(npu_inst_pe_1_3_3_N75) );
  AND2_X1 npu_inst_pe_1_3_3_U128 ( .A1(npu_inst_pe_1_3_3_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_3__3__2_), .ZN(
        npu_inst_pe_1_3_3_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_3_U127 ( .A(npu_inst_int_data_res_3__3__3_), .B(
        npu_inst_pe_1_3_3_add_79_carry_3_), .Z(npu_inst_pe_1_3_3_N76) );
  AND2_X1 npu_inst_pe_1_3_3_U126 ( .A1(npu_inst_pe_1_3_3_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_3__3__3_), .ZN(
        npu_inst_pe_1_3_3_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_3_U125 ( .A(npu_inst_int_data_res_3__3__4_), .B(
        npu_inst_pe_1_3_3_add_79_carry_4_), .Z(npu_inst_pe_1_3_3_N77) );
  AND2_X1 npu_inst_pe_1_3_3_U124 ( .A1(npu_inst_pe_1_3_3_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_3__3__4_), .ZN(
        npu_inst_pe_1_3_3_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_3_U123 ( .A(npu_inst_int_data_res_3__3__5_), .B(
        npu_inst_pe_1_3_3_add_79_carry_5_), .Z(npu_inst_pe_1_3_3_N78) );
  AND2_X1 npu_inst_pe_1_3_3_U122 ( .A1(npu_inst_pe_1_3_3_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_3__3__5_), .ZN(
        npu_inst_pe_1_3_3_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_3_U121 ( .A(npu_inst_int_data_res_3__3__6_), .B(
        npu_inst_pe_1_3_3_add_79_carry_6_), .Z(npu_inst_pe_1_3_3_N79) );
  AND2_X1 npu_inst_pe_1_3_3_U120 ( .A1(npu_inst_pe_1_3_3_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_3__3__6_), .ZN(
        npu_inst_pe_1_3_3_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_3_U119 ( .A(npu_inst_int_data_res_3__3__7_), .B(
        npu_inst_pe_1_3_3_add_79_carry_7_), .Z(npu_inst_pe_1_3_3_N80) );
  XNOR2_X1 npu_inst_pe_1_3_3_U118 ( .A(npu_inst_pe_1_3_3_sub_77_carry_2_), .B(
        npu_inst_int_data_res_3__3__2_), .ZN(npu_inst_pe_1_3_3_N67) );
  OR2_X1 npu_inst_pe_1_3_3_U117 ( .A1(npu_inst_int_data_res_3__3__2_), .A2(
        npu_inst_pe_1_3_3_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_3_3_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_3_U116 ( .A(npu_inst_pe_1_3_3_sub_77_carry_3_), .B(
        npu_inst_int_data_res_3__3__3_), .ZN(npu_inst_pe_1_3_3_N68) );
  OR2_X1 npu_inst_pe_1_3_3_U115 ( .A1(npu_inst_int_data_res_3__3__3_), .A2(
        npu_inst_pe_1_3_3_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_3_3_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_3_U114 ( .A(npu_inst_pe_1_3_3_sub_77_carry_4_), .B(
        npu_inst_int_data_res_3__3__4_), .ZN(npu_inst_pe_1_3_3_N69) );
  OR2_X1 npu_inst_pe_1_3_3_U113 ( .A1(npu_inst_int_data_res_3__3__4_), .A2(
        npu_inst_pe_1_3_3_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_3_3_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_3_U112 ( .A(npu_inst_pe_1_3_3_sub_77_carry_5_), .B(
        npu_inst_int_data_res_3__3__5_), .ZN(npu_inst_pe_1_3_3_N70) );
  OR2_X1 npu_inst_pe_1_3_3_U111 ( .A1(npu_inst_int_data_res_3__3__5_), .A2(
        npu_inst_pe_1_3_3_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_3_3_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_3_U110 ( .A(npu_inst_pe_1_3_3_sub_77_carry_6_), .B(
        npu_inst_int_data_res_3__3__6_), .ZN(npu_inst_pe_1_3_3_N71) );
  OR2_X1 npu_inst_pe_1_3_3_U109 ( .A1(npu_inst_int_data_res_3__3__6_), .A2(
        npu_inst_pe_1_3_3_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_3_3_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_3_U108 ( .A(npu_inst_int_data_res_3__3__7_), .B(
        npu_inst_pe_1_3_3_sub_77_carry_7_), .ZN(npu_inst_pe_1_3_3_N72) );
  INV_X1 npu_inst_pe_1_3_3_U107 ( .A(npu_inst_n60), .ZN(npu_inst_pe_1_3_3_n6)
         );
  INV_X1 npu_inst_pe_1_3_3_U106 ( .A(npu_inst_pe_1_3_3_n6), .ZN(
        npu_inst_pe_1_3_3_n5) );
  INV_X1 npu_inst_pe_1_3_3_U105 ( .A(npu_inst_n39), .ZN(npu_inst_pe_1_3_3_n2)
         );
  AOI22_X1 npu_inst_pe_1_3_3_U104 ( .A1(npu_inst_int_data_y_4__3__0_), .A2(
        npu_inst_pe_1_3_3_n58), .B1(npu_inst_pe_1_3_3_n118), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_3_n57) );
  INV_X1 npu_inst_pe_1_3_3_U103 ( .A(npu_inst_pe_1_3_3_n57), .ZN(
        npu_inst_pe_1_3_3_n107) );
  AOI22_X1 npu_inst_pe_1_3_3_U102 ( .A1(npu_inst_int_data_y_4__3__0_), .A2(
        npu_inst_pe_1_3_3_n54), .B1(npu_inst_pe_1_3_3_n117), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_3_n53) );
  INV_X1 npu_inst_pe_1_3_3_U99 ( .A(npu_inst_pe_1_3_3_n53), .ZN(
        npu_inst_pe_1_3_3_n108) );
  AOI22_X1 npu_inst_pe_1_3_3_U98 ( .A1(npu_inst_int_data_y_4__3__0_), .A2(
        npu_inst_pe_1_3_3_n50), .B1(npu_inst_pe_1_3_3_n116), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_3_n49) );
  INV_X1 npu_inst_pe_1_3_3_U97 ( .A(npu_inst_pe_1_3_3_n49), .ZN(
        npu_inst_pe_1_3_3_n109) );
  AOI22_X1 npu_inst_pe_1_3_3_U96 ( .A1(npu_inst_int_data_y_4__3__0_), .A2(
        npu_inst_pe_1_3_3_n46), .B1(npu_inst_pe_1_3_3_n115), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_3_n45) );
  INV_X1 npu_inst_pe_1_3_3_U95 ( .A(npu_inst_pe_1_3_3_n45), .ZN(
        npu_inst_pe_1_3_3_n110) );
  AOI22_X1 npu_inst_pe_1_3_3_U94 ( .A1(npu_inst_int_data_y_4__3__0_), .A2(
        npu_inst_pe_1_3_3_n42), .B1(npu_inst_pe_1_3_3_n114), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_3_n41) );
  INV_X1 npu_inst_pe_1_3_3_U93 ( .A(npu_inst_pe_1_3_3_n41), .ZN(
        npu_inst_pe_1_3_3_n111) );
  AOI22_X1 npu_inst_pe_1_3_3_U92 ( .A1(npu_inst_int_data_y_4__3__1_), .A2(
        npu_inst_pe_1_3_3_n58), .B1(npu_inst_pe_1_3_3_n118), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_3_n59) );
  INV_X1 npu_inst_pe_1_3_3_U91 ( .A(npu_inst_pe_1_3_3_n59), .ZN(
        npu_inst_pe_1_3_3_n101) );
  AOI22_X1 npu_inst_pe_1_3_3_U90 ( .A1(npu_inst_int_data_y_4__3__1_), .A2(
        npu_inst_pe_1_3_3_n54), .B1(npu_inst_pe_1_3_3_n117), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_3_n55) );
  INV_X1 npu_inst_pe_1_3_3_U89 ( .A(npu_inst_pe_1_3_3_n55), .ZN(
        npu_inst_pe_1_3_3_n102) );
  AOI22_X1 npu_inst_pe_1_3_3_U88 ( .A1(npu_inst_int_data_y_4__3__1_), .A2(
        npu_inst_pe_1_3_3_n50), .B1(npu_inst_pe_1_3_3_n116), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_3_n51) );
  INV_X1 npu_inst_pe_1_3_3_U87 ( .A(npu_inst_pe_1_3_3_n51), .ZN(
        npu_inst_pe_1_3_3_n103) );
  AOI22_X1 npu_inst_pe_1_3_3_U86 ( .A1(npu_inst_int_data_y_4__3__1_), .A2(
        npu_inst_pe_1_3_3_n46), .B1(npu_inst_pe_1_3_3_n115), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_3_n47) );
  INV_X1 npu_inst_pe_1_3_3_U85 ( .A(npu_inst_pe_1_3_3_n47), .ZN(
        npu_inst_pe_1_3_3_n104) );
  AOI22_X1 npu_inst_pe_1_3_3_U84 ( .A1(npu_inst_int_data_y_4__3__1_), .A2(
        npu_inst_pe_1_3_3_n42), .B1(npu_inst_pe_1_3_3_n114), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_3_n43) );
  INV_X1 npu_inst_pe_1_3_3_U83 ( .A(npu_inst_pe_1_3_3_n43), .ZN(
        npu_inst_pe_1_3_3_n105) );
  AOI22_X1 npu_inst_pe_1_3_3_U82 ( .A1(npu_inst_pe_1_3_3_n38), .A2(
        npu_inst_int_data_y_4__3__1_), .B1(npu_inst_pe_1_3_3_n113), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_3_n39) );
  INV_X1 npu_inst_pe_1_3_3_U81 ( .A(npu_inst_pe_1_3_3_n39), .ZN(
        npu_inst_pe_1_3_3_n106) );
  AND2_X1 npu_inst_pe_1_3_3_U80 ( .A1(npu_inst_pe_1_3_3_N93), .A2(npu_inst_n39), .ZN(npu_inst_int_data_y_3__3__0_) );
  NAND2_X1 npu_inst_pe_1_3_3_U79 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_3_n60), .ZN(npu_inst_pe_1_3_3_n74) );
  OAI21_X1 npu_inst_pe_1_3_3_U78 ( .B1(npu_inst_pe_1_3_3_n63), .B2(
        npu_inst_pe_1_3_3_n60), .A(npu_inst_pe_1_3_3_n74), .ZN(
        npu_inst_pe_1_3_3_n97) );
  NAND2_X1 npu_inst_pe_1_3_3_U77 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_3_n60), .ZN(npu_inst_pe_1_3_3_n73) );
  OAI21_X1 npu_inst_pe_1_3_3_U76 ( .B1(npu_inst_pe_1_3_3_n61), .B2(
        npu_inst_pe_1_3_3_n60), .A(npu_inst_pe_1_3_3_n73), .ZN(
        npu_inst_pe_1_3_3_n96) );
  NAND2_X1 npu_inst_pe_1_3_3_U75 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_3_n56), .ZN(npu_inst_pe_1_3_3_n72) );
  OAI21_X1 npu_inst_pe_1_3_3_U74 ( .B1(npu_inst_pe_1_3_3_n63), .B2(
        npu_inst_pe_1_3_3_n56), .A(npu_inst_pe_1_3_3_n72), .ZN(
        npu_inst_pe_1_3_3_n95) );
  NAND2_X1 npu_inst_pe_1_3_3_U73 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_3_n56), .ZN(npu_inst_pe_1_3_3_n71) );
  OAI21_X1 npu_inst_pe_1_3_3_U72 ( .B1(npu_inst_pe_1_3_3_n61), .B2(
        npu_inst_pe_1_3_3_n56), .A(npu_inst_pe_1_3_3_n71), .ZN(
        npu_inst_pe_1_3_3_n94) );
  NAND2_X1 npu_inst_pe_1_3_3_U71 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_3_n52), .ZN(npu_inst_pe_1_3_3_n70) );
  OAI21_X1 npu_inst_pe_1_3_3_U70 ( .B1(npu_inst_pe_1_3_3_n63), .B2(
        npu_inst_pe_1_3_3_n52), .A(npu_inst_pe_1_3_3_n70), .ZN(
        npu_inst_pe_1_3_3_n93) );
  NAND2_X1 npu_inst_pe_1_3_3_U69 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_3_n52), .ZN(npu_inst_pe_1_3_3_n69) );
  OAI21_X1 npu_inst_pe_1_3_3_U68 ( .B1(npu_inst_pe_1_3_3_n61), .B2(
        npu_inst_pe_1_3_3_n52), .A(npu_inst_pe_1_3_3_n69), .ZN(
        npu_inst_pe_1_3_3_n92) );
  NAND2_X1 npu_inst_pe_1_3_3_U67 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_3_n48), .ZN(npu_inst_pe_1_3_3_n68) );
  OAI21_X1 npu_inst_pe_1_3_3_U66 ( .B1(npu_inst_pe_1_3_3_n63), .B2(
        npu_inst_pe_1_3_3_n48), .A(npu_inst_pe_1_3_3_n68), .ZN(
        npu_inst_pe_1_3_3_n91) );
  NAND2_X1 npu_inst_pe_1_3_3_U65 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_3_n48), .ZN(npu_inst_pe_1_3_3_n67) );
  OAI21_X1 npu_inst_pe_1_3_3_U64 ( .B1(npu_inst_pe_1_3_3_n61), .B2(
        npu_inst_pe_1_3_3_n48), .A(npu_inst_pe_1_3_3_n67), .ZN(
        npu_inst_pe_1_3_3_n90) );
  NAND2_X1 npu_inst_pe_1_3_3_U63 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_3_n44), .ZN(npu_inst_pe_1_3_3_n66) );
  OAI21_X1 npu_inst_pe_1_3_3_U62 ( .B1(npu_inst_pe_1_3_3_n63), .B2(
        npu_inst_pe_1_3_3_n44), .A(npu_inst_pe_1_3_3_n66), .ZN(
        npu_inst_pe_1_3_3_n89) );
  NAND2_X1 npu_inst_pe_1_3_3_U61 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_3_n44), .ZN(npu_inst_pe_1_3_3_n65) );
  OAI21_X1 npu_inst_pe_1_3_3_U60 ( .B1(npu_inst_pe_1_3_3_n61), .B2(
        npu_inst_pe_1_3_3_n44), .A(npu_inst_pe_1_3_3_n65), .ZN(
        npu_inst_pe_1_3_3_n88) );
  NAND2_X1 npu_inst_pe_1_3_3_U59 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_3_n40), .ZN(npu_inst_pe_1_3_3_n64) );
  OAI21_X1 npu_inst_pe_1_3_3_U58 ( .B1(npu_inst_pe_1_3_3_n63), .B2(
        npu_inst_pe_1_3_3_n40), .A(npu_inst_pe_1_3_3_n64), .ZN(
        npu_inst_pe_1_3_3_n87) );
  NAND2_X1 npu_inst_pe_1_3_3_U57 ( .A1(npu_inst_pe_1_3_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_3_n40), .ZN(npu_inst_pe_1_3_3_n62) );
  OAI21_X1 npu_inst_pe_1_3_3_U56 ( .B1(npu_inst_pe_1_3_3_n61), .B2(
        npu_inst_pe_1_3_3_n40), .A(npu_inst_pe_1_3_3_n62), .ZN(
        npu_inst_pe_1_3_3_n86) );
  AOI22_X1 npu_inst_pe_1_3_3_U55 ( .A1(npu_inst_pe_1_3_3_n38), .A2(
        npu_inst_int_data_y_4__3__0_), .B1(npu_inst_pe_1_3_3_n113), .B2(
        npu_inst_pe_1_3_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_3_n37) );
  INV_X1 npu_inst_pe_1_3_3_U54 ( .A(npu_inst_pe_1_3_3_n37), .ZN(
        npu_inst_pe_1_3_3_n112) );
  AND2_X1 npu_inst_pe_1_3_3_U53 ( .A1(npu_inst_n39), .A2(npu_inst_pe_1_3_3_N94), .ZN(npu_inst_int_data_y_3__3__1_) );
  AOI222_X1 npu_inst_pe_1_3_3_U52 ( .A1(npu_inst_int_data_res_4__3__0_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N73), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N65), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n84) );
  INV_X1 npu_inst_pe_1_3_3_U51 ( .A(npu_inst_pe_1_3_3_n84), .ZN(
        npu_inst_pe_1_3_3_n100) );
  AOI222_X1 npu_inst_pe_1_3_3_U50 ( .A1(npu_inst_pe_1_3_3_n1), .A2(
        npu_inst_int_data_res_4__3__7_), .B1(npu_inst_pe_1_3_3_N80), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N72), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n75) );
  INV_X1 npu_inst_pe_1_3_3_U49 ( .A(npu_inst_pe_1_3_3_n75), .ZN(
        npu_inst_pe_1_3_3_n32) );
  AOI222_X1 npu_inst_pe_1_3_3_U48 ( .A1(npu_inst_int_data_res_4__3__1_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N74), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N66), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n83) );
  INV_X1 npu_inst_pe_1_3_3_U47 ( .A(npu_inst_pe_1_3_3_n83), .ZN(
        npu_inst_pe_1_3_3_n99) );
  AOI222_X1 npu_inst_pe_1_3_3_U46 ( .A1(npu_inst_int_data_res_4__3__3_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N76), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N68), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n81) );
  INV_X1 npu_inst_pe_1_3_3_U45 ( .A(npu_inst_pe_1_3_3_n81), .ZN(
        npu_inst_pe_1_3_3_n36) );
  AOI222_X1 npu_inst_pe_1_3_3_U44 ( .A1(npu_inst_int_data_res_4__3__4_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N77), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N69), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n80) );
  INV_X1 npu_inst_pe_1_3_3_U43 ( .A(npu_inst_pe_1_3_3_n80), .ZN(
        npu_inst_pe_1_3_3_n35) );
  AOI222_X1 npu_inst_pe_1_3_3_U42 ( .A1(npu_inst_int_data_res_4__3__5_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N78), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N70), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n79) );
  INV_X1 npu_inst_pe_1_3_3_U41 ( .A(npu_inst_pe_1_3_3_n79), .ZN(
        npu_inst_pe_1_3_3_n34) );
  AOI222_X1 npu_inst_pe_1_3_3_U40 ( .A1(npu_inst_int_data_res_4__3__6_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N79), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N71), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n78) );
  INV_X1 npu_inst_pe_1_3_3_U39 ( .A(npu_inst_pe_1_3_3_n78), .ZN(
        npu_inst_pe_1_3_3_n33) );
  AND2_X1 npu_inst_pe_1_3_3_U38 ( .A1(npu_inst_int_data_x_3__3__1_), .A2(
        npu_inst_pe_1_3_3_int_q_weight_1_), .ZN(npu_inst_pe_1_3_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_3_U37 ( .A1(npu_inst_int_data_x_3__3__0_), .A2(
        npu_inst_pe_1_3_3_int_q_weight_1_), .ZN(npu_inst_pe_1_3_3_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_3_3_U36 ( .A(npu_inst_pe_1_3_3_int_data_1_), .ZN(
        npu_inst_pe_1_3_3_n13) );
  NOR3_X1 npu_inst_pe_1_3_3_U35 ( .A1(npu_inst_pe_1_3_3_n26), .A2(npu_inst_n39), .A3(npu_inst_int_ckg[36]), .ZN(npu_inst_pe_1_3_3_n85) );
  OR2_X1 npu_inst_pe_1_3_3_U34 ( .A1(npu_inst_pe_1_3_3_n85), .A2(
        npu_inst_pe_1_3_3_n1), .ZN(npu_inst_pe_1_3_3_N84) );
  AOI222_X1 npu_inst_pe_1_3_3_U33 ( .A1(npu_inst_int_data_res_4__3__2_), .A2(
        npu_inst_pe_1_3_3_n1), .B1(npu_inst_pe_1_3_3_N75), .B2(
        npu_inst_pe_1_3_3_n76), .C1(npu_inst_pe_1_3_3_N67), .C2(
        npu_inst_pe_1_3_3_n77), .ZN(npu_inst_pe_1_3_3_n82) );
  INV_X1 npu_inst_pe_1_3_3_U32 ( .A(npu_inst_pe_1_3_3_n82), .ZN(
        npu_inst_pe_1_3_3_n98) );
  AOI22_X1 npu_inst_pe_1_3_3_U31 ( .A1(npu_inst_n39), .A2(
        npu_inst_int_data_y_4__3__1_), .B1(npu_inst_pe_1_3_3_n2), .B2(
        npu_inst_int_data_x_3__4__1_), .ZN(npu_inst_pe_1_3_3_n63) );
  AOI22_X1 npu_inst_pe_1_3_3_U30 ( .A1(npu_inst_n39), .A2(
        npu_inst_int_data_y_4__3__0_), .B1(npu_inst_pe_1_3_3_n2), .B2(
        npu_inst_int_data_x_3__4__0_), .ZN(npu_inst_pe_1_3_3_n61) );
  INV_X1 npu_inst_pe_1_3_3_U29 ( .A(npu_inst_pe_1_3_3_int_data_0_), .ZN(
        npu_inst_pe_1_3_3_n12) );
  INV_X1 npu_inst_pe_1_3_3_U28 ( .A(npu_inst_n52), .ZN(npu_inst_pe_1_3_3_n4)
         );
  OR3_X1 npu_inst_pe_1_3_3_U27 ( .A1(npu_inst_pe_1_3_3_n5), .A2(
        npu_inst_pe_1_3_3_n7), .A3(npu_inst_pe_1_3_3_n4), .ZN(
        npu_inst_pe_1_3_3_n56) );
  OR3_X1 npu_inst_pe_1_3_3_U26 ( .A1(npu_inst_pe_1_3_3_n4), .A2(
        npu_inst_pe_1_3_3_n7), .A3(npu_inst_pe_1_3_3_n6), .ZN(
        npu_inst_pe_1_3_3_n48) );
  INV_X1 npu_inst_pe_1_3_3_U25 ( .A(npu_inst_pe_1_3_3_n4), .ZN(
        npu_inst_pe_1_3_3_n3) );
  OR3_X1 npu_inst_pe_1_3_3_U24 ( .A1(npu_inst_pe_1_3_3_n3), .A2(
        npu_inst_pe_1_3_3_n7), .A3(npu_inst_pe_1_3_3_n6), .ZN(
        npu_inst_pe_1_3_3_n52) );
  OR3_X1 npu_inst_pe_1_3_3_U23 ( .A1(npu_inst_pe_1_3_3_n5), .A2(
        npu_inst_pe_1_3_3_n7), .A3(npu_inst_pe_1_3_3_n3), .ZN(
        npu_inst_pe_1_3_3_n60) );
  BUF_X1 npu_inst_pe_1_3_3_U22 ( .A(npu_inst_n23), .Z(npu_inst_pe_1_3_3_n1) );
  NOR2_X1 npu_inst_pe_1_3_3_U21 ( .A1(npu_inst_pe_1_3_3_n60), .A2(
        npu_inst_pe_1_3_3_n2), .ZN(npu_inst_pe_1_3_3_n58) );
  NOR2_X1 npu_inst_pe_1_3_3_U20 ( .A1(npu_inst_pe_1_3_3_n56), .A2(
        npu_inst_pe_1_3_3_n2), .ZN(npu_inst_pe_1_3_3_n54) );
  NOR2_X1 npu_inst_pe_1_3_3_U19 ( .A1(npu_inst_pe_1_3_3_n52), .A2(
        npu_inst_pe_1_3_3_n2), .ZN(npu_inst_pe_1_3_3_n50) );
  NOR2_X1 npu_inst_pe_1_3_3_U18 ( .A1(npu_inst_pe_1_3_3_n48), .A2(
        npu_inst_pe_1_3_3_n2), .ZN(npu_inst_pe_1_3_3_n46) );
  NOR2_X1 npu_inst_pe_1_3_3_U17 ( .A1(npu_inst_pe_1_3_3_n40), .A2(
        npu_inst_pe_1_3_3_n2), .ZN(npu_inst_pe_1_3_3_n38) );
  NOR2_X1 npu_inst_pe_1_3_3_U16 ( .A1(npu_inst_pe_1_3_3_n44), .A2(
        npu_inst_pe_1_3_3_n2), .ZN(npu_inst_pe_1_3_3_n42) );
  BUF_X1 npu_inst_pe_1_3_3_U15 ( .A(npu_inst_n83), .Z(npu_inst_pe_1_3_3_n7) );
  INV_X1 npu_inst_pe_1_3_3_U14 ( .A(npu_inst_n107), .ZN(npu_inst_pe_1_3_3_n11)
         );
  INV_X1 npu_inst_pe_1_3_3_U13 ( .A(npu_inst_pe_1_3_3_n38), .ZN(
        npu_inst_pe_1_3_3_n113) );
  INV_X1 npu_inst_pe_1_3_3_U12 ( .A(npu_inst_pe_1_3_3_n58), .ZN(
        npu_inst_pe_1_3_3_n118) );
  INV_X1 npu_inst_pe_1_3_3_U11 ( .A(npu_inst_pe_1_3_3_n54), .ZN(
        npu_inst_pe_1_3_3_n117) );
  INV_X1 npu_inst_pe_1_3_3_U10 ( .A(npu_inst_pe_1_3_3_n50), .ZN(
        npu_inst_pe_1_3_3_n116) );
  INV_X1 npu_inst_pe_1_3_3_U9 ( .A(npu_inst_pe_1_3_3_n46), .ZN(
        npu_inst_pe_1_3_3_n115) );
  INV_X1 npu_inst_pe_1_3_3_U8 ( .A(npu_inst_pe_1_3_3_n42), .ZN(
        npu_inst_pe_1_3_3_n114) );
  BUF_X1 npu_inst_pe_1_3_3_U7 ( .A(npu_inst_pe_1_3_3_n11), .Z(
        npu_inst_pe_1_3_3_n10) );
  BUF_X1 npu_inst_pe_1_3_3_U6 ( .A(npu_inst_pe_1_3_3_n11), .Z(
        npu_inst_pe_1_3_3_n9) );
  BUF_X1 npu_inst_pe_1_3_3_U5 ( .A(npu_inst_pe_1_3_3_n11), .Z(
        npu_inst_pe_1_3_3_n8) );
  NOR2_X1 npu_inst_pe_1_3_3_U4 ( .A1(npu_inst_pe_1_3_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_3_n1), .ZN(npu_inst_pe_1_3_3_n76) );
  NOR2_X1 npu_inst_pe_1_3_3_U3 ( .A1(npu_inst_pe_1_3_3_n27), .A2(
        npu_inst_pe_1_3_3_n1), .ZN(npu_inst_pe_1_3_3_n77) );
  FA_X1 npu_inst_pe_1_3_3_sub_77_U2_1 ( .A(npu_inst_int_data_res_3__3__1_), 
        .B(npu_inst_pe_1_3_3_n13), .CI(npu_inst_pe_1_3_3_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_3_3_sub_77_carry_2_), .S(npu_inst_pe_1_3_3_N66) );
  FA_X1 npu_inst_pe_1_3_3_add_79_U1_1 ( .A(npu_inst_int_data_res_3__3__1_), 
        .B(npu_inst_pe_1_3_3_int_data_1_), .CI(
        npu_inst_pe_1_3_3_add_79_carry_1_), .CO(
        npu_inst_pe_1_3_3_add_79_carry_2_), .S(npu_inst_pe_1_3_3_N74) );
  NAND3_X1 npu_inst_pe_1_3_3_U101 ( .A1(npu_inst_pe_1_3_3_n4), .A2(
        npu_inst_pe_1_3_3_n6), .A3(npu_inst_pe_1_3_3_n7), .ZN(
        npu_inst_pe_1_3_3_n44) );
  NAND3_X1 npu_inst_pe_1_3_3_U100 ( .A1(npu_inst_pe_1_3_3_n3), .A2(
        npu_inst_pe_1_3_3_n6), .A3(npu_inst_pe_1_3_3_n7), .ZN(
        npu_inst_pe_1_3_3_n40) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_3_n33), .CK(
        npu_inst_pe_1_3_3_net3857), .RN(npu_inst_pe_1_3_3_n8), .Q(
        npu_inst_int_data_res_3__3__6_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_3_n34), .CK(
        npu_inst_pe_1_3_3_net3857), .RN(npu_inst_pe_1_3_3_n8), .Q(
        npu_inst_int_data_res_3__3__5_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_3_n35), .CK(
        npu_inst_pe_1_3_3_net3857), .RN(npu_inst_pe_1_3_3_n8), .Q(
        npu_inst_int_data_res_3__3__4_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_3_n36), .CK(
        npu_inst_pe_1_3_3_net3857), .RN(npu_inst_pe_1_3_3_n8), .Q(
        npu_inst_int_data_res_3__3__3_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_3_n98), .CK(
        npu_inst_pe_1_3_3_net3857), .RN(npu_inst_pe_1_3_3_n8), .Q(
        npu_inst_int_data_res_3__3__2_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_3_n99), .CK(
        npu_inst_pe_1_3_3_net3857), .RN(npu_inst_pe_1_3_3_n8), .Q(
        npu_inst_int_data_res_3__3__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_3_n32), .CK(
        npu_inst_pe_1_3_3_net3857), .RN(npu_inst_pe_1_3_3_n8), .Q(
        npu_inst_int_data_res_3__3__7_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_3_n100), 
        .CK(npu_inst_pe_1_3_3_net3857), .RN(npu_inst_pe_1_3_3_n8), .Q(
        npu_inst_int_data_res_3__3__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_weight_reg_0_ ( .D(npu_inst_n93), .CK(
        npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n8), .Q(
        npu_inst_pe_1_3_3_int_q_weight_0_), .QN(npu_inst_pe_1_3_3_n27) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_weight_reg_1_ ( .D(npu_inst_n99), .CK(
        npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n8), .Q(
        npu_inst_pe_1_3_3_int_q_weight_1_), .QN(npu_inst_pe_1_3_3_n26) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_3_n112), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n8), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_3_n106), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n8), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_3_n111), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_3_n105), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_3_n110), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_3_n104), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_3_n109), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_3_n103), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_3_n108), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_3_n102), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_3_n107), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_3_n101), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_3_n86), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_3_n87), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n9), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_3_n88), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_3_n89), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_3_n90), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_3_n91), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_3_n92), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_3_n93), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_3_n94), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_3_n95), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_3_n96), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_3_n97), 
        .CK(npu_inst_pe_1_3_3_net3863), .RN(npu_inst_pe_1_3_3_n10), .Q(
        npu_inst_pe_1_3_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_3_net3857) );
  CLKGATETST_X1 npu_inst_pe_1_3_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n46), .SE(1'b0), .GCK(npu_inst_pe_1_3_3_net3863) );
  MUX2_X1 npu_inst_pe_1_3_4_U152 ( .A(npu_inst_pe_1_3_4_n30), .B(
        npu_inst_pe_1_3_4_n25), .S(npu_inst_pe_1_3_4_n6), .Z(
        npu_inst_pe_1_3_4_N93) );
  MUX2_X1 npu_inst_pe_1_3_4_U151 ( .A(npu_inst_pe_1_3_4_n29), .B(
        npu_inst_pe_1_3_4_n28), .S(npu_inst_n59), .Z(npu_inst_pe_1_3_4_n30) );
  MUX2_X1 npu_inst_pe_1_3_4_U150 ( .A(npu_inst_pe_1_3_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_4_n3), .Z(
        npu_inst_pe_1_3_4_n29) );
  MUX2_X1 npu_inst_pe_1_3_4_U149 ( .A(npu_inst_pe_1_3_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_4_n3), .Z(
        npu_inst_pe_1_3_4_n28) );
  MUX2_X1 npu_inst_pe_1_3_4_U148 ( .A(npu_inst_pe_1_3_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_4_n3), .Z(
        npu_inst_pe_1_3_4_n25) );
  MUX2_X1 npu_inst_pe_1_3_4_U147 ( .A(npu_inst_pe_1_3_4_n24), .B(
        npu_inst_pe_1_3_4_n21), .S(npu_inst_pe_1_3_4_n6), .Z(
        npu_inst_pe_1_3_4_N94) );
  MUX2_X1 npu_inst_pe_1_3_4_U146 ( .A(npu_inst_pe_1_3_4_n23), .B(
        npu_inst_pe_1_3_4_n22), .S(npu_inst_n59), .Z(npu_inst_pe_1_3_4_n24) );
  MUX2_X1 npu_inst_pe_1_3_4_U145 ( .A(npu_inst_pe_1_3_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_4_n3), .Z(
        npu_inst_pe_1_3_4_n23) );
  MUX2_X1 npu_inst_pe_1_3_4_U144 ( .A(npu_inst_pe_1_3_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_4_n3), .Z(
        npu_inst_pe_1_3_4_n22) );
  MUX2_X1 npu_inst_pe_1_3_4_U143 ( .A(npu_inst_pe_1_3_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_4_n3), .Z(
        npu_inst_pe_1_3_4_n21) );
  MUX2_X1 npu_inst_pe_1_3_4_U142 ( .A(npu_inst_pe_1_3_4_n20), .B(
        npu_inst_pe_1_3_4_n17), .S(npu_inst_pe_1_3_4_n6), .Z(
        npu_inst_int_data_x_3__4__1_) );
  MUX2_X1 npu_inst_pe_1_3_4_U141 ( .A(npu_inst_pe_1_3_4_n19), .B(
        npu_inst_pe_1_3_4_n18), .S(npu_inst_n59), .Z(npu_inst_pe_1_3_4_n20) );
  MUX2_X1 npu_inst_pe_1_3_4_U140 ( .A(npu_inst_pe_1_3_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_4_n3), .Z(
        npu_inst_pe_1_3_4_n19) );
  MUX2_X1 npu_inst_pe_1_3_4_U139 ( .A(npu_inst_pe_1_3_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_4_n3), .Z(
        npu_inst_pe_1_3_4_n18) );
  MUX2_X1 npu_inst_pe_1_3_4_U138 ( .A(npu_inst_pe_1_3_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_4_n3), .Z(
        npu_inst_pe_1_3_4_n17) );
  MUX2_X1 npu_inst_pe_1_3_4_U137 ( .A(npu_inst_pe_1_3_4_n16), .B(
        npu_inst_pe_1_3_4_n13), .S(npu_inst_pe_1_3_4_n6), .Z(
        npu_inst_int_data_x_3__4__0_) );
  MUX2_X1 npu_inst_pe_1_3_4_U136 ( .A(npu_inst_pe_1_3_4_n15), .B(
        npu_inst_pe_1_3_4_n14), .S(npu_inst_n59), .Z(npu_inst_pe_1_3_4_n16) );
  MUX2_X1 npu_inst_pe_1_3_4_U135 ( .A(npu_inst_pe_1_3_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_4_n3), .Z(
        npu_inst_pe_1_3_4_n15) );
  MUX2_X1 npu_inst_pe_1_3_4_U134 ( .A(npu_inst_pe_1_3_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_4_n3), .Z(
        npu_inst_pe_1_3_4_n14) );
  MUX2_X1 npu_inst_pe_1_3_4_U133 ( .A(npu_inst_pe_1_3_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_4_n3), .Z(
        npu_inst_pe_1_3_4_n13) );
  XOR2_X1 npu_inst_pe_1_3_4_U132 ( .A(npu_inst_pe_1_3_4_int_data_0_), .B(
        npu_inst_int_data_res_3__4__0_), .Z(npu_inst_pe_1_3_4_N73) );
  AND2_X1 npu_inst_pe_1_3_4_U131 ( .A1(npu_inst_int_data_res_3__4__0_), .A2(
        npu_inst_pe_1_3_4_int_data_0_), .ZN(npu_inst_pe_1_3_4_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_4_U130 ( .A(npu_inst_int_data_res_3__4__0_), .B(
        npu_inst_pe_1_3_4_n11), .ZN(npu_inst_pe_1_3_4_N65) );
  OR2_X1 npu_inst_pe_1_3_4_U129 ( .A1(npu_inst_pe_1_3_4_n11), .A2(
        npu_inst_int_data_res_3__4__0_), .ZN(npu_inst_pe_1_3_4_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_4_U128 ( .A(npu_inst_int_data_res_3__4__2_), .B(
        npu_inst_pe_1_3_4_add_79_carry_2_), .Z(npu_inst_pe_1_3_4_N75) );
  AND2_X1 npu_inst_pe_1_3_4_U127 ( .A1(npu_inst_pe_1_3_4_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_3__4__2_), .ZN(
        npu_inst_pe_1_3_4_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_4_U126 ( .A(npu_inst_int_data_res_3__4__3_), .B(
        npu_inst_pe_1_3_4_add_79_carry_3_), .Z(npu_inst_pe_1_3_4_N76) );
  AND2_X1 npu_inst_pe_1_3_4_U125 ( .A1(npu_inst_pe_1_3_4_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_3__4__3_), .ZN(
        npu_inst_pe_1_3_4_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_4_U124 ( .A(npu_inst_int_data_res_3__4__4_), .B(
        npu_inst_pe_1_3_4_add_79_carry_4_), .Z(npu_inst_pe_1_3_4_N77) );
  AND2_X1 npu_inst_pe_1_3_4_U123 ( .A1(npu_inst_pe_1_3_4_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_3__4__4_), .ZN(
        npu_inst_pe_1_3_4_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_4_U122 ( .A(npu_inst_int_data_res_3__4__5_), .B(
        npu_inst_pe_1_3_4_add_79_carry_5_), .Z(npu_inst_pe_1_3_4_N78) );
  AND2_X1 npu_inst_pe_1_3_4_U121 ( .A1(npu_inst_pe_1_3_4_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_3__4__5_), .ZN(
        npu_inst_pe_1_3_4_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_4_U120 ( .A(npu_inst_int_data_res_3__4__6_), .B(
        npu_inst_pe_1_3_4_add_79_carry_6_), .Z(npu_inst_pe_1_3_4_N79) );
  AND2_X1 npu_inst_pe_1_3_4_U119 ( .A1(npu_inst_pe_1_3_4_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_3__4__6_), .ZN(
        npu_inst_pe_1_3_4_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_4_U118 ( .A(npu_inst_int_data_res_3__4__7_), .B(
        npu_inst_pe_1_3_4_add_79_carry_7_), .Z(npu_inst_pe_1_3_4_N80) );
  XNOR2_X1 npu_inst_pe_1_3_4_U117 ( .A(npu_inst_pe_1_3_4_sub_77_carry_2_), .B(
        npu_inst_int_data_res_3__4__2_), .ZN(npu_inst_pe_1_3_4_N67) );
  OR2_X1 npu_inst_pe_1_3_4_U116 ( .A1(npu_inst_int_data_res_3__4__2_), .A2(
        npu_inst_pe_1_3_4_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_3_4_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_4_U115 ( .A(npu_inst_pe_1_3_4_sub_77_carry_3_), .B(
        npu_inst_int_data_res_3__4__3_), .ZN(npu_inst_pe_1_3_4_N68) );
  OR2_X1 npu_inst_pe_1_3_4_U114 ( .A1(npu_inst_int_data_res_3__4__3_), .A2(
        npu_inst_pe_1_3_4_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_3_4_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_4_U113 ( .A(npu_inst_pe_1_3_4_sub_77_carry_4_), .B(
        npu_inst_int_data_res_3__4__4_), .ZN(npu_inst_pe_1_3_4_N69) );
  OR2_X1 npu_inst_pe_1_3_4_U112 ( .A1(npu_inst_int_data_res_3__4__4_), .A2(
        npu_inst_pe_1_3_4_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_3_4_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_4_U111 ( .A(npu_inst_pe_1_3_4_sub_77_carry_5_), .B(
        npu_inst_int_data_res_3__4__5_), .ZN(npu_inst_pe_1_3_4_N70) );
  OR2_X1 npu_inst_pe_1_3_4_U110 ( .A1(npu_inst_int_data_res_3__4__5_), .A2(
        npu_inst_pe_1_3_4_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_3_4_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_4_U109 ( .A(npu_inst_pe_1_3_4_sub_77_carry_6_), .B(
        npu_inst_int_data_res_3__4__6_), .ZN(npu_inst_pe_1_3_4_N71) );
  OR2_X1 npu_inst_pe_1_3_4_U108 ( .A1(npu_inst_int_data_res_3__4__6_), .A2(
        npu_inst_pe_1_3_4_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_3_4_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_4_U107 ( .A(npu_inst_int_data_res_3__4__7_), .B(
        npu_inst_pe_1_3_4_sub_77_carry_7_), .ZN(npu_inst_pe_1_3_4_N72) );
  INV_X1 npu_inst_pe_1_3_4_U106 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_3_4_n5)
         );
  INV_X1 npu_inst_pe_1_3_4_U105 ( .A(npu_inst_n39), .ZN(npu_inst_pe_1_3_4_n2)
         );
  AOI22_X1 npu_inst_pe_1_3_4_U104 ( .A1(npu_inst_int_data_y_4__4__0_), .A2(
        npu_inst_pe_1_3_4_n58), .B1(npu_inst_pe_1_3_4_n117), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_4_n57) );
  INV_X1 npu_inst_pe_1_3_4_U103 ( .A(npu_inst_pe_1_3_4_n57), .ZN(
        npu_inst_pe_1_3_4_n106) );
  AOI22_X1 npu_inst_pe_1_3_4_U102 ( .A1(npu_inst_int_data_y_4__4__0_), .A2(
        npu_inst_pe_1_3_4_n54), .B1(npu_inst_pe_1_3_4_n116), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_4_n53) );
  INV_X1 npu_inst_pe_1_3_4_U99 ( .A(npu_inst_pe_1_3_4_n53), .ZN(
        npu_inst_pe_1_3_4_n107) );
  AOI22_X1 npu_inst_pe_1_3_4_U98 ( .A1(npu_inst_int_data_y_4__4__0_), .A2(
        npu_inst_pe_1_3_4_n50), .B1(npu_inst_pe_1_3_4_n115), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_4_n49) );
  INV_X1 npu_inst_pe_1_3_4_U97 ( .A(npu_inst_pe_1_3_4_n49), .ZN(
        npu_inst_pe_1_3_4_n108) );
  AOI22_X1 npu_inst_pe_1_3_4_U96 ( .A1(npu_inst_int_data_y_4__4__0_), .A2(
        npu_inst_pe_1_3_4_n46), .B1(npu_inst_pe_1_3_4_n114), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_4_n45) );
  INV_X1 npu_inst_pe_1_3_4_U95 ( .A(npu_inst_pe_1_3_4_n45), .ZN(
        npu_inst_pe_1_3_4_n109) );
  AOI22_X1 npu_inst_pe_1_3_4_U94 ( .A1(npu_inst_int_data_y_4__4__0_), .A2(
        npu_inst_pe_1_3_4_n42), .B1(npu_inst_pe_1_3_4_n113), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_4_n41) );
  INV_X1 npu_inst_pe_1_3_4_U93 ( .A(npu_inst_pe_1_3_4_n41), .ZN(
        npu_inst_pe_1_3_4_n110) );
  AOI22_X1 npu_inst_pe_1_3_4_U92 ( .A1(npu_inst_int_data_y_4__4__1_), .A2(
        npu_inst_pe_1_3_4_n58), .B1(npu_inst_pe_1_3_4_n117), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_4_n59) );
  INV_X1 npu_inst_pe_1_3_4_U91 ( .A(npu_inst_pe_1_3_4_n59), .ZN(
        npu_inst_pe_1_3_4_n100) );
  AOI22_X1 npu_inst_pe_1_3_4_U90 ( .A1(npu_inst_int_data_y_4__4__1_), .A2(
        npu_inst_pe_1_3_4_n54), .B1(npu_inst_pe_1_3_4_n116), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_4_n55) );
  INV_X1 npu_inst_pe_1_3_4_U89 ( .A(npu_inst_pe_1_3_4_n55), .ZN(
        npu_inst_pe_1_3_4_n101) );
  AOI22_X1 npu_inst_pe_1_3_4_U88 ( .A1(npu_inst_int_data_y_4__4__1_), .A2(
        npu_inst_pe_1_3_4_n50), .B1(npu_inst_pe_1_3_4_n115), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_4_n51) );
  INV_X1 npu_inst_pe_1_3_4_U87 ( .A(npu_inst_pe_1_3_4_n51), .ZN(
        npu_inst_pe_1_3_4_n102) );
  AOI22_X1 npu_inst_pe_1_3_4_U86 ( .A1(npu_inst_int_data_y_4__4__1_), .A2(
        npu_inst_pe_1_3_4_n46), .B1(npu_inst_pe_1_3_4_n114), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_4_n47) );
  INV_X1 npu_inst_pe_1_3_4_U85 ( .A(npu_inst_pe_1_3_4_n47), .ZN(
        npu_inst_pe_1_3_4_n103) );
  AOI22_X1 npu_inst_pe_1_3_4_U84 ( .A1(npu_inst_int_data_y_4__4__1_), .A2(
        npu_inst_pe_1_3_4_n42), .B1(npu_inst_pe_1_3_4_n113), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_4_n43) );
  INV_X1 npu_inst_pe_1_3_4_U83 ( .A(npu_inst_pe_1_3_4_n43), .ZN(
        npu_inst_pe_1_3_4_n104) );
  AOI22_X1 npu_inst_pe_1_3_4_U82 ( .A1(npu_inst_pe_1_3_4_n38), .A2(
        npu_inst_int_data_y_4__4__1_), .B1(npu_inst_pe_1_3_4_n112), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_4_n39) );
  INV_X1 npu_inst_pe_1_3_4_U81 ( .A(npu_inst_pe_1_3_4_n39), .ZN(
        npu_inst_pe_1_3_4_n105) );
  AND2_X1 npu_inst_pe_1_3_4_U80 ( .A1(npu_inst_pe_1_3_4_N93), .A2(npu_inst_n39), .ZN(npu_inst_int_data_y_3__4__0_) );
  NAND2_X1 npu_inst_pe_1_3_4_U79 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_4_n60), .ZN(npu_inst_pe_1_3_4_n74) );
  OAI21_X1 npu_inst_pe_1_3_4_U78 ( .B1(npu_inst_pe_1_3_4_n63), .B2(
        npu_inst_pe_1_3_4_n60), .A(npu_inst_pe_1_3_4_n74), .ZN(
        npu_inst_pe_1_3_4_n97) );
  NAND2_X1 npu_inst_pe_1_3_4_U77 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_4_n60), .ZN(npu_inst_pe_1_3_4_n73) );
  OAI21_X1 npu_inst_pe_1_3_4_U76 ( .B1(npu_inst_pe_1_3_4_n61), .B2(
        npu_inst_pe_1_3_4_n60), .A(npu_inst_pe_1_3_4_n73), .ZN(
        npu_inst_pe_1_3_4_n96) );
  NAND2_X1 npu_inst_pe_1_3_4_U75 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_4_n56), .ZN(npu_inst_pe_1_3_4_n72) );
  OAI21_X1 npu_inst_pe_1_3_4_U74 ( .B1(npu_inst_pe_1_3_4_n63), .B2(
        npu_inst_pe_1_3_4_n56), .A(npu_inst_pe_1_3_4_n72), .ZN(
        npu_inst_pe_1_3_4_n95) );
  NAND2_X1 npu_inst_pe_1_3_4_U73 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_4_n56), .ZN(npu_inst_pe_1_3_4_n71) );
  OAI21_X1 npu_inst_pe_1_3_4_U72 ( .B1(npu_inst_pe_1_3_4_n61), .B2(
        npu_inst_pe_1_3_4_n56), .A(npu_inst_pe_1_3_4_n71), .ZN(
        npu_inst_pe_1_3_4_n94) );
  NAND2_X1 npu_inst_pe_1_3_4_U71 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_4_n52), .ZN(npu_inst_pe_1_3_4_n70) );
  OAI21_X1 npu_inst_pe_1_3_4_U70 ( .B1(npu_inst_pe_1_3_4_n63), .B2(
        npu_inst_pe_1_3_4_n52), .A(npu_inst_pe_1_3_4_n70), .ZN(
        npu_inst_pe_1_3_4_n93) );
  NAND2_X1 npu_inst_pe_1_3_4_U69 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_4_n52), .ZN(npu_inst_pe_1_3_4_n69) );
  OAI21_X1 npu_inst_pe_1_3_4_U68 ( .B1(npu_inst_pe_1_3_4_n61), .B2(
        npu_inst_pe_1_3_4_n52), .A(npu_inst_pe_1_3_4_n69), .ZN(
        npu_inst_pe_1_3_4_n92) );
  NAND2_X1 npu_inst_pe_1_3_4_U67 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_4_n48), .ZN(npu_inst_pe_1_3_4_n68) );
  OAI21_X1 npu_inst_pe_1_3_4_U66 ( .B1(npu_inst_pe_1_3_4_n63), .B2(
        npu_inst_pe_1_3_4_n48), .A(npu_inst_pe_1_3_4_n68), .ZN(
        npu_inst_pe_1_3_4_n91) );
  NAND2_X1 npu_inst_pe_1_3_4_U65 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_4_n48), .ZN(npu_inst_pe_1_3_4_n67) );
  OAI21_X1 npu_inst_pe_1_3_4_U64 ( .B1(npu_inst_pe_1_3_4_n61), .B2(
        npu_inst_pe_1_3_4_n48), .A(npu_inst_pe_1_3_4_n67), .ZN(
        npu_inst_pe_1_3_4_n90) );
  NAND2_X1 npu_inst_pe_1_3_4_U63 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_4_n44), .ZN(npu_inst_pe_1_3_4_n66) );
  OAI21_X1 npu_inst_pe_1_3_4_U62 ( .B1(npu_inst_pe_1_3_4_n63), .B2(
        npu_inst_pe_1_3_4_n44), .A(npu_inst_pe_1_3_4_n66), .ZN(
        npu_inst_pe_1_3_4_n89) );
  NAND2_X1 npu_inst_pe_1_3_4_U61 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_4_n44), .ZN(npu_inst_pe_1_3_4_n65) );
  OAI21_X1 npu_inst_pe_1_3_4_U60 ( .B1(npu_inst_pe_1_3_4_n61), .B2(
        npu_inst_pe_1_3_4_n44), .A(npu_inst_pe_1_3_4_n65), .ZN(
        npu_inst_pe_1_3_4_n88) );
  NAND2_X1 npu_inst_pe_1_3_4_U59 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_4_n40), .ZN(npu_inst_pe_1_3_4_n64) );
  OAI21_X1 npu_inst_pe_1_3_4_U58 ( .B1(npu_inst_pe_1_3_4_n63), .B2(
        npu_inst_pe_1_3_4_n40), .A(npu_inst_pe_1_3_4_n64), .ZN(
        npu_inst_pe_1_3_4_n87) );
  NAND2_X1 npu_inst_pe_1_3_4_U57 ( .A1(npu_inst_pe_1_3_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_4_n40), .ZN(npu_inst_pe_1_3_4_n62) );
  OAI21_X1 npu_inst_pe_1_3_4_U56 ( .B1(npu_inst_pe_1_3_4_n61), .B2(
        npu_inst_pe_1_3_4_n40), .A(npu_inst_pe_1_3_4_n62), .ZN(
        npu_inst_pe_1_3_4_n86) );
  AOI22_X1 npu_inst_pe_1_3_4_U55 ( .A1(npu_inst_pe_1_3_4_n38), .A2(
        npu_inst_int_data_y_4__4__0_), .B1(npu_inst_pe_1_3_4_n112), .B2(
        npu_inst_pe_1_3_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_4_n37) );
  INV_X1 npu_inst_pe_1_3_4_U54 ( .A(npu_inst_pe_1_3_4_n37), .ZN(
        npu_inst_pe_1_3_4_n111) );
  AND2_X1 npu_inst_pe_1_3_4_U53 ( .A1(npu_inst_n39), .A2(npu_inst_pe_1_3_4_N94), .ZN(npu_inst_int_data_y_3__4__1_) );
  AOI222_X1 npu_inst_pe_1_3_4_U52 ( .A1(npu_inst_int_data_res_4__4__0_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N73), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N65), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n84) );
  INV_X1 npu_inst_pe_1_3_4_U51 ( .A(npu_inst_pe_1_3_4_n84), .ZN(
        npu_inst_pe_1_3_4_n99) );
  AOI222_X1 npu_inst_pe_1_3_4_U50 ( .A1(npu_inst_pe_1_3_4_n1), .A2(
        npu_inst_int_data_res_4__4__7_), .B1(npu_inst_pe_1_3_4_N80), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N72), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n75) );
  INV_X1 npu_inst_pe_1_3_4_U49 ( .A(npu_inst_pe_1_3_4_n75), .ZN(
        npu_inst_pe_1_3_4_n31) );
  AOI222_X1 npu_inst_pe_1_3_4_U48 ( .A1(npu_inst_int_data_res_4__4__1_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N74), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N66), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n83) );
  INV_X1 npu_inst_pe_1_3_4_U47 ( .A(npu_inst_pe_1_3_4_n83), .ZN(
        npu_inst_pe_1_3_4_n98) );
  AOI222_X1 npu_inst_pe_1_3_4_U46 ( .A1(npu_inst_int_data_res_4__4__3_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N76), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N68), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n81) );
  INV_X1 npu_inst_pe_1_3_4_U45 ( .A(npu_inst_pe_1_3_4_n81), .ZN(
        npu_inst_pe_1_3_4_n35) );
  AOI222_X1 npu_inst_pe_1_3_4_U44 ( .A1(npu_inst_int_data_res_4__4__4_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N77), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N69), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n80) );
  INV_X1 npu_inst_pe_1_3_4_U43 ( .A(npu_inst_pe_1_3_4_n80), .ZN(
        npu_inst_pe_1_3_4_n34) );
  AOI222_X1 npu_inst_pe_1_3_4_U42 ( .A1(npu_inst_int_data_res_4__4__5_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N78), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N70), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n79) );
  INV_X1 npu_inst_pe_1_3_4_U41 ( .A(npu_inst_pe_1_3_4_n79), .ZN(
        npu_inst_pe_1_3_4_n33) );
  AOI222_X1 npu_inst_pe_1_3_4_U40 ( .A1(npu_inst_int_data_res_4__4__6_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N79), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N71), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n78) );
  INV_X1 npu_inst_pe_1_3_4_U39 ( .A(npu_inst_pe_1_3_4_n78), .ZN(
        npu_inst_pe_1_3_4_n32) );
  AND2_X1 npu_inst_pe_1_3_4_U38 ( .A1(npu_inst_int_data_x_3__4__1_), .A2(
        npu_inst_pe_1_3_4_int_q_weight_1_), .ZN(npu_inst_pe_1_3_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_4_U37 ( .A1(npu_inst_int_data_x_3__4__0_), .A2(
        npu_inst_pe_1_3_4_int_q_weight_1_), .ZN(npu_inst_pe_1_3_4_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_3_4_U36 ( .A(npu_inst_pe_1_3_4_int_data_1_), .ZN(
        npu_inst_pe_1_3_4_n12) );
  NOR3_X1 npu_inst_pe_1_3_4_U35 ( .A1(npu_inst_pe_1_3_4_n26), .A2(npu_inst_n39), .A3(npu_inst_int_ckg[35]), .ZN(npu_inst_pe_1_3_4_n85) );
  OR2_X1 npu_inst_pe_1_3_4_U34 ( .A1(npu_inst_pe_1_3_4_n85), .A2(
        npu_inst_pe_1_3_4_n1), .ZN(npu_inst_pe_1_3_4_N84) );
  AOI222_X1 npu_inst_pe_1_3_4_U33 ( .A1(npu_inst_int_data_res_4__4__2_), .A2(
        npu_inst_pe_1_3_4_n1), .B1(npu_inst_pe_1_3_4_N75), .B2(
        npu_inst_pe_1_3_4_n76), .C1(npu_inst_pe_1_3_4_N67), .C2(
        npu_inst_pe_1_3_4_n77), .ZN(npu_inst_pe_1_3_4_n82) );
  INV_X1 npu_inst_pe_1_3_4_U32 ( .A(npu_inst_pe_1_3_4_n82), .ZN(
        npu_inst_pe_1_3_4_n36) );
  AOI22_X1 npu_inst_pe_1_3_4_U31 ( .A1(npu_inst_n39), .A2(
        npu_inst_int_data_y_4__4__1_), .B1(npu_inst_pe_1_3_4_n2), .B2(
        npu_inst_int_data_x_3__5__1_), .ZN(npu_inst_pe_1_3_4_n63) );
  AOI22_X1 npu_inst_pe_1_3_4_U30 ( .A1(npu_inst_n39), .A2(
        npu_inst_int_data_y_4__4__0_), .B1(npu_inst_pe_1_3_4_n2), .B2(
        npu_inst_int_data_x_3__5__0_), .ZN(npu_inst_pe_1_3_4_n61) );
  INV_X1 npu_inst_pe_1_3_4_U29 ( .A(npu_inst_pe_1_3_4_int_data_0_), .ZN(
        npu_inst_pe_1_3_4_n11) );
  INV_X1 npu_inst_pe_1_3_4_U28 ( .A(npu_inst_n51), .ZN(npu_inst_pe_1_3_4_n4)
         );
  OR3_X1 npu_inst_pe_1_3_4_U27 ( .A1(npu_inst_n59), .A2(npu_inst_pe_1_3_4_n6), 
        .A3(npu_inst_pe_1_3_4_n4), .ZN(npu_inst_pe_1_3_4_n56) );
  OR3_X1 npu_inst_pe_1_3_4_U26 ( .A1(npu_inst_pe_1_3_4_n4), .A2(
        npu_inst_pe_1_3_4_n6), .A3(npu_inst_pe_1_3_4_n5), .ZN(
        npu_inst_pe_1_3_4_n48) );
  INV_X1 npu_inst_pe_1_3_4_U25 ( .A(npu_inst_pe_1_3_4_n4), .ZN(
        npu_inst_pe_1_3_4_n3) );
  OR3_X1 npu_inst_pe_1_3_4_U24 ( .A1(npu_inst_pe_1_3_4_n3), .A2(
        npu_inst_pe_1_3_4_n6), .A3(npu_inst_pe_1_3_4_n5), .ZN(
        npu_inst_pe_1_3_4_n52) );
  OR3_X1 npu_inst_pe_1_3_4_U23 ( .A1(npu_inst_n59), .A2(npu_inst_pe_1_3_4_n6), 
        .A3(npu_inst_pe_1_3_4_n3), .ZN(npu_inst_pe_1_3_4_n60) );
  BUF_X1 npu_inst_pe_1_3_4_U22 ( .A(npu_inst_n22), .Z(npu_inst_pe_1_3_4_n1) );
  NOR2_X1 npu_inst_pe_1_3_4_U21 ( .A1(npu_inst_pe_1_3_4_n60), .A2(
        npu_inst_pe_1_3_4_n2), .ZN(npu_inst_pe_1_3_4_n58) );
  NOR2_X1 npu_inst_pe_1_3_4_U20 ( .A1(npu_inst_pe_1_3_4_n56), .A2(
        npu_inst_pe_1_3_4_n2), .ZN(npu_inst_pe_1_3_4_n54) );
  NOR2_X1 npu_inst_pe_1_3_4_U19 ( .A1(npu_inst_pe_1_3_4_n52), .A2(
        npu_inst_pe_1_3_4_n2), .ZN(npu_inst_pe_1_3_4_n50) );
  NOR2_X1 npu_inst_pe_1_3_4_U18 ( .A1(npu_inst_pe_1_3_4_n48), .A2(
        npu_inst_pe_1_3_4_n2), .ZN(npu_inst_pe_1_3_4_n46) );
  NOR2_X1 npu_inst_pe_1_3_4_U17 ( .A1(npu_inst_pe_1_3_4_n40), .A2(
        npu_inst_pe_1_3_4_n2), .ZN(npu_inst_pe_1_3_4_n38) );
  NOR2_X1 npu_inst_pe_1_3_4_U16 ( .A1(npu_inst_pe_1_3_4_n44), .A2(
        npu_inst_pe_1_3_4_n2), .ZN(npu_inst_pe_1_3_4_n42) );
  BUF_X1 npu_inst_pe_1_3_4_U15 ( .A(npu_inst_n82), .Z(npu_inst_pe_1_3_4_n6) );
  INV_X1 npu_inst_pe_1_3_4_U14 ( .A(npu_inst_n106), .ZN(npu_inst_pe_1_3_4_n10)
         );
  INV_X1 npu_inst_pe_1_3_4_U13 ( .A(npu_inst_pe_1_3_4_n38), .ZN(
        npu_inst_pe_1_3_4_n112) );
  INV_X1 npu_inst_pe_1_3_4_U12 ( .A(npu_inst_pe_1_3_4_n58), .ZN(
        npu_inst_pe_1_3_4_n117) );
  INV_X1 npu_inst_pe_1_3_4_U11 ( .A(npu_inst_pe_1_3_4_n54), .ZN(
        npu_inst_pe_1_3_4_n116) );
  INV_X1 npu_inst_pe_1_3_4_U10 ( .A(npu_inst_pe_1_3_4_n50), .ZN(
        npu_inst_pe_1_3_4_n115) );
  INV_X1 npu_inst_pe_1_3_4_U9 ( .A(npu_inst_pe_1_3_4_n46), .ZN(
        npu_inst_pe_1_3_4_n114) );
  INV_X1 npu_inst_pe_1_3_4_U8 ( .A(npu_inst_pe_1_3_4_n42), .ZN(
        npu_inst_pe_1_3_4_n113) );
  BUF_X1 npu_inst_pe_1_3_4_U7 ( .A(npu_inst_pe_1_3_4_n10), .Z(
        npu_inst_pe_1_3_4_n9) );
  BUF_X1 npu_inst_pe_1_3_4_U6 ( .A(npu_inst_pe_1_3_4_n10), .Z(
        npu_inst_pe_1_3_4_n8) );
  BUF_X1 npu_inst_pe_1_3_4_U5 ( .A(npu_inst_pe_1_3_4_n10), .Z(
        npu_inst_pe_1_3_4_n7) );
  NOR2_X1 npu_inst_pe_1_3_4_U4 ( .A1(npu_inst_pe_1_3_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_4_n1), .ZN(npu_inst_pe_1_3_4_n76) );
  NOR2_X1 npu_inst_pe_1_3_4_U3 ( .A1(npu_inst_pe_1_3_4_n27), .A2(
        npu_inst_pe_1_3_4_n1), .ZN(npu_inst_pe_1_3_4_n77) );
  FA_X1 npu_inst_pe_1_3_4_sub_77_U2_1 ( .A(npu_inst_int_data_res_3__4__1_), 
        .B(npu_inst_pe_1_3_4_n12), .CI(npu_inst_pe_1_3_4_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_3_4_sub_77_carry_2_), .S(npu_inst_pe_1_3_4_N66) );
  FA_X1 npu_inst_pe_1_3_4_add_79_U1_1 ( .A(npu_inst_int_data_res_3__4__1_), 
        .B(npu_inst_pe_1_3_4_int_data_1_), .CI(
        npu_inst_pe_1_3_4_add_79_carry_1_), .CO(
        npu_inst_pe_1_3_4_add_79_carry_2_), .S(npu_inst_pe_1_3_4_N74) );
  NAND3_X1 npu_inst_pe_1_3_4_U101 ( .A1(npu_inst_pe_1_3_4_n4), .A2(
        npu_inst_pe_1_3_4_n5), .A3(npu_inst_pe_1_3_4_n6), .ZN(
        npu_inst_pe_1_3_4_n44) );
  NAND3_X1 npu_inst_pe_1_3_4_U100 ( .A1(npu_inst_pe_1_3_4_n3), .A2(
        npu_inst_pe_1_3_4_n5), .A3(npu_inst_pe_1_3_4_n6), .ZN(
        npu_inst_pe_1_3_4_n40) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_4_n32), .CK(
        npu_inst_pe_1_3_4_net3834), .RN(npu_inst_pe_1_3_4_n7), .Q(
        npu_inst_int_data_res_3__4__6_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_4_n33), .CK(
        npu_inst_pe_1_3_4_net3834), .RN(npu_inst_pe_1_3_4_n7), .Q(
        npu_inst_int_data_res_3__4__5_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_4_n34), .CK(
        npu_inst_pe_1_3_4_net3834), .RN(npu_inst_pe_1_3_4_n7), .Q(
        npu_inst_int_data_res_3__4__4_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_4_n35), .CK(
        npu_inst_pe_1_3_4_net3834), .RN(npu_inst_pe_1_3_4_n7), .Q(
        npu_inst_int_data_res_3__4__3_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_4_n36), .CK(
        npu_inst_pe_1_3_4_net3834), .RN(npu_inst_pe_1_3_4_n7), .Q(
        npu_inst_int_data_res_3__4__2_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_4_n98), .CK(
        npu_inst_pe_1_3_4_net3834), .RN(npu_inst_pe_1_3_4_n7), .Q(
        npu_inst_int_data_res_3__4__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_4_n31), .CK(
        npu_inst_pe_1_3_4_net3834), .RN(npu_inst_pe_1_3_4_n7), .Q(
        npu_inst_int_data_res_3__4__7_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_4_n99), .CK(
        npu_inst_pe_1_3_4_net3834), .RN(npu_inst_pe_1_3_4_n7), .Q(
        npu_inst_int_data_res_3__4__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_weight_reg_0_ ( .D(npu_inst_n92), .CK(
        npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n7), .Q(
        npu_inst_pe_1_3_4_int_q_weight_0_), .QN(npu_inst_pe_1_3_4_n27) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_weight_reg_1_ ( .D(npu_inst_n98), .CK(
        npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n7), .Q(
        npu_inst_pe_1_3_4_int_q_weight_1_), .QN(npu_inst_pe_1_3_4_n26) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_4_n111), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n7), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_4_n105), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n7), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_4_n110), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_4_n104), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_4_n109), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_4_n103), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_4_n108), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_4_n102), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_4_n107), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_4_n101), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_4_n106), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_4_n100), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_4_n86), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_4_n87), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n8), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_4_n88), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_4_n89), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_4_n90), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_4_n91), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_4_n92), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_4_n93), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_4_n94), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_4_n95), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_4_n96), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_4_n97), 
        .CK(npu_inst_pe_1_3_4_net3840), .RN(npu_inst_pe_1_3_4_n9), .Q(
        npu_inst_pe_1_3_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_4_net3834) );
  CLKGATETST_X1 npu_inst_pe_1_3_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n46), .SE(1'b0), .GCK(npu_inst_pe_1_3_4_net3840) );
  MUX2_X1 npu_inst_pe_1_3_5_U153 ( .A(npu_inst_pe_1_3_5_n31), .B(
        npu_inst_pe_1_3_5_n28), .S(npu_inst_pe_1_3_5_n7), .Z(
        npu_inst_pe_1_3_5_N93) );
  MUX2_X1 npu_inst_pe_1_3_5_U152 ( .A(npu_inst_pe_1_3_5_n30), .B(
        npu_inst_pe_1_3_5_n29), .S(npu_inst_pe_1_3_5_n5), .Z(
        npu_inst_pe_1_3_5_n31) );
  MUX2_X1 npu_inst_pe_1_3_5_U151 ( .A(npu_inst_pe_1_3_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_5_n3), .Z(
        npu_inst_pe_1_3_5_n30) );
  MUX2_X1 npu_inst_pe_1_3_5_U150 ( .A(npu_inst_pe_1_3_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_5_n3), .Z(
        npu_inst_pe_1_3_5_n29) );
  MUX2_X1 npu_inst_pe_1_3_5_U149 ( .A(npu_inst_pe_1_3_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_5_n3), .Z(
        npu_inst_pe_1_3_5_n28) );
  MUX2_X1 npu_inst_pe_1_3_5_U148 ( .A(npu_inst_pe_1_3_5_n25), .B(
        npu_inst_pe_1_3_5_n22), .S(npu_inst_pe_1_3_5_n7), .Z(
        npu_inst_pe_1_3_5_N94) );
  MUX2_X1 npu_inst_pe_1_3_5_U147 ( .A(npu_inst_pe_1_3_5_n24), .B(
        npu_inst_pe_1_3_5_n23), .S(npu_inst_pe_1_3_5_n5), .Z(
        npu_inst_pe_1_3_5_n25) );
  MUX2_X1 npu_inst_pe_1_3_5_U146 ( .A(npu_inst_pe_1_3_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_5_n3), .Z(
        npu_inst_pe_1_3_5_n24) );
  MUX2_X1 npu_inst_pe_1_3_5_U145 ( .A(npu_inst_pe_1_3_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_5_n3), .Z(
        npu_inst_pe_1_3_5_n23) );
  MUX2_X1 npu_inst_pe_1_3_5_U144 ( .A(npu_inst_pe_1_3_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_5_n3), .Z(
        npu_inst_pe_1_3_5_n22) );
  MUX2_X1 npu_inst_pe_1_3_5_U143 ( .A(npu_inst_pe_1_3_5_n21), .B(
        npu_inst_pe_1_3_5_n18), .S(npu_inst_pe_1_3_5_n7), .Z(
        npu_inst_int_data_x_3__5__1_) );
  MUX2_X1 npu_inst_pe_1_3_5_U142 ( .A(npu_inst_pe_1_3_5_n20), .B(
        npu_inst_pe_1_3_5_n19), .S(npu_inst_pe_1_3_5_n5), .Z(
        npu_inst_pe_1_3_5_n21) );
  MUX2_X1 npu_inst_pe_1_3_5_U141 ( .A(npu_inst_pe_1_3_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_5_n3), .Z(
        npu_inst_pe_1_3_5_n20) );
  MUX2_X1 npu_inst_pe_1_3_5_U140 ( .A(npu_inst_pe_1_3_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_5_n3), .Z(
        npu_inst_pe_1_3_5_n19) );
  MUX2_X1 npu_inst_pe_1_3_5_U139 ( .A(npu_inst_pe_1_3_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_5_n3), .Z(
        npu_inst_pe_1_3_5_n18) );
  MUX2_X1 npu_inst_pe_1_3_5_U138 ( .A(npu_inst_pe_1_3_5_n17), .B(
        npu_inst_pe_1_3_5_n14), .S(npu_inst_pe_1_3_5_n7), .Z(
        npu_inst_int_data_x_3__5__0_) );
  MUX2_X1 npu_inst_pe_1_3_5_U137 ( .A(npu_inst_pe_1_3_5_n16), .B(
        npu_inst_pe_1_3_5_n15), .S(npu_inst_pe_1_3_5_n5), .Z(
        npu_inst_pe_1_3_5_n17) );
  MUX2_X1 npu_inst_pe_1_3_5_U136 ( .A(npu_inst_pe_1_3_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_5_n3), .Z(
        npu_inst_pe_1_3_5_n16) );
  MUX2_X1 npu_inst_pe_1_3_5_U135 ( .A(npu_inst_pe_1_3_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_5_n3), .Z(
        npu_inst_pe_1_3_5_n15) );
  MUX2_X1 npu_inst_pe_1_3_5_U134 ( .A(npu_inst_pe_1_3_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_5_n3), .Z(
        npu_inst_pe_1_3_5_n14) );
  XOR2_X1 npu_inst_pe_1_3_5_U133 ( .A(npu_inst_pe_1_3_5_int_data_0_), .B(
        npu_inst_int_data_res_3__5__0_), .Z(npu_inst_pe_1_3_5_N73) );
  AND2_X1 npu_inst_pe_1_3_5_U132 ( .A1(npu_inst_int_data_res_3__5__0_), .A2(
        npu_inst_pe_1_3_5_int_data_0_), .ZN(npu_inst_pe_1_3_5_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_5_U131 ( .A(npu_inst_int_data_res_3__5__0_), .B(
        npu_inst_pe_1_3_5_n12), .ZN(npu_inst_pe_1_3_5_N65) );
  OR2_X1 npu_inst_pe_1_3_5_U130 ( .A1(npu_inst_pe_1_3_5_n12), .A2(
        npu_inst_int_data_res_3__5__0_), .ZN(npu_inst_pe_1_3_5_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_5_U129 ( .A(npu_inst_int_data_res_3__5__2_), .B(
        npu_inst_pe_1_3_5_add_79_carry_2_), .Z(npu_inst_pe_1_3_5_N75) );
  AND2_X1 npu_inst_pe_1_3_5_U128 ( .A1(npu_inst_pe_1_3_5_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_3__5__2_), .ZN(
        npu_inst_pe_1_3_5_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_5_U127 ( .A(npu_inst_int_data_res_3__5__3_), .B(
        npu_inst_pe_1_3_5_add_79_carry_3_), .Z(npu_inst_pe_1_3_5_N76) );
  AND2_X1 npu_inst_pe_1_3_5_U126 ( .A1(npu_inst_pe_1_3_5_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_3__5__3_), .ZN(
        npu_inst_pe_1_3_5_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_5_U125 ( .A(npu_inst_int_data_res_3__5__4_), .B(
        npu_inst_pe_1_3_5_add_79_carry_4_), .Z(npu_inst_pe_1_3_5_N77) );
  AND2_X1 npu_inst_pe_1_3_5_U124 ( .A1(npu_inst_pe_1_3_5_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_3__5__4_), .ZN(
        npu_inst_pe_1_3_5_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_5_U123 ( .A(npu_inst_int_data_res_3__5__5_), .B(
        npu_inst_pe_1_3_5_add_79_carry_5_), .Z(npu_inst_pe_1_3_5_N78) );
  AND2_X1 npu_inst_pe_1_3_5_U122 ( .A1(npu_inst_pe_1_3_5_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_3__5__5_), .ZN(
        npu_inst_pe_1_3_5_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_5_U121 ( .A(npu_inst_int_data_res_3__5__6_), .B(
        npu_inst_pe_1_3_5_add_79_carry_6_), .Z(npu_inst_pe_1_3_5_N79) );
  AND2_X1 npu_inst_pe_1_3_5_U120 ( .A1(npu_inst_pe_1_3_5_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_3__5__6_), .ZN(
        npu_inst_pe_1_3_5_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_5_U119 ( .A(npu_inst_int_data_res_3__5__7_), .B(
        npu_inst_pe_1_3_5_add_79_carry_7_), .Z(npu_inst_pe_1_3_5_N80) );
  XNOR2_X1 npu_inst_pe_1_3_5_U118 ( .A(npu_inst_pe_1_3_5_sub_77_carry_2_), .B(
        npu_inst_int_data_res_3__5__2_), .ZN(npu_inst_pe_1_3_5_N67) );
  OR2_X1 npu_inst_pe_1_3_5_U117 ( .A1(npu_inst_int_data_res_3__5__2_), .A2(
        npu_inst_pe_1_3_5_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_3_5_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_5_U116 ( .A(npu_inst_pe_1_3_5_sub_77_carry_3_), .B(
        npu_inst_int_data_res_3__5__3_), .ZN(npu_inst_pe_1_3_5_N68) );
  OR2_X1 npu_inst_pe_1_3_5_U115 ( .A1(npu_inst_int_data_res_3__5__3_), .A2(
        npu_inst_pe_1_3_5_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_3_5_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_5_U114 ( .A(npu_inst_pe_1_3_5_sub_77_carry_4_), .B(
        npu_inst_int_data_res_3__5__4_), .ZN(npu_inst_pe_1_3_5_N69) );
  OR2_X1 npu_inst_pe_1_3_5_U113 ( .A1(npu_inst_int_data_res_3__5__4_), .A2(
        npu_inst_pe_1_3_5_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_3_5_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_5_U112 ( .A(npu_inst_pe_1_3_5_sub_77_carry_5_), .B(
        npu_inst_int_data_res_3__5__5_), .ZN(npu_inst_pe_1_3_5_N70) );
  OR2_X1 npu_inst_pe_1_3_5_U111 ( .A1(npu_inst_int_data_res_3__5__5_), .A2(
        npu_inst_pe_1_3_5_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_3_5_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_5_U110 ( .A(npu_inst_pe_1_3_5_sub_77_carry_6_), .B(
        npu_inst_int_data_res_3__5__6_), .ZN(npu_inst_pe_1_3_5_N71) );
  OR2_X1 npu_inst_pe_1_3_5_U109 ( .A1(npu_inst_int_data_res_3__5__6_), .A2(
        npu_inst_pe_1_3_5_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_3_5_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_5_U108 ( .A(npu_inst_int_data_res_3__5__7_), .B(
        npu_inst_pe_1_3_5_sub_77_carry_7_), .ZN(npu_inst_pe_1_3_5_N72) );
  INV_X1 npu_inst_pe_1_3_5_U107 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_3_5_n6)
         );
  INV_X1 npu_inst_pe_1_3_5_U106 ( .A(npu_inst_pe_1_3_5_n6), .ZN(
        npu_inst_pe_1_3_5_n5) );
  INV_X1 npu_inst_pe_1_3_5_U105 ( .A(npu_inst_n38), .ZN(npu_inst_pe_1_3_5_n2)
         );
  AOI22_X1 npu_inst_pe_1_3_5_U104 ( .A1(npu_inst_int_data_y_4__5__0_), .A2(
        npu_inst_pe_1_3_5_n58), .B1(npu_inst_pe_1_3_5_n118), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_5_n57) );
  INV_X1 npu_inst_pe_1_3_5_U103 ( .A(npu_inst_pe_1_3_5_n57), .ZN(
        npu_inst_pe_1_3_5_n107) );
  AOI22_X1 npu_inst_pe_1_3_5_U102 ( .A1(npu_inst_int_data_y_4__5__0_), .A2(
        npu_inst_pe_1_3_5_n54), .B1(npu_inst_pe_1_3_5_n117), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_5_n53) );
  INV_X1 npu_inst_pe_1_3_5_U99 ( .A(npu_inst_pe_1_3_5_n53), .ZN(
        npu_inst_pe_1_3_5_n108) );
  AOI22_X1 npu_inst_pe_1_3_5_U98 ( .A1(npu_inst_int_data_y_4__5__0_), .A2(
        npu_inst_pe_1_3_5_n50), .B1(npu_inst_pe_1_3_5_n116), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_5_n49) );
  INV_X1 npu_inst_pe_1_3_5_U97 ( .A(npu_inst_pe_1_3_5_n49), .ZN(
        npu_inst_pe_1_3_5_n109) );
  AOI22_X1 npu_inst_pe_1_3_5_U96 ( .A1(npu_inst_int_data_y_4__5__0_), .A2(
        npu_inst_pe_1_3_5_n46), .B1(npu_inst_pe_1_3_5_n115), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_5_n45) );
  INV_X1 npu_inst_pe_1_3_5_U95 ( .A(npu_inst_pe_1_3_5_n45), .ZN(
        npu_inst_pe_1_3_5_n110) );
  AOI22_X1 npu_inst_pe_1_3_5_U94 ( .A1(npu_inst_int_data_y_4__5__0_), .A2(
        npu_inst_pe_1_3_5_n42), .B1(npu_inst_pe_1_3_5_n114), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_5_n41) );
  INV_X1 npu_inst_pe_1_3_5_U93 ( .A(npu_inst_pe_1_3_5_n41), .ZN(
        npu_inst_pe_1_3_5_n111) );
  AOI22_X1 npu_inst_pe_1_3_5_U92 ( .A1(npu_inst_int_data_y_4__5__1_), .A2(
        npu_inst_pe_1_3_5_n58), .B1(npu_inst_pe_1_3_5_n118), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_5_n59) );
  INV_X1 npu_inst_pe_1_3_5_U91 ( .A(npu_inst_pe_1_3_5_n59), .ZN(
        npu_inst_pe_1_3_5_n101) );
  AOI22_X1 npu_inst_pe_1_3_5_U90 ( .A1(npu_inst_int_data_y_4__5__1_), .A2(
        npu_inst_pe_1_3_5_n54), .B1(npu_inst_pe_1_3_5_n117), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_5_n55) );
  INV_X1 npu_inst_pe_1_3_5_U89 ( .A(npu_inst_pe_1_3_5_n55), .ZN(
        npu_inst_pe_1_3_5_n102) );
  AOI22_X1 npu_inst_pe_1_3_5_U88 ( .A1(npu_inst_int_data_y_4__5__1_), .A2(
        npu_inst_pe_1_3_5_n50), .B1(npu_inst_pe_1_3_5_n116), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_5_n51) );
  INV_X1 npu_inst_pe_1_3_5_U87 ( .A(npu_inst_pe_1_3_5_n51), .ZN(
        npu_inst_pe_1_3_5_n103) );
  AOI22_X1 npu_inst_pe_1_3_5_U86 ( .A1(npu_inst_int_data_y_4__5__1_), .A2(
        npu_inst_pe_1_3_5_n46), .B1(npu_inst_pe_1_3_5_n115), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_5_n47) );
  INV_X1 npu_inst_pe_1_3_5_U85 ( .A(npu_inst_pe_1_3_5_n47), .ZN(
        npu_inst_pe_1_3_5_n104) );
  AOI22_X1 npu_inst_pe_1_3_5_U84 ( .A1(npu_inst_int_data_y_4__5__1_), .A2(
        npu_inst_pe_1_3_5_n42), .B1(npu_inst_pe_1_3_5_n114), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_5_n43) );
  INV_X1 npu_inst_pe_1_3_5_U83 ( .A(npu_inst_pe_1_3_5_n43), .ZN(
        npu_inst_pe_1_3_5_n105) );
  AOI22_X1 npu_inst_pe_1_3_5_U82 ( .A1(npu_inst_pe_1_3_5_n38), .A2(
        npu_inst_int_data_y_4__5__1_), .B1(npu_inst_pe_1_3_5_n113), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_5_n39) );
  INV_X1 npu_inst_pe_1_3_5_U81 ( .A(npu_inst_pe_1_3_5_n39), .ZN(
        npu_inst_pe_1_3_5_n106) );
  AND2_X1 npu_inst_pe_1_3_5_U80 ( .A1(npu_inst_pe_1_3_5_N93), .A2(npu_inst_n38), .ZN(npu_inst_int_data_y_3__5__0_) );
  NAND2_X1 npu_inst_pe_1_3_5_U79 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_5_n60), .ZN(npu_inst_pe_1_3_5_n74) );
  OAI21_X1 npu_inst_pe_1_3_5_U78 ( .B1(npu_inst_pe_1_3_5_n63), .B2(
        npu_inst_pe_1_3_5_n60), .A(npu_inst_pe_1_3_5_n74), .ZN(
        npu_inst_pe_1_3_5_n97) );
  NAND2_X1 npu_inst_pe_1_3_5_U77 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_5_n60), .ZN(npu_inst_pe_1_3_5_n73) );
  OAI21_X1 npu_inst_pe_1_3_5_U76 ( .B1(npu_inst_pe_1_3_5_n61), .B2(
        npu_inst_pe_1_3_5_n60), .A(npu_inst_pe_1_3_5_n73), .ZN(
        npu_inst_pe_1_3_5_n96) );
  NAND2_X1 npu_inst_pe_1_3_5_U75 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_5_n56), .ZN(npu_inst_pe_1_3_5_n72) );
  OAI21_X1 npu_inst_pe_1_3_5_U74 ( .B1(npu_inst_pe_1_3_5_n63), .B2(
        npu_inst_pe_1_3_5_n56), .A(npu_inst_pe_1_3_5_n72), .ZN(
        npu_inst_pe_1_3_5_n95) );
  NAND2_X1 npu_inst_pe_1_3_5_U73 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_5_n56), .ZN(npu_inst_pe_1_3_5_n71) );
  OAI21_X1 npu_inst_pe_1_3_5_U72 ( .B1(npu_inst_pe_1_3_5_n61), .B2(
        npu_inst_pe_1_3_5_n56), .A(npu_inst_pe_1_3_5_n71), .ZN(
        npu_inst_pe_1_3_5_n94) );
  NAND2_X1 npu_inst_pe_1_3_5_U71 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_5_n52), .ZN(npu_inst_pe_1_3_5_n70) );
  OAI21_X1 npu_inst_pe_1_3_5_U70 ( .B1(npu_inst_pe_1_3_5_n63), .B2(
        npu_inst_pe_1_3_5_n52), .A(npu_inst_pe_1_3_5_n70), .ZN(
        npu_inst_pe_1_3_5_n93) );
  NAND2_X1 npu_inst_pe_1_3_5_U69 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_5_n52), .ZN(npu_inst_pe_1_3_5_n69) );
  OAI21_X1 npu_inst_pe_1_3_5_U68 ( .B1(npu_inst_pe_1_3_5_n61), .B2(
        npu_inst_pe_1_3_5_n52), .A(npu_inst_pe_1_3_5_n69), .ZN(
        npu_inst_pe_1_3_5_n92) );
  NAND2_X1 npu_inst_pe_1_3_5_U67 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_5_n48), .ZN(npu_inst_pe_1_3_5_n68) );
  OAI21_X1 npu_inst_pe_1_3_5_U66 ( .B1(npu_inst_pe_1_3_5_n63), .B2(
        npu_inst_pe_1_3_5_n48), .A(npu_inst_pe_1_3_5_n68), .ZN(
        npu_inst_pe_1_3_5_n91) );
  NAND2_X1 npu_inst_pe_1_3_5_U65 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_5_n48), .ZN(npu_inst_pe_1_3_5_n67) );
  OAI21_X1 npu_inst_pe_1_3_5_U64 ( .B1(npu_inst_pe_1_3_5_n61), .B2(
        npu_inst_pe_1_3_5_n48), .A(npu_inst_pe_1_3_5_n67), .ZN(
        npu_inst_pe_1_3_5_n90) );
  NAND2_X1 npu_inst_pe_1_3_5_U63 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_5_n44), .ZN(npu_inst_pe_1_3_5_n66) );
  OAI21_X1 npu_inst_pe_1_3_5_U62 ( .B1(npu_inst_pe_1_3_5_n63), .B2(
        npu_inst_pe_1_3_5_n44), .A(npu_inst_pe_1_3_5_n66), .ZN(
        npu_inst_pe_1_3_5_n89) );
  NAND2_X1 npu_inst_pe_1_3_5_U61 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_5_n44), .ZN(npu_inst_pe_1_3_5_n65) );
  OAI21_X1 npu_inst_pe_1_3_5_U60 ( .B1(npu_inst_pe_1_3_5_n61), .B2(
        npu_inst_pe_1_3_5_n44), .A(npu_inst_pe_1_3_5_n65), .ZN(
        npu_inst_pe_1_3_5_n88) );
  NAND2_X1 npu_inst_pe_1_3_5_U59 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_5_n40), .ZN(npu_inst_pe_1_3_5_n64) );
  OAI21_X1 npu_inst_pe_1_3_5_U58 ( .B1(npu_inst_pe_1_3_5_n63), .B2(
        npu_inst_pe_1_3_5_n40), .A(npu_inst_pe_1_3_5_n64), .ZN(
        npu_inst_pe_1_3_5_n87) );
  NAND2_X1 npu_inst_pe_1_3_5_U57 ( .A1(npu_inst_pe_1_3_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_5_n40), .ZN(npu_inst_pe_1_3_5_n62) );
  OAI21_X1 npu_inst_pe_1_3_5_U56 ( .B1(npu_inst_pe_1_3_5_n61), .B2(
        npu_inst_pe_1_3_5_n40), .A(npu_inst_pe_1_3_5_n62), .ZN(
        npu_inst_pe_1_3_5_n86) );
  AOI22_X1 npu_inst_pe_1_3_5_U55 ( .A1(npu_inst_pe_1_3_5_n38), .A2(
        npu_inst_int_data_y_4__5__0_), .B1(npu_inst_pe_1_3_5_n113), .B2(
        npu_inst_pe_1_3_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_5_n37) );
  INV_X1 npu_inst_pe_1_3_5_U54 ( .A(npu_inst_pe_1_3_5_n37), .ZN(
        npu_inst_pe_1_3_5_n112) );
  AND2_X1 npu_inst_pe_1_3_5_U53 ( .A1(npu_inst_n38), .A2(npu_inst_pe_1_3_5_N94), .ZN(npu_inst_int_data_y_3__5__1_) );
  AOI222_X1 npu_inst_pe_1_3_5_U52 ( .A1(npu_inst_int_data_res_4__5__0_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N73), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N65), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n84) );
  INV_X1 npu_inst_pe_1_3_5_U51 ( .A(npu_inst_pe_1_3_5_n84), .ZN(
        npu_inst_pe_1_3_5_n100) );
  AOI222_X1 npu_inst_pe_1_3_5_U50 ( .A1(npu_inst_pe_1_3_5_n1), .A2(
        npu_inst_int_data_res_4__5__7_), .B1(npu_inst_pe_1_3_5_N80), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N72), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n75) );
  INV_X1 npu_inst_pe_1_3_5_U49 ( .A(npu_inst_pe_1_3_5_n75), .ZN(
        npu_inst_pe_1_3_5_n32) );
  AOI222_X1 npu_inst_pe_1_3_5_U48 ( .A1(npu_inst_int_data_res_4__5__1_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N74), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N66), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n83) );
  INV_X1 npu_inst_pe_1_3_5_U47 ( .A(npu_inst_pe_1_3_5_n83), .ZN(
        npu_inst_pe_1_3_5_n99) );
  AOI222_X1 npu_inst_pe_1_3_5_U46 ( .A1(npu_inst_int_data_res_4__5__3_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N76), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N68), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n81) );
  INV_X1 npu_inst_pe_1_3_5_U45 ( .A(npu_inst_pe_1_3_5_n81), .ZN(
        npu_inst_pe_1_3_5_n36) );
  AOI222_X1 npu_inst_pe_1_3_5_U44 ( .A1(npu_inst_int_data_res_4__5__4_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N77), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N69), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n80) );
  INV_X1 npu_inst_pe_1_3_5_U43 ( .A(npu_inst_pe_1_3_5_n80), .ZN(
        npu_inst_pe_1_3_5_n35) );
  AOI222_X1 npu_inst_pe_1_3_5_U42 ( .A1(npu_inst_int_data_res_4__5__5_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N78), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N70), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n79) );
  INV_X1 npu_inst_pe_1_3_5_U41 ( .A(npu_inst_pe_1_3_5_n79), .ZN(
        npu_inst_pe_1_3_5_n34) );
  AOI222_X1 npu_inst_pe_1_3_5_U40 ( .A1(npu_inst_int_data_res_4__5__6_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N79), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N71), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n78) );
  INV_X1 npu_inst_pe_1_3_5_U39 ( .A(npu_inst_pe_1_3_5_n78), .ZN(
        npu_inst_pe_1_3_5_n33) );
  AND2_X1 npu_inst_pe_1_3_5_U38 ( .A1(npu_inst_int_data_x_3__5__1_), .A2(
        npu_inst_pe_1_3_5_int_q_weight_1_), .ZN(npu_inst_pe_1_3_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_5_U37 ( .A1(npu_inst_int_data_x_3__5__0_), .A2(
        npu_inst_pe_1_3_5_int_q_weight_1_), .ZN(npu_inst_pe_1_3_5_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_3_5_U36 ( .A(npu_inst_pe_1_3_5_int_data_1_), .ZN(
        npu_inst_pe_1_3_5_n13) );
  NOR3_X1 npu_inst_pe_1_3_5_U35 ( .A1(npu_inst_pe_1_3_5_n26), .A2(npu_inst_n38), .A3(npu_inst_int_ckg[34]), .ZN(npu_inst_pe_1_3_5_n85) );
  OR2_X1 npu_inst_pe_1_3_5_U34 ( .A1(npu_inst_pe_1_3_5_n85), .A2(
        npu_inst_pe_1_3_5_n1), .ZN(npu_inst_pe_1_3_5_N84) );
  AOI222_X1 npu_inst_pe_1_3_5_U33 ( .A1(npu_inst_int_data_res_4__5__2_), .A2(
        npu_inst_pe_1_3_5_n1), .B1(npu_inst_pe_1_3_5_N75), .B2(
        npu_inst_pe_1_3_5_n76), .C1(npu_inst_pe_1_3_5_N67), .C2(
        npu_inst_pe_1_3_5_n77), .ZN(npu_inst_pe_1_3_5_n82) );
  INV_X1 npu_inst_pe_1_3_5_U32 ( .A(npu_inst_pe_1_3_5_n82), .ZN(
        npu_inst_pe_1_3_5_n98) );
  AOI22_X1 npu_inst_pe_1_3_5_U31 ( .A1(npu_inst_n38), .A2(
        npu_inst_int_data_y_4__5__1_), .B1(npu_inst_pe_1_3_5_n2), .B2(
        npu_inst_int_data_x_3__6__1_), .ZN(npu_inst_pe_1_3_5_n63) );
  AOI22_X1 npu_inst_pe_1_3_5_U30 ( .A1(npu_inst_n38), .A2(
        npu_inst_int_data_y_4__5__0_), .B1(npu_inst_pe_1_3_5_n2), .B2(
        npu_inst_int_data_x_3__6__0_), .ZN(npu_inst_pe_1_3_5_n61) );
  INV_X1 npu_inst_pe_1_3_5_U29 ( .A(npu_inst_pe_1_3_5_int_data_0_), .ZN(
        npu_inst_pe_1_3_5_n12) );
  INV_X1 npu_inst_pe_1_3_5_U28 ( .A(npu_inst_n51), .ZN(npu_inst_pe_1_3_5_n4)
         );
  OR3_X1 npu_inst_pe_1_3_5_U27 ( .A1(npu_inst_pe_1_3_5_n5), .A2(
        npu_inst_pe_1_3_5_n7), .A3(npu_inst_pe_1_3_5_n4), .ZN(
        npu_inst_pe_1_3_5_n56) );
  OR3_X1 npu_inst_pe_1_3_5_U26 ( .A1(npu_inst_pe_1_3_5_n4), .A2(
        npu_inst_pe_1_3_5_n7), .A3(npu_inst_pe_1_3_5_n6), .ZN(
        npu_inst_pe_1_3_5_n48) );
  INV_X1 npu_inst_pe_1_3_5_U25 ( .A(npu_inst_pe_1_3_5_n4), .ZN(
        npu_inst_pe_1_3_5_n3) );
  OR3_X1 npu_inst_pe_1_3_5_U24 ( .A1(npu_inst_pe_1_3_5_n3), .A2(
        npu_inst_pe_1_3_5_n7), .A3(npu_inst_pe_1_3_5_n6), .ZN(
        npu_inst_pe_1_3_5_n52) );
  OR3_X1 npu_inst_pe_1_3_5_U23 ( .A1(npu_inst_pe_1_3_5_n5), .A2(
        npu_inst_pe_1_3_5_n7), .A3(npu_inst_pe_1_3_5_n3), .ZN(
        npu_inst_pe_1_3_5_n60) );
  BUF_X1 npu_inst_pe_1_3_5_U22 ( .A(npu_inst_n22), .Z(npu_inst_pe_1_3_5_n1) );
  NOR2_X1 npu_inst_pe_1_3_5_U21 ( .A1(npu_inst_pe_1_3_5_n60), .A2(
        npu_inst_pe_1_3_5_n2), .ZN(npu_inst_pe_1_3_5_n58) );
  NOR2_X1 npu_inst_pe_1_3_5_U20 ( .A1(npu_inst_pe_1_3_5_n56), .A2(
        npu_inst_pe_1_3_5_n2), .ZN(npu_inst_pe_1_3_5_n54) );
  NOR2_X1 npu_inst_pe_1_3_5_U19 ( .A1(npu_inst_pe_1_3_5_n52), .A2(
        npu_inst_pe_1_3_5_n2), .ZN(npu_inst_pe_1_3_5_n50) );
  NOR2_X1 npu_inst_pe_1_3_5_U18 ( .A1(npu_inst_pe_1_3_5_n48), .A2(
        npu_inst_pe_1_3_5_n2), .ZN(npu_inst_pe_1_3_5_n46) );
  NOR2_X1 npu_inst_pe_1_3_5_U17 ( .A1(npu_inst_pe_1_3_5_n40), .A2(
        npu_inst_pe_1_3_5_n2), .ZN(npu_inst_pe_1_3_5_n38) );
  NOR2_X1 npu_inst_pe_1_3_5_U16 ( .A1(npu_inst_pe_1_3_5_n44), .A2(
        npu_inst_pe_1_3_5_n2), .ZN(npu_inst_pe_1_3_5_n42) );
  BUF_X1 npu_inst_pe_1_3_5_U15 ( .A(npu_inst_n82), .Z(npu_inst_pe_1_3_5_n7) );
  INV_X1 npu_inst_pe_1_3_5_U14 ( .A(npu_inst_n106), .ZN(npu_inst_pe_1_3_5_n11)
         );
  INV_X1 npu_inst_pe_1_3_5_U13 ( .A(npu_inst_pe_1_3_5_n38), .ZN(
        npu_inst_pe_1_3_5_n113) );
  INV_X1 npu_inst_pe_1_3_5_U12 ( .A(npu_inst_pe_1_3_5_n58), .ZN(
        npu_inst_pe_1_3_5_n118) );
  INV_X1 npu_inst_pe_1_3_5_U11 ( .A(npu_inst_pe_1_3_5_n54), .ZN(
        npu_inst_pe_1_3_5_n117) );
  INV_X1 npu_inst_pe_1_3_5_U10 ( .A(npu_inst_pe_1_3_5_n50), .ZN(
        npu_inst_pe_1_3_5_n116) );
  INV_X1 npu_inst_pe_1_3_5_U9 ( .A(npu_inst_pe_1_3_5_n46), .ZN(
        npu_inst_pe_1_3_5_n115) );
  INV_X1 npu_inst_pe_1_3_5_U8 ( .A(npu_inst_pe_1_3_5_n42), .ZN(
        npu_inst_pe_1_3_5_n114) );
  BUF_X1 npu_inst_pe_1_3_5_U7 ( .A(npu_inst_pe_1_3_5_n11), .Z(
        npu_inst_pe_1_3_5_n10) );
  BUF_X1 npu_inst_pe_1_3_5_U6 ( .A(npu_inst_pe_1_3_5_n11), .Z(
        npu_inst_pe_1_3_5_n9) );
  BUF_X1 npu_inst_pe_1_3_5_U5 ( .A(npu_inst_pe_1_3_5_n11), .Z(
        npu_inst_pe_1_3_5_n8) );
  NOR2_X1 npu_inst_pe_1_3_5_U4 ( .A1(npu_inst_pe_1_3_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_5_n1), .ZN(npu_inst_pe_1_3_5_n76) );
  NOR2_X1 npu_inst_pe_1_3_5_U3 ( .A1(npu_inst_pe_1_3_5_n27), .A2(
        npu_inst_pe_1_3_5_n1), .ZN(npu_inst_pe_1_3_5_n77) );
  FA_X1 npu_inst_pe_1_3_5_sub_77_U2_1 ( .A(npu_inst_int_data_res_3__5__1_), 
        .B(npu_inst_pe_1_3_5_n13), .CI(npu_inst_pe_1_3_5_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_3_5_sub_77_carry_2_), .S(npu_inst_pe_1_3_5_N66) );
  FA_X1 npu_inst_pe_1_3_5_add_79_U1_1 ( .A(npu_inst_int_data_res_3__5__1_), 
        .B(npu_inst_pe_1_3_5_int_data_1_), .CI(
        npu_inst_pe_1_3_5_add_79_carry_1_), .CO(
        npu_inst_pe_1_3_5_add_79_carry_2_), .S(npu_inst_pe_1_3_5_N74) );
  NAND3_X1 npu_inst_pe_1_3_5_U101 ( .A1(npu_inst_pe_1_3_5_n4), .A2(
        npu_inst_pe_1_3_5_n6), .A3(npu_inst_pe_1_3_5_n7), .ZN(
        npu_inst_pe_1_3_5_n44) );
  NAND3_X1 npu_inst_pe_1_3_5_U100 ( .A1(npu_inst_pe_1_3_5_n3), .A2(
        npu_inst_pe_1_3_5_n6), .A3(npu_inst_pe_1_3_5_n7), .ZN(
        npu_inst_pe_1_3_5_n40) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_5_n33), .CK(
        npu_inst_pe_1_3_5_net3811), .RN(npu_inst_pe_1_3_5_n8), .Q(
        npu_inst_int_data_res_3__5__6_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_5_n34), .CK(
        npu_inst_pe_1_3_5_net3811), .RN(npu_inst_pe_1_3_5_n8), .Q(
        npu_inst_int_data_res_3__5__5_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_5_n35), .CK(
        npu_inst_pe_1_3_5_net3811), .RN(npu_inst_pe_1_3_5_n8), .Q(
        npu_inst_int_data_res_3__5__4_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_5_n36), .CK(
        npu_inst_pe_1_3_5_net3811), .RN(npu_inst_pe_1_3_5_n8), .Q(
        npu_inst_int_data_res_3__5__3_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_5_n98), .CK(
        npu_inst_pe_1_3_5_net3811), .RN(npu_inst_pe_1_3_5_n8), .Q(
        npu_inst_int_data_res_3__5__2_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_5_n99), .CK(
        npu_inst_pe_1_3_5_net3811), .RN(npu_inst_pe_1_3_5_n8), .Q(
        npu_inst_int_data_res_3__5__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_5_n32), .CK(
        npu_inst_pe_1_3_5_net3811), .RN(npu_inst_pe_1_3_5_n8), .Q(
        npu_inst_int_data_res_3__5__7_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_5_n100), 
        .CK(npu_inst_pe_1_3_5_net3811), .RN(npu_inst_pe_1_3_5_n8), .Q(
        npu_inst_int_data_res_3__5__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_weight_reg_0_ ( .D(npu_inst_n92), .CK(
        npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n8), .Q(
        npu_inst_pe_1_3_5_int_q_weight_0_), .QN(npu_inst_pe_1_3_5_n27) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_weight_reg_1_ ( .D(npu_inst_n98), .CK(
        npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n8), .Q(
        npu_inst_pe_1_3_5_int_q_weight_1_), .QN(npu_inst_pe_1_3_5_n26) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_5_n112), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n8), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_5_n106), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n8), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_5_n111), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_5_n105), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_5_n110), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_5_n104), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_5_n109), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_5_n103), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_5_n108), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_5_n102), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_5_n107), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_5_n101), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_5_n86), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_5_n87), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n9), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_5_n88), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_5_n89), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_5_n90), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_5_n91), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_5_n92), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_5_n93), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_5_n94), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_5_n95), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_5_n96), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_5_n97), 
        .CK(npu_inst_pe_1_3_5_net3817), .RN(npu_inst_pe_1_3_5_n10), .Q(
        npu_inst_pe_1_3_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_5_net3811) );
  CLKGATETST_X1 npu_inst_pe_1_3_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n46), .SE(1'b0), .GCK(npu_inst_pe_1_3_5_net3817) );
  MUX2_X1 npu_inst_pe_1_3_6_U153 ( .A(npu_inst_pe_1_3_6_n31), .B(
        npu_inst_pe_1_3_6_n28), .S(npu_inst_pe_1_3_6_n7), .Z(
        npu_inst_pe_1_3_6_N93) );
  MUX2_X1 npu_inst_pe_1_3_6_U152 ( .A(npu_inst_pe_1_3_6_n30), .B(
        npu_inst_pe_1_3_6_n29), .S(npu_inst_pe_1_3_6_n5), .Z(
        npu_inst_pe_1_3_6_n31) );
  MUX2_X1 npu_inst_pe_1_3_6_U151 ( .A(npu_inst_pe_1_3_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_6_n3), .Z(
        npu_inst_pe_1_3_6_n30) );
  MUX2_X1 npu_inst_pe_1_3_6_U150 ( .A(npu_inst_pe_1_3_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_6_n3), .Z(
        npu_inst_pe_1_3_6_n29) );
  MUX2_X1 npu_inst_pe_1_3_6_U149 ( .A(npu_inst_pe_1_3_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_6_n3), .Z(
        npu_inst_pe_1_3_6_n28) );
  MUX2_X1 npu_inst_pe_1_3_6_U148 ( .A(npu_inst_pe_1_3_6_n25), .B(
        npu_inst_pe_1_3_6_n22), .S(npu_inst_pe_1_3_6_n7), .Z(
        npu_inst_pe_1_3_6_N94) );
  MUX2_X1 npu_inst_pe_1_3_6_U147 ( .A(npu_inst_pe_1_3_6_n24), .B(
        npu_inst_pe_1_3_6_n23), .S(npu_inst_pe_1_3_6_n5), .Z(
        npu_inst_pe_1_3_6_n25) );
  MUX2_X1 npu_inst_pe_1_3_6_U146 ( .A(npu_inst_pe_1_3_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_6_n3), .Z(
        npu_inst_pe_1_3_6_n24) );
  MUX2_X1 npu_inst_pe_1_3_6_U145 ( .A(npu_inst_pe_1_3_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_6_n3), .Z(
        npu_inst_pe_1_3_6_n23) );
  MUX2_X1 npu_inst_pe_1_3_6_U144 ( .A(npu_inst_pe_1_3_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_6_n3), .Z(
        npu_inst_pe_1_3_6_n22) );
  MUX2_X1 npu_inst_pe_1_3_6_U143 ( .A(npu_inst_pe_1_3_6_n21), .B(
        npu_inst_pe_1_3_6_n18), .S(npu_inst_pe_1_3_6_n7), .Z(
        npu_inst_int_data_x_3__6__1_) );
  MUX2_X1 npu_inst_pe_1_3_6_U142 ( .A(npu_inst_pe_1_3_6_n20), .B(
        npu_inst_pe_1_3_6_n19), .S(npu_inst_pe_1_3_6_n5), .Z(
        npu_inst_pe_1_3_6_n21) );
  MUX2_X1 npu_inst_pe_1_3_6_U141 ( .A(npu_inst_pe_1_3_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_6_n3), .Z(
        npu_inst_pe_1_3_6_n20) );
  MUX2_X1 npu_inst_pe_1_3_6_U140 ( .A(npu_inst_pe_1_3_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_6_n3), .Z(
        npu_inst_pe_1_3_6_n19) );
  MUX2_X1 npu_inst_pe_1_3_6_U139 ( .A(npu_inst_pe_1_3_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_6_n3), .Z(
        npu_inst_pe_1_3_6_n18) );
  MUX2_X1 npu_inst_pe_1_3_6_U138 ( .A(npu_inst_pe_1_3_6_n17), .B(
        npu_inst_pe_1_3_6_n14), .S(npu_inst_pe_1_3_6_n7), .Z(
        npu_inst_int_data_x_3__6__0_) );
  MUX2_X1 npu_inst_pe_1_3_6_U137 ( .A(npu_inst_pe_1_3_6_n16), .B(
        npu_inst_pe_1_3_6_n15), .S(npu_inst_pe_1_3_6_n5), .Z(
        npu_inst_pe_1_3_6_n17) );
  MUX2_X1 npu_inst_pe_1_3_6_U136 ( .A(npu_inst_pe_1_3_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_6_n3), .Z(
        npu_inst_pe_1_3_6_n16) );
  MUX2_X1 npu_inst_pe_1_3_6_U135 ( .A(npu_inst_pe_1_3_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_6_n3), .Z(
        npu_inst_pe_1_3_6_n15) );
  MUX2_X1 npu_inst_pe_1_3_6_U134 ( .A(npu_inst_pe_1_3_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_6_n3), .Z(
        npu_inst_pe_1_3_6_n14) );
  XOR2_X1 npu_inst_pe_1_3_6_U133 ( .A(npu_inst_pe_1_3_6_int_data_0_), .B(
        npu_inst_int_data_res_3__6__0_), .Z(npu_inst_pe_1_3_6_N73) );
  AND2_X1 npu_inst_pe_1_3_6_U132 ( .A1(npu_inst_int_data_res_3__6__0_), .A2(
        npu_inst_pe_1_3_6_int_data_0_), .ZN(npu_inst_pe_1_3_6_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_6_U131 ( .A(npu_inst_int_data_res_3__6__0_), .B(
        npu_inst_pe_1_3_6_n12), .ZN(npu_inst_pe_1_3_6_N65) );
  OR2_X1 npu_inst_pe_1_3_6_U130 ( .A1(npu_inst_pe_1_3_6_n12), .A2(
        npu_inst_int_data_res_3__6__0_), .ZN(npu_inst_pe_1_3_6_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_6_U129 ( .A(npu_inst_int_data_res_3__6__2_), .B(
        npu_inst_pe_1_3_6_add_79_carry_2_), .Z(npu_inst_pe_1_3_6_N75) );
  AND2_X1 npu_inst_pe_1_3_6_U128 ( .A1(npu_inst_pe_1_3_6_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_3__6__2_), .ZN(
        npu_inst_pe_1_3_6_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_6_U127 ( .A(npu_inst_int_data_res_3__6__3_), .B(
        npu_inst_pe_1_3_6_add_79_carry_3_), .Z(npu_inst_pe_1_3_6_N76) );
  AND2_X1 npu_inst_pe_1_3_6_U126 ( .A1(npu_inst_pe_1_3_6_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_3__6__3_), .ZN(
        npu_inst_pe_1_3_6_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_6_U125 ( .A(npu_inst_int_data_res_3__6__4_), .B(
        npu_inst_pe_1_3_6_add_79_carry_4_), .Z(npu_inst_pe_1_3_6_N77) );
  AND2_X1 npu_inst_pe_1_3_6_U124 ( .A1(npu_inst_pe_1_3_6_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_3__6__4_), .ZN(
        npu_inst_pe_1_3_6_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_6_U123 ( .A(npu_inst_int_data_res_3__6__5_), .B(
        npu_inst_pe_1_3_6_add_79_carry_5_), .Z(npu_inst_pe_1_3_6_N78) );
  AND2_X1 npu_inst_pe_1_3_6_U122 ( .A1(npu_inst_pe_1_3_6_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_3__6__5_), .ZN(
        npu_inst_pe_1_3_6_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_6_U121 ( .A(npu_inst_int_data_res_3__6__6_), .B(
        npu_inst_pe_1_3_6_add_79_carry_6_), .Z(npu_inst_pe_1_3_6_N79) );
  AND2_X1 npu_inst_pe_1_3_6_U120 ( .A1(npu_inst_pe_1_3_6_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_3__6__6_), .ZN(
        npu_inst_pe_1_3_6_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_6_U119 ( .A(npu_inst_int_data_res_3__6__7_), .B(
        npu_inst_pe_1_3_6_add_79_carry_7_), .Z(npu_inst_pe_1_3_6_N80) );
  XNOR2_X1 npu_inst_pe_1_3_6_U118 ( .A(npu_inst_pe_1_3_6_sub_77_carry_2_), .B(
        npu_inst_int_data_res_3__6__2_), .ZN(npu_inst_pe_1_3_6_N67) );
  OR2_X1 npu_inst_pe_1_3_6_U117 ( .A1(npu_inst_int_data_res_3__6__2_), .A2(
        npu_inst_pe_1_3_6_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_3_6_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_6_U116 ( .A(npu_inst_pe_1_3_6_sub_77_carry_3_), .B(
        npu_inst_int_data_res_3__6__3_), .ZN(npu_inst_pe_1_3_6_N68) );
  OR2_X1 npu_inst_pe_1_3_6_U115 ( .A1(npu_inst_int_data_res_3__6__3_), .A2(
        npu_inst_pe_1_3_6_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_3_6_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_6_U114 ( .A(npu_inst_pe_1_3_6_sub_77_carry_4_), .B(
        npu_inst_int_data_res_3__6__4_), .ZN(npu_inst_pe_1_3_6_N69) );
  OR2_X1 npu_inst_pe_1_3_6_U113 ( .A1(npu_inst_int_data_res_3__6__4_), .A2(
        npu_inst_pe_1_3_6_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_3_6_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_6_U112 ( .A(npu_inst_pe_1_3_6_sub_77_carry_5_), .B(
        npu_inst_int_data_res_3__6__5_), .ZN(npu_inst_pe_1_3_6_N70) );
  OR2_X1 npu_inst_pe_1_3_6_U111 ( .A1(npu_inst_int_data_res_3__6__5_), .A2(
        npu_inst_pe_1_3_6_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_3_6_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_6_U110 ( .A(npu_inst_pe_1_3_6_sub_77_carry_6_), .B(
        npu_inst_int_data_res_3__6__6_), .ZN(npu_inst_pe_1_3_6_N71) );
  OR2_X1 npu_inst_pe_1_3_6_U109 ( .A1(npu_inst_int_data_res_3__6__6_), .A2(
        npu_inst_pe_1_3_6_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_3_6_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_6_U108 ( .A(npu_inst_int_data_res_3__6__7_), .B(
        npu_inst_pe_1_3_6_sub_77_carry_7_), .ZN(npu_inst_pe_1_3_6_N72) );
  INV_X1 npu_inst_pe_1_3_6_U107 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_3_6_n6)
         );
  INV_X1 npu_inst_pe_1_3_6_U106 ( .A(npu_inst_pe_1_3_6_n6), .ZN(
        npu_inst_pe_1_3_6_n5) );
  INV_X1 npu_inst_pe_1_3_6_U105 ( .A(npu_inst_n38), .ZN(npu_inst_pe_1_3_6_n2)
         );
  AOI22_X1 npu_inst_pe_1_3_6_U104 ( .A1(npu_inst_int_data_y_4__6__0_), .A2(
        npu_inst_pe_1_3_6_n58), .B1(npu_inst_pe_1_3_6_n118), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_6_n57) );
  INV_X1 npu_inst_pe_1_3_6_U103 ( .A(npu_inst_pe_1_3_6_n57), .ZN(
        npu_inst_pe_1_3_6_n107) );
  AOI22_X1 npu_inst_pe_1_3_6_U102 ( .A1(npu_inst_int_data_y_4__6__0_), .A2(
        npu_inst_pe_1_3_6_n54), .B1(npu_inst_pe_1_3_6_n117), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_6_n53) );
  INV_X1 npu_inst_pe_1_3_6_U99 ( .A(npu_inst_pe_1_3_6_n53), .ZN(
        npu_inst_pe_1_3_6_n108) );
  AOI22_X1 npu_inst_pe_1_3_6_U98 ( .A1(npu_inst_int_data_y_4__6__0_), .A2(
        npu_inst_pe_1_3_6_n50), .B1(npu_inst_pe_1_3_6_n116), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_6_n49) );
  INV_X1 npu_inst_pe_1_3_6_U97 ( .A(npu_inst_pe_1_3_6_n49), .ZN(
        npu_inst_pe_1_3_6_n109) );
  AOI22_X1 npu_inst_pe_1_3_6_U96 ( .A1(npu_inst_int_data_y_4__6__0_), .A2(
        npu_inst_pe_1_3_6_n46), .B1(npu_inst_pe_1_3_6_n115), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_6_n45) );
  INV_X1 npu_inst_pe_1_3_6_U95 ( .A(npu_inst_pe_1_3_6_n45), .ZN(
        npu_inst_pe_1_3_6_n110) );
  AOI22_X1 npu_inst_pe_1_3_6_U94 ( .A1(npu_inst_int_data_y_4__6__0_), .A2(
        npu_inst_pe_1_3_6_n42), .B1(npu_inst_pe_1_3_6_n114), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_6_n41) );
  INV_X1 npu_inst_pe_1_3_6_U93 ( .A(npu_inst_pe_1_3_6_n41), .ZN(
        npu_inst_pe_1_3_6_n111) );
  AOI22_X1 npu_inst_pe_1_3_6_U92 ( .A1(npu_inst_int_data_y_4__6__1_), .A2(
        npu_inst_pe_1_3_6_n58), .B1(npu_inst_pe_1_3_6_n118), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_6_n59) );
  INV_X1 npu_inst_pe_1_3_6_U91 ( .A(npu_inst_pe_1_3_6_n59), .ZN(
        npu_inst_pe_1_3_6_n101) );
  AOI22_X1 npu_inst_pe_1_3_6_U90 ( .A1(npu_inst_int_data_y_4__6__1_), .A2(
        npu_inst_pe_1_3_6_n54), .B1(npu_inst_pe_1_3_6_n117), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_6_n55) );
  INV_X1 npu_inst_pe_1_3_6_U89 ( .A(npu_inst_pe_1_3_6_n55), .ZN(
        npu_inst_pe_1_3_6_n102) );
  AOI22_X1 npu_inst_pe_1_3_6_U88 ( .A1(npu_inst_int_data_y_4__6__1_), .A2(
        npu_inst_pe_1_3_6_n50), .B1(npu_inst_pe_1_3_6_n116), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_6_n51) );
  INV_X1 npu_inst_pe_1_3_6_U87 ( .A(npu_inst_pe_1_3_6_n51), .ZN(
        npu_inst_pe_1_3_6_n103) );
  AOI22_X1 npu_inst_pe_1_3_6_U86 ( .A1(npu_inst_int_data_y_4__6__1_), .A2(
        npu_inst_pe_1_3_6_n46), .B1(npu_inst_pe_1_3_6_n115), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_6_n47) );
  INV_X1 npu_inst_pe_1_3_6_U85 ( .A(npu_inst_pe_1_3_6_n47), .ZN(
        npu_inst_pe_1_3_6_n104) );
  AOI22_X1 npu_inst_pe_1_3_6_U84 ( .A1(npu_inst_int_data_y_4__6__1_), .A2(
        npu_inst_pe_1_3_6_n42), .B1(npu_inst_pe_1_3_6_n114), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_6_n43) );
  INV_X1 npu_inst_pe_1_3_6_U83 ( .A(npu_inst_pe_1_3_6_n43), .ZN(
        npu_inst_pe_1_3_6_n105) );
  AOI22_X1 npu_inst_pe_1_3_6_U82 ( .A1(npu_inst_pe_1_3_6_n38), .A2(
        npu_inst_int_data_y_4__6__1_), .B1(npu_inst_pe_1_3_6_n113), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_6_n39) );
  INV_X1 npu_inst_pe_1_3_6_U81 ( .A(npu_inst_pe_1_3_6_n39), .ZN(
        npu_inst_pe_1_3_6_n106) );
  AND2_X1 npu_inst_pe_1_3_6_U80 ( .A1(npu_inst_pe_1_3_6_N93), .A2(npu_inst_n38), .ZN(npu_inst_int_data_y_3__6__0_) );
  NAND2_X1 npu_inst_pe_1_3_6_U79 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_6_n60), .ZN(npu_inst_pe_1_3_6_n74) );
  OAI21_X1 npu_inst_pe_1_3_6_U78 ( .B1(npu_inst_pe_1_3_6_n63), .B2(
        npu_inst_pe_1_3_6_n60), .A(npu_inst_pe_1_3_6_n74), .ZN(
        npu_inst_pe_1_3_6_n97) );
  NAND2_X1 npu_inst_pe_1_3_6_U77 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_6_n60), .ZN(npu_inst_pe_1_3_6_n73) );
  OAI21_X1 npu_inst_pe_1_3_6_U76 ( .B1(npu_inst_pe_1_3_6_n61), .B2(
        npu_inst_pe_1_3_6_n60), .A(npu_inst_pe_1_3_6_n73), .ZN(
        npu_inst_pe_1_3_6_n96) );
  NAND2_X1 npu_inst_pe_1_3_6_U75 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_6_n56), .ZN(npu_inst_pe_1_3_6_n72) );
  OAI21_X1 npu_inst_pe_1_3_6_U74 ( .B1(npu_inst_pe_1_3_6_n63), .B2(
        npu_inst_pe_1_3_6_n56), .A(npu_inst_pe_1_3_6_n72), .ZN(
        npu_inst_pe_1_3_6_n95) );
  NAND2_X1 npu_inst_pe_1_3_6_U73 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_6_n56), .ZN(npu_inst_pe_1_3_6_n71) );
  OAI21_X1 npu_inst_pe_1_3_6_U72 ( .B1(npu_inst_pe_1_3_6_n61), .B2(
        npu_inst_pe_1_3_6_n56), .A(npu_inst_pe_1_3_6_n71), .ZN(
        npu_inst_pe_1_3_6_n94) );
  NAND2_X1 npu_inst_pe_1_3_6_U71 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_6_n52), .ZN(npu_inst_pe_1_3_6_n70) );
  OAI21_X1 npu_inst_pe_1_3_6_U70 ( .B1(npu_inst_pe_1_3_6_n63), .B2(
        npu_inst_pe_1_3_6_n52), .A(npu_inst_pe_1_3_6_n70), .ZN(
        npu_inst_pe_1_3_6_n93) );
  NAND2_X1 npu_inst_pe_1_3_6_U69 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_6_n52), .ZN(npu_inst_pe_1_3_6_n69) );
  OAI21_X1 npu_inst_pe_1_3_6_U68 ( .B1(npu_inst_pe_1_3_6_n61), .B2(
        npu_inst_pe_1_3_6_n52), .A(npu_inst_pe_1_3_6_n69), .ZN(
        npu_inst_pe_1_3_6_n92) );
  NAND2_X1 npu_inst_pe_1_3_6_U67 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_6_n48), .ZN(npu_inst_pe_1_3_6_n68) );
  OAI21_X1 npu_inst_pe_1_3_6_U66 ( .B1(npu_inst_pe_1_3_6_n63), .B2(
        npu_inst_pe_1_3_6_n48), .A(npu_inst_pe_1_3_6_n68), .ZN(
        npu_inst_pe_1_3_6_n91) );
  NAND2_X1 npu_inst_pe_1_3_6_U65 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_6_n48), .ZN(npu_inst_pe_1_3_6_n67) );
  OAI21_X1 npu_inst_pe_1_3_6_U64 ( .B1(npu_inst_pe_1_3_6_n61), .B2(
        npu_inst_pe_1_3_6_n48), .A(npu_inst_pe_1_3_6_n67), .ZN(
        npu_inst_pe_1_3_6_n90) );
  NAND2_X1 npu_inst_pe_1_3_6_U63 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_6_n44), .ZN(npu_inst_pe_1_3_6_n66) );
  OAI21_X1 npu_inst_pe_1_3_6_U62 ( .B1(npu_inst_pe_1_3_6_n63), .B2(
        npu_inst_pe_1_3_6_n44), .A(npu_inst_pe_1_3_6_n66), .ZN(
        npu_inst_pe_1_3_6_n89) );
  NAND2_X1 npu_inst_pe_1_3_6_U61 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_6_n44), .ZN(npu_inst_pe_1_3_6_n65) );
  OAI21_X1 npu_inst_pe_1_3_6_U60 ( .B1(npu_inst_pe_1_3_6_n61), .B2(
        npu_inst_pe_1_3_6_n44), .A(npu_inst_pe_1_3_6_n65), .ZN(
        npu_inst_pe_1_3_6_n88) );
  NAND2_X1 npu_inst_pe_1_3_6_U59 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_6_n40), .ZN(npu_inst_pe_1_3_6_n64) );
  OAI21_X1 npu_inst_pe_1_3_6_U58 ( .B1(npu_inst_pe_1_3_6_n63), .B2(
        npu_inst_pe_1_3_6_n40), .A(npu_inst_pe_1_3_6_n64), .ZN(
        npu_inst_pe_1_3_6_n87) );
  NAND2_X1 npu_inst_pe_1_3_6_U57 ( .A1(npu_inst_pe_1_3_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_6_n40), .ZN(npu_inst_pe_1_3_6_n62) );
  OAI21_X1 npu_inst_pe_1_3_6_U56 ( .B1(npu_inst_pe_1_3_6_n61), .B2(
        npu_inst_pe_1_3_6_n40), .A(npu_inst_pe_1_3_6_n62), .ZN(
        npu_inst_pe_1_3_6_n86) );
  AOI22_X1 npu_inst_pe_1_3_6_U55 ( .A1(npu_inst_pe_1_3_6_n38), .A2(
        npu_inst_int_data_y_4__6__0_), .B1(npu_inst_pe_1_3_6_n113), .B2(
        npu_inst_pe_1_3_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_6_n37) );
  INV_X1 npu_inst_pe_1_3_6_U54 ( .A(npu_inst_pe_1_3_6_n37), .ZN(
        npu_inst_pe_1_3_6_n112) );
  AND2_X1 npu_inst_pe_1_3_6_U53 ( .A1(npu_inst_n38), .A2(npu_inst_pe_1_3_6_N94), .ZN(npu_inst_int_data_y_3__6__1_) );
  AOI222_X1 npu_inst_pe_1_3_6_U52 ( .A1(npu_inst_int_data_res_4__6__0_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N73), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N65), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n84) );
  INV_X1 npu_inst_pe_1_3_6_U51 ( .A(npu_inst_pe_1_3_6_n84), .ZN(
        npu_inst_pe_1_3_6_n100) );
  AOI222_X1 npu_inst_pe_1_3_6_U50 ( .A1(npu_inst_pe_1_3_6_n1), .A2(
        npu_inst_int_data_res_4__6__7_), .B1(npu_inst_pe_1_3_6_N80), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N72), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n75) );
  INV_X1 npu_inst_pe_1_3_6_U49 ( .A(npu_inst_pe_1_3_6_n75), .ZN(
        npu_inst_pe_1_3_6_n32) );
  AOI222_X1 npu_inst_pe_1_3_6_U48 ( .A1(npu_inst_int_data_res_4__6__1_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N74), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N66), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n83) );
  INV_X1 npu_inst_pe_1_3_6_U47 ( .A(npu_inst_pe_1_3_6_n83), .ZN(
        npu_inst_pe_1_3_6_n99) );
  AOI222_X1 npu_inst_pe_1_3_6_U46 ( .A1(npu_inst_int_data_res_4__6__3_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N76), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N68), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n81) );
  INV_X1 npu_inst_pe_1_3_6_U45 ( .A(npu_inst_pe_1_3_6_n81), .ZN(
        npu_inst_pe_1_3_6_n36) );
  AOI222_X1 npu_inst_pe_1_3_6_U44 ( .A1(npu_inst_int_data_res_4__6__4_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N77), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N69), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n80) );
  INV_X1 npu_inst_pe_1_3_6_U43 ( .A(npu_inst_pe_1_3_6_n80), .ZN(
        npu_inst_pe_1_3_6_n35) );
  AOI222_X1 npu_inst_pe_1_3_6_U42 ( .A1(npu_inst_int_data_res_4__6__5_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N78), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N70), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n79) );
  INV_X1 npu_inst_pe_1_3_6_U41 ( .A(npu_inst_pe_1_3_6_n79), .ZN(
        npu_inst_pe_1_3_6_n34) );
  AOI222_X1 npu_inst_pe_1_3_6_U40 ( .A1(npu_inst_int_data_res_4__6__6_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N79), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N71), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n78) );
  INV_X1 npu_inst_pe_1_3_6_U39 ( .A(npu_inst_pe_1_3_6_n78), .ZN(
        npu_inst_pe_1_3_6_n33) );
  AND2_X1 npu_inst_pe_1_3_6_U38 ( .A1(npu_inst_int_data_x_3__6__1_), .A2(
        npu_inst_pe_1_3_6_int_q_weight_1_), .ZN(npu_inst_pe_1_3_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_6_U37 ( .A1(npu_inst_int_data_x_3__6__0_), .A2(
        npu_inst_pe_1_3_6_int_q_weight_1_), .ZN(npu_inst_pe_1_3_6_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_3_6_U36 ( .A(npu_inst_pe_1_3_6_int_data_1_), .ZN(
        npu_inst_pe_1_3_6_n13) );
  NOR3_X1 npu_inst_pe_1_3_6_U35 ( .A1(npu_inst_pe_1_3_6_n26), .A2(npu_inst_n38), .A3(npu_inst_int_ckg[33]), .ZN(npu_inst_pe_1_3_6_n85) );
  OR2_X1 npu_inst_pe_1_3_6_U34 ( .A1(npu_inst_pe_1_3_6_n85), .A2(
        npu_inst_pe_1_3_6_n1), .ZN(npu_inst_pe_1_3_6_N84) );
  AOI222_X1 npu_inst_pe_1_3_6_U33 ( .A1(npu_inst_int_data_res_4__6__2_), .A2(
        npu_inst_pe_1_3_6_n1), .B1(npu_inst_pe_1_3_6_N75), .B2(
        npu_inst_pe_1_3_6_n76), .C1(npu_inst_pe_1_3_6_N67), .C2(
        npu_inst_pe_1_3_6_n77), .ZN(npu_inst_pe_1_3_6_n82) );
  INV_X1 npu_inst_pe_1_3_6_U32 ( .A(npu_inst_pe_1_3_6_n82), .ZN(
        npu_inst_pe_1_3_6_n98) );
  AOI22_X1 npu_inst_pe_1_3_6_U31 ( .A1(npu_inst_n38), .A2(
        npu_inst_int_data_y_4__6__1_), .B1(npu_inst_pe_1_3_6_n2), .B2(
        npu_inst_int_data_x_3__7__1_), .ZN(npu_inst_pe_1_3_6_n63) );
  AOI22_X1 npu_inst_pe_1_3_6_U30 ( .A1(npu_inst_n38), .A2(
        npu_inst_int_data_y_4__6__0_), .B1(npu_inst_pe_1_3_6_n2), .B2(
        npu_inst_int_data_x_3__7__0_), .ZN(npu_inst_pe_1_3_6_n61) );
  INV_X1 npu_inst_pe_1_3_6_U29 ( .A(npu_inst_pe_1_3_6_int_data_0_), .ZN(
        npu_inst_pe_1_3_6_n12) );
  INV_X1 npu_inst_pe_1_3_6_U28 ( .A(npu_inst_n51), .ZN(npu_inst_pe_1_3_6_n4)
         );
  OR3_X1 npu_inst_pe_1_3_6_U27 ( .A1(npu_inst_pe_1_3_6_n5), .A2(
        npu_inst_pe_1_3_6_n7), .A3(npu_inst_pe_1_3_6_n4), .ZN(
        npu_inst_pe_1_3_6_n56) );
  OR3_X1 npu_inst_pe_1_3_6_U26 ( .A1(npu_inst_pe_1_3_6_n4), .A2(
        npu_inst_pe_1_3_6_n7), .A3(npu_inst_pe_1_3_6_n6), .ZN(
        npu_inst_pe_1_3_6_n48) );
  INV_X1 npu_inst_pe_1_3_6_U25 ( .A(npu_inst_pe_1_3_6_n4), .ZN(
        npu_inst_pe_1_3_6_n3) );
  OR3_X1 npu_inst_pe_1_3_6_U24 ( .A1(npu_inst_pe_1_3_6_n3), .A2(
        npu_inst_pe_1_3_6_n7), .A3(npu_inst_pe_1_3_6_n6), .ZN(
        npu_inst_pe_1_3_6_n52) );
  OR3_X1 npu_inst_pe_1_3_6_U23 ( .A1(npu_inst_pe_1_3_6_n5), .A2(
        npu_inst_pe_1_3_6_n7), .A3(npu_inst_pe_1_3_6_n3), .ZN(
        npu_inst_pe_1_3_6_n60) );
  BUF_X1 npu_inst_pe_1_3_6_U22 ( .A(npu_inst_n22), .Z(npu_inst_pe_1_3_6_n1) );
  NOR2_X1 npu_inst_pe_1_3_6_U21 ( .A1(npu_inst_pe_1_3_6_n60), .A2(
        npu_inst_pe_1_3_6_n2), .ZN(npu_inst_pe_1_3_6_n58) );
  NOR2_X1 npu_inst_pe_1_3_6_U20 ( .A1(npu_inst_pe_1_3_6_n56), .A2(
        npu_inst_pe_1_3_6_n2), .ZN(npu_inst_pe_1_3_6_n54) );
  NOR2_X1 npu_inst_pe_1_3_6_U19 ( .A1(npu_inst_pe_1_3_6_n52), .A2(
        npu_inst_pe_1_3_6_n2), .ZN(npu_inst_pe_1_3_6_n50) );
  NOR2_X1 npu_inst_pe_1_3_6_U18 ( .A1(npu_inst_pe_1_3_6_n48), .A2(
        npu_inst_pe_1_3_6_n2), .ZN(npu_inst_pe_1_3_6_n46) );
  NOR2_X1 npu_inst_pe_1_3_6_U17 ( .A1(npu_inst_pe_1_3_6_n40), .A2(
        npu_inst_pe_1_3_6_n2), .ZN(npu_inst_pe_1_3_6_n38) );
  NOR2_X1 npu_inst_pe_1_3_6_U16 ( .A1(npu_inst_pe_1_3_6_n44), .A2(
        npu_inst_pe_1_3_6_n2), .ZN(npu_inst_pe_1_3_6_n42) );
  BUF_X1 npu_inst_pe_1_3_6_U15 ( .A(npu_inst_n82), .Z(npu_inst_pe_1_3_6_n7) );
  INV_X1 npu_inst_pe_1_3_6_U14 ( .A(npu_inst_n106), .ZN(npu_inst_pe_1_3_6_n11)
         );
  INV_X1 npu_inst_pe_1_3_6_U13 ( .A(npu_inst_pe_1_3_6_n38), .ZN(
        npu_inst_pe_1_3_6_n113) );
  INV_X1 npu_inst_pe_1_3_6_U12 ( .A(npu_inst_pe_1_3_6_n58), .ZN(
        npu_inst_pe_1_3_6_n118) );
  INV_X1 npu_inst_pe_1_3_6_U11 ( .A(npu_inst_pe_1_3_6_n54), .ZN(
        npu_inst_pe_1_3_6_n117) );
  INV_X1 npu_inst_pe_1_3_6_U10 ( .A(npu_inst_pe_1_3_6_n50), .ZN(
        npu_inst_pe_1_3_6_n116) );
  INV_X1 npu_inst_pe_1_3_6_U9 ( .A(npu_inst_pe_1_3_6_n46), .ZN(
        npu_inst_pe_1_3_6_n115) );
  INV_X1 npu_inst_pe_1_3_6_U8 ( .A(npu_inst_pe_1_3_6_n42), .ZN(
        npu_inst_pe_1_3_6_n114) );
  BUF_X1 npu_inst_pe_1_3_6_U7 ( .A(npu_inst_pe_1_3_6_n11), .Z(
        npu_inst_pe_1_3_6_n10) );
  BUF_X1 npu_inst_pe_1_3_6_U6 ( .A(npu_inst_pe_1_3_6_n11), .Z(
        npu_inst_pe_1_3_6_n9) );
  BUF_X1 npu_inst_pe_1_3_6_U5 ( .A(npu_inst_pe_1_3_6_n11), .Z(
        npu_inst_pe_1_3_6_n8) );
  NOR2_X1 npu_inst_pe_1_3_6_U4 ( .A1(npu_inst_pe_1_3_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_6_n1), .ZN(npu_inst_pe_1_3_6_n76) );
  NOR2_X1 npu_inst_pe_1_3_6_U3 ( .A1(npu_inst_pe_1_3_6_n27), .A2(
        npu_inst_pe_1_3_6_n1), .ZN(npu_inst_pe_1_3_6_n77) );
  FA_X1 npu_inst_pe_1_3_6_sub_77_U2_1 ( .A(npu_inst_int_data_res_3__6__1_), 
        .B(npu_inst_pe_1_3_6_n13), .CI(npu_inst_pe_1_3_6_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_3_6_sub_77_carry_2_), .S(npu_inst_pe_1_3_6_N66) );
  FA_X1 npu_inst_pe_1_3_6_add_79_U1_1 ( .A(npu_inst_int_data_res_3__6__1_), 
        .B(npu_inst_pe_1_3_6_int_data_1_), .CI(
        npu_inst_pe_1_3_6_add_79_carry_1_), .CO(
        npu_inst_pe_1_3_6_add_79_carry_2_), .S(npu_inst_pe_1_3_6_N74) );
  NAND3_X1 npu_inst_pe_1_3_6_U101 ( .A1(npu_inst_pe_1_3_6_n4), .A2(
        npu_inst_pe_1_3_6_n6), .A3(npu_inst_pe_1_3_6_n7), .ZN(
        npu_inst_pe_1_3_6_n44) );
  NAND3_X1 npu_inst_pe_1_3_6_U100 ( .A1(npu_inst_pe_1_3_6_n3), .A2(
        npu_inst_pe_1_3_6_n6), .A3(npu_inst_pe_1_3_6_n7), .ZN(
        npu_inst_pe_1_3_6_n40) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_6_n33), .CK(
        npu_inst_pe_1_3_6_net3788), .RN(npu_inst_pe_1_3_6_n8), .Q(
        npu_inst_int_data_res_3__6__6_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_6_n34), .CK(
        npu_inst_pe_1_3_6_net3788), .RN(npu_inst_pe_1_3_6_n8), .Q(
        npu_inst_int_data_res_3__6__5_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_6_n35), .CK(
        npu_inst_pe_1_3_6_net3788), .RN(npu_inst_pe_1_3_6_n8), .Q(
        npu_inst_int_data_res_3__6__4_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_6_n36), .CK(
        npu_inst_pe_1_3_6_net3788), .RN(npu_inst_pe_1_3_6_n8), .Q(
        npu_inst_int_data_res_3__6__3_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_6_n98), .CK(
        npu_inst_pe_1_3_6_net3788), .RN(npu_inst_pe_1_3_6_n8), .Q(
        npu_inst_int_data_res_3__6__2_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_6_n99), .CK(
        npu_inst_pe_1_3_6_net3788), .RN(npu_inst_pe_1_3_6_n8), .Q(
        npu_inst_int_data_res_3__6__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_6_n32), .CK(
        npu_inst_pe_1_3_6_net3788), .RN(npu_inst_pe_1_3_6_n8), .Q(
        npu_inst_int_data_res_3__6__7_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_6_n100), 
        .CK(npu_inst_pe_1_3_6_net3788), .RN(npu_inst_pe_1_3_6_n8), .Q(
        npu_inst_int_data_res_3__6__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_weight_reg_0_ ( .D(npu_inst_n92), .CK(
        npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n8), .Q(
        npu_inst_pe_1_3_6_int_q_weight_0_), .QN(npu_inst_pe_1_3_6_n27) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_weight_reg_1_ ( .D(npu_inst_n98), .CK(
        npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n8), .Q(
        npu_inst_pe_1_3_6_int_q_weight_1_), .QN(npu_inst_pe_1_3_6_n26) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_6_n112), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n8), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_6_n106), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n8), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_6_n111), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_6_n105), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_6_n110), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_6_n104), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_6_n109), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_6_n103), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_6_n108), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_6_n102), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_6_n107), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_6_n101), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_6_n86), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_6_n87), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n9), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_6_n88), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_6_n89), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_6_n90), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_6_n91), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_6_n92), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_6_n93), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_6_n94), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_6_n95), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_6_n96), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_6_n97), 
        .CK(npu_inst_pe_1_3_6_net3794), .RN(npu_inst_pe_1_3_6_n10), .Q(
        npu_inst_pe_1_3_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_6_net3788) );
  CLKGATETST_X1 npu_inst_pe_1_3_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n46), .SE(1'b0), .GCK(npu_inst_pe_1_3_6_net3794) );
  MUX2_X1 npu_inst_pe_1_3_7_U153 ( .A(npu_inst_pe_1_3_7_n31), .B(
        npu_inst_pe_1_3_7_n28), .S(npu_inst_pe_1_3_7_n7), .Z(
        npu_inst_pe_1_3_7_N93) );
  MUX2_X1 npu_inst_pe_1_3_7_U152 ( .A(npu_inst_pe_1_3_7_n30), .B(
        npu_inst_pe_1_3_7_n29), .S(npu_inst_pe_1_3_7_n5), .Z(
        npu_inst_pe_1_3_7_n31) );
  MUX2_X1 npu_inst_pe_1_3_7_U151 ( .A(npu_inst_pe_1_3_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_3_7_n3), .Z(
        npu_inst_pe_1_3_7_n30) );
  MUX2_X1 npu_inst_pe_1_3_7_U150 ( .A(npu_inst_pe_1_3_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_3_7_n3), .Z(
        npu_inst_pe_1_3_7_n29) );
  MUX2_X1 npu_inst_pe_1_3_7_U149 ( .A(npu_inst_pe_1_3_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_3_7_n3), .Z(
        npu_inst_pe_1_3_7_n28) );
  MUX2_X1 npu_inst_pe_1_3_7_U148 ( .A(npu_inst_pe_1_3_7_n25), .B(
        npu_inst_pe_1_3_7_n22), .S(npu_inst_pe_1_3_7_n7), .Z(
        npu_inst_pe_1_3_7_N94) );
  MUX2_X1 npu_inst_pe_1_3_7_U147 ( .A(npu_inst_pe_1_3_7_n24), .B(
        npu_inst_pe_1_3_7_n23), .S(npu_inst_pe_1_3_7_n5), .Z(
        npu_inst_pe_1_3_7_n25) );
  MUX2_X1 npu_inst_pe_1_3_7_U146 ( .A(npu_inst_pe_1_3_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_3_7_n3), .Z(
        npu_inst_pe_1_3_7_n24) );
  MUX2_X1 npu_inst_pe_1_3_7_U145 ( .A(npu_inst_pe_1_3_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_3_7_n3), .Z(
        npu_inst_pe_1_3_7_n23) );
  MUX2_X1 npu_inst_pe_1_3_7_U144 ( .A(npu_inst_pe_1_3_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_3_7_n3), .Z(
        npu_inst_pe_1_3_7_n22) );
  MUX2_X1 npu_inst_pe_1_3_7_U143 ( .A(npu_inst_pe_1_3_7_n21), .B(
        npu_inst_pe_1_3_7_n18), .S(npu_inst_pe_1_3_7_n7), .Z(
        npu_inst_int_data_x_3__7__1_) );
  MUX2_X1 npu_inst_pe_1_3_7_U142 ( .A(npu_inst_pe_1_3_7_n20), .B(
        npu_inst_pe_1_3_7_n19), .S(npu_inst_pe_1_3_7_n5), .Z(
        npu_inst_pe_1_3_7_n21) );
  MUX2_X1 npu_inst_pe_1_3_7_U141 ( .A(npu_inst_pe_1_3_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_3_7_n3), .Z(
        npu_inst_pe_1_3_7_n20) );
  MUX2_X1 npu_inst_pe_1_3_7_U140 ( .A(npu_inst_pe_1_3_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_3_7_n3), .Z(
        npu_inst_pe_1_3_7_n19) );
  MUX2_X1 npu_inst_pe_1_3_7_U139 ( .A(npu_inst_pe_1_3_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_3_7_n3), .Z(
        npu_inst_pe_1_3_7_n18) );
  MUX2_X1 npu_inst_pe_1_3_7_U138 ( .A(npu_inst_pe_1_3_7_n17), .B(
        npu_inst_pe_1_3_7_n14), .S(npu_inst_pe_1_3_7_n7), .Z(
        npu_inst_int_data_x_3__7__0_) );
  MUX2_X1 npu_inst_pe_1_3_7_U137 ( .A(npu_inst_pe_1_3_7_n16), .B(
        npu_inst_pe_1_3_7_n15), .S(npu_inst_pe_1_3_7_n5), .Z(
        npu_inst_pe_1_3_7_n17) );
  MUX2_X1 npu_inst_pe_1_3_7_U136 ( .A(npu_inst_pe_1_3_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_3_7_n3), .Z(
        npu_inst_pe_1_3_7_n16) );
  MUX2_X1 npu_inst_pe_1_3_7_U135 ( .A(npu_inst_pe_1_3_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_3_7_n3), .Z(
        npu_inst_pe_1_3_7_n15) );
  MUX2_X1 npu_inst_pe_1_3_7_U134 ( .A(npu_inst_pe_1_3_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_3_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_3_7_n3), .Z(
        npu_inst_pe_1_3_7_n14) );
  XOR2_X1 npu_inst_pe_1_3_7_U133 ( .A(npu_inst_pe_1_3_7_int_data_0_), .B(
        npu_inst_int_data_res_3__7__0_), .Z(npu_inst_pe_1_3_7_N73) );
  AND2_X1 npu_inst_pe_1_3_7_U132 ( .A1(npu_inst_int_data_res_3__7__0_), .A2(
        npu_inst_pe_1_3_7_int_data_0_), .ZN(npu_inst_pe_1_3_7_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_3_7_U131 ( .A(npu_inst_int_data_res_3__7__0_), .B(
        npu_inst_pe_1_3_7_n12), .ZN(npu_inst_pe_1_3_7_N65) );
  OR2_X1 npu_inst_pe_1_3_7_U130 ( .A1(npu_inst_pe_1_3_7_n12), .A2(
        npu_inst_int_data_res_3__7__0_), .ZN(npu_inst_pe_1_3_7_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_3_7_U129 ( .A(npu_inst_int_data_res_3__7__2_), .B(
        npu_inst_pe_1_3_7_add_79_carry_2_), .Z(npu_inst_pe_1_3_7_N75) );
  AND2_X1 npu_inst_pe_1_3_7_U128 ( .A1(npu_inst_pe_1_3_7_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_3__7__2_), .ZN(
        npu_inst_pe_1_3_7_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_3_7_U127 ( .A(npu_inst_int_data_res_3__7__3_), .B(
        npu_inst_pe_1_3_7_add_79_carry_3_), .Z(npu_inst_pe_1_3_7_N76) );
  AND2_X1 npu_inst_pe_1_3_7_U126 ( .A1(npu_inst_pe_1_3_7_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_3__7__3_), .ZN(
        npu_inst_pe_1_3_7_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_3_7_U125 ( .A(npu_inst_int_data_res_3__7__4_), .B(
        npu_inst_pe_1_3_7_add_79_carry_4_), .Z(npu_inst_pe_1_3_7_N77) );
  AND2_X1 npu_inst_pe_1_3_7_U124 ( .A1(npu_inst_pe_1_3_7_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_3__7__4_), .ZN(
        npu_inst_pe_1_3_7_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_3_7_U123 ( .A(npu_inst_int_data_res_3__7__5_), .B(
        npu_inst_pe_1_3_7_add_79_carry_5_), .Z(npu_inst_pe_1_3_7_N78) );
  AND2_X1 npu_inst_pe_1_3_7_U122 ( .A1(npu_inst_pe_1_3_7_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_3__7__5_), .ZN(
        npu_inst_pe_1_3_7_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_3_7_U121 ( .A(npu_inst_int_data_res_3__7__6_), .B(
        npu_inst_pe_1_3_7_add_79_carry_6_), .Z(npu_inst_pe_1_3_7_N79) );
  AND2_X1 npu_inst_pe_1_3_7_U120 ( .A1(npu_inst_pe_1_3_7_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_3__7__6_), .ZN(
        npu_inst_pe_1_3_7_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_3_7_U119 ( .A(npu_inst_int_data_res_3__7__7_), .B(
        npu_inst_pe_1_3_7_add_79_carry_7_), .Z(npu_inst_pe_1_3_7_N80) );
  XNOR2_X1 npu_inst_pe_1_3_7_U118 ( .A(npu_inst_pe_1_3_7_sub_77_carry_2_), .B(
        npu_inst_int_data_res_3__7__2_), .ZN(npu_inst_pe_1_3_7_N67) );
  OR2_X1 npu_inst_pe_1_3_7_U117 ( .A1(npu_inst_int_data_res_3__7__2_), .A2(
        npu_inst_pe_1_3_7_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_3_7_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_3_7_U116 ( .A(npu_inst_pe_1_3_7_sub_77_carry_3_), .B(
        npu_inst_int_data_res_3__7__3_), .ZN(npu_inst_pe_1_3_7_N68) );
  OR2_X1 npu_inst_pe_1_3_7_U115 ( .A1(npu_inst_int_data_res_3__7__3_), .A2(
        npu_inst_pe_1_3_7_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_3_7_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_3_7_U114 ( .A(npu_inst_pe_1_3_7_sub_77_carry_4_), .B(
        npu_inst_int_data_res_3__7__4_), .ZN(npu_inst_pe_1_3_7_N69) );
  OR2_X1 npu_inst_pe_1_3_7_U113 ( .A1(npu_inst_int_data_res_3__7__4_), .A2(
        npu_inst_pe_1_3_7_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_3_7_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_3_7_U112 ( .A(npu_inst_pe_1_3_7_sub_77_carry_5_), .B(
        npu_inst_int_data_res_3__7__5_), .ZN(npu_inst_pe_1_3_7_N70) );
  OR2_X1 npu_inst_pe_1_3_7_U111 ( .A1(npu_inst_int_data_res_3__7__5_), .A2(
        npu_inst_pe_1_3_7_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_3_7_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_3_7_U110 ( .A(npu_inst_pe_1_3_7_sub_77_carry_6_), .B(
        npu_inst_int_data_res_3__7__6_), .ZN(npu_inst_pe_1_3_7_N71) );
  OR2_X1 npu_inst_pe_1_3_7_U109 ( .A1(npu_inst_int_data_res_3__7__6_), .A2(
        npu_inst_pe_1_3_7_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_3_7_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_3_7_U108 ( .A(npu_inst_int_data_res_3__7__7_), .B(
        npu_inst_pe_1_3_7_sub_77_carry_7_), .ZN(npu_inst_pe_1_3_7_N72) );
  INV_X1 npu_inst_pe_1_3_7_U107 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_3_7_n6)
         );
  INV_X1 npu_inst_pe_1_3_7_U106 ( .A(npu_inst_pe_1_3_7_n6), .ZN(
        npu_inst_pe_1_3_7_n5) );
  INV_X1 npu_inst_pe_1_3_7_U105 ( .A(npu_inst_n38), .ZN(npu_inst_pe_1_3_7_n2)
         );
  AOI22_X1 npu_inst_pe_1_3_7_U104 ( .A1(npu_inst_int_data_y_4__7__0_), .A2(
        npu_inst_pe_1_3_7_n58), .B1(npu_inst_pe_1_3_7_n118), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_3_7_n57) );
  INV_X1 npu_inst_pe_1_3_7_U103 ( .A(npu_inst_pe_1_3_7_n57), .ZN(
        npu_inst_pe_1_3_7_n107) );
  AOI22_X1 npu_inst_pe_1_3_7_U102 ( .A1(npu_inst_int_data_y_4__7__0_), .A2(
        npu_inst_pe_1_3_7_n54), .B1(npu_inst_pe_1_3_7_n117), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_3_7_n53) );
  INV_X1 npu_inst_pe_1_3_7_U99 ( .A(npu_inst_pe_1_3_7_n53), .ZN(
        npu_inst_pe_1_3_7_n108) );
  AOI22_X1 npu_inst_pe_1_3_7_U98 ( .A1(npu_inst_int_data_y_4__7__0_), .A2(
        npu_inst_pe_1_3_7_n50), .B1(npu_inst_pe_1_3_7_n116), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_3_7_n49) );
  INV_X1 npu_inst_pe_1_3_7_U97 ( .A(npu_inst_pe_1_3_7_n49), .ZN(
        npu_inst_pe_1_3_7_n109) );
  AOI22_X1 npu_inst_pe_1_3_7_U96 ( .A1(npu_inst_int_data_y_4__7__0_), .A2(
        npu_inst_pe_1_3_7_n46), .B1(npu_inst_pe_1_3_7_n115), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_3_7_n45) );
  INV_X1 npu_inst_pe_1_3_7_U95 ( .A(npu_inst_pe_1_3_7_n45), .ZN(
        npu_inst_pe_1_3_7_n110) );
  AOI22_X1 npu_inst_pe_1_3_7_U94 ( .A1(npu_inst_int_data_y_4__7__0_), .A2(
        npu_inst_pe_1_3_7_n42), .B1(npu_inst_pe_1_3_7_n114), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_3_7_n41) );
  INV_X1 npu_inst_pe_1_3_7_U93 ( .A(npu_inst_pe_1_3_7_n41), .ZN(
        npu_inst_pe_1_3_7_n111) );
  AOI22_X1 npu_inst_pe_1_3_7_U92 ( .A1(npu_inst_int_data_y_4__7__1_), .A2(
        npu_inst_pe_1_3_7_n58), .B1(npu_inst_pe_1_3_7_n118), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_3_7_n59) );
  INV_X1 npu_inst_pe_1_3_7_U91 ( .A(npu_inst_pe_1_3_7_n59), .ZN(
        npu_inst_pe_1_3_7_n101) );
  AOI22_X1 npu_inst_pe_1_3_7_U90 ( .A1(npu_inst_int_data_y_4__7__1_), .A2(
        npu_inst_pe_1_3_7_n54), .B1(npu_inst_pe_1_3_7_n117), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_3_7_n55) );
  INV_X1 npu_inst_pe_1_3_7_U89 ( .A(npu_inst_pe_1_3_7_n55), .ZN(
        npu_inst_pe_1_3_7_n102) );
  AOI22_X1 npu_inst_pe_1_3_7_U88 ( .A1(npu_inst_int_data_y_4__7__1_), .A2(
        npu_inst_pe_1_3_7_n50), .B1(npu_inst_pe_1_3_7_n116), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_3_7_n51) );
  INV_X1 npu_inst_pe_1_3_7_U87 ( .A(npu_inst_pe_1_3_7_n51), .ZN(
        npu_inst_pe_1_3_7_n103) );
  AOI22_X1 npu_inst_pe_1_3_7_U86 ( .A1(npu_inst_int_data_y_4__7__1_), .A2(
        npu_inst_pe_1_3_7_n46), .B1(npu_inst_pe_1_3_7_n115), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_3_7_n47) );
  INV_X1 npu_inst_pe_1_3_7_U85 ( .A(npu_inst_pe_1_3_7_n47), .ZN(
        npu_inst_pe_1_3_7_n104) );
  AOI22_X1 npu_inst_pe_1_3_7_U84 ( .A1(npu_inst_int_data_y_4__7__1_), .A2(
        npu_inst_pe_1_3_7_n42), .B1(npu_inst_pe_1_3_7_n114), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_3_7_n43) );
  INV_X1 npu_inst_pe_1_3_7_U83 ( .A(npu_inst_pe_1_3_7_n43), .ZN(
        npu_inst_pe_1_3_7_n105) );
  AOI22_X1 npu_inst_pe_1_3_7_U82 ( .A1(npu_inst_pe_1_3_7_n38), .A2(
        npu_inst_int_data_y_4__7__1_), .B1(npu_inst_pe_1_3_7_n113), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_3_7_n39) );
  INV_X1 npu_inst_pe_1_3_7_U81 ( .A(npu_inst_pe_1_3_7_n39), .ZN(
        npu_inst_pe_1_3_7_n106) );
  AND2_X1 npu_inst_pe_1_3_7_U80 ( .A1(npu_inst_pe_1_3_7_N93), .A2(npu_inst_n38), .ZN(npu_inst_int_data_y_3__7__0_) );
  AOI22_X1 npu_inst_pe_1_3_7_U79 ( .A1(npu_inst_pe_1_3_7_n38), .A2(
        npu_inst_int_data_y_4__7__0_), .B1(npu_inst_pe_1_3_7_n113), .B2(
        npu_inst_pe_1_3_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_3_7_n37) );
  INV_X1 npu_inst_pe_1_3_7_U78 ( .A(npu_inst_pe_1_3_7_n37), .ZN(
        npu_inst_pe_1_3_7_n112) );
  AND2_X1 npu_inst_pe_1_3_7_U77 ( .A1(npu_inst_n38), .A2(npu_inst_pe_1_3_7_N94), .ZN(npu_inst_int_data_y_3__7__1_) );
  AOI222_X1 npu_inst_pe_1_3_7_U76 ( .A1(npu_inst_int_data_res_4__7__0_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N73), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N65), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n84) );
  INV_X1 npu_inst_pe_1_3_7_U75 ( .A(npu_inst_pe_1_3_7_n84), .ZN(
        npu_inst_pe_1_3_7_n100) );
  AOI222_X1 npu_inst_pe_1_3_7_U74 ( .A1(npu_inst_pe_1_3_7_n1), .A2(
        npu_inst_int_data_res_4__7__7_), .B1(npu_inst_pe_1_3_7_N80), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N72), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n75) );
  INV_X1 npu_inst_pe_1_3_7_U73 ( .A(npu_inst_pe_1_3_7_n75), .ZN(
        npu_inst_pe_1_3_7_n32) );
  AOI222_X1 npu_inst_pe_1_3_7_U72 ( .A1(npu_inst_int_data_res_4__7__1_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N74), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N66), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n83) );
  INV_X1 npu_inst_pe_1_3_7_U71 ( .A(npu_inst_pe_1_3_7_n83), .ZN(
        npu_inst_pe_1_3_7_n99) );
  AOI222_X1 npu_inst_pe_1_3_7_U70 ( .A1(npu_inst_int_data_res_4__7__3_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N76), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N68), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n81) );
  INV_X1 npu_inst_pe_1_3_7_U69 ( .A(npu_inst_pe_1_3_7_n81), .ZN(
        npu_inst_pe_1_3_7_n36) );
  AOI222_X1 npu_inst_pe_1_3_7_U68 ( .A1(npu_inst_int_data_res_4__7__4_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N77), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N69), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n80) );
  INV_X1 npu_inst_pe_1_3_7_U67 ( .A(npu_inst_pe_1_3_7_n80), .ZN(
        npu_inst_pe_1_3_7_n35) );
  AOI222_X1 npu_inst_pe_1_3_7_U66 ( .A1(npu_inst_int_data_res_4__7__5_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N78), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N70), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n79) );
  INV_X1 npu_inst_pe_1_3_7_U65 ( .A(npu_inst_pe_1_3_7_n79), .ZN(
        npu_inst_pe_1_3_7_n34) );
  AOI222_X1 npu_inst_pe_1_3_7_U64 ( .A1(npu_inst_int_data_res_4__7__6_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N79), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N71), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n78) );
  INV_X1 npu_inst_pe_1_3_7_U63 ( .A(npu_inst_pe_1_3_7_n78), .ZN(
        npu_inst_pe_1_3_7_n33) );
  AND2_X1 npu_inst_pe_1_3_7_U62 ( .A1(npu_inst_int_data_x_3__7__1_), .A2(
        npu_inst_pe_1_3_7_int_q_weight_1_), .ZN(npu_inst_pe_1_3_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_3_7_U61 ( .A1(npu_inst_int_data_x_3__7__0_), .A2(
        npu_inst_pe_1_3_7_int_q_weight_1_), .ZN(npu_inst_pe_1_3_7_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_3_7_U60 ( .A(npu_inst_pe_1_3_7_int_data_1_), .ZN(
        npu_inst_pe_1_3_7_n13) );
  NAND2_X1 npu_inst_pe_1_3_7_U59 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_3_7_n60), .ZN(npu_inst_pe_1_3_7_n74) );
  OAI21_X1 npu_inst_pe_1_3_7_U58 ( .B1(npu_inst_pe_1_3_7_n63), .B2(
        npu_inst_pe_1_3_7_n60), .A(npu_inst_pe_1_3_7_n74), .ZN(
        npu_inst_pe_1_3_7_n97) );
  NAND2_X1 npu_inst_pe_1_3_7_U57 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_3_7_n60), .ZN(npu_inst_pe_1_3_7_n73) );
  OAI21_X1 npu_inst_pe_1_3_7_U56 ( .B1(npu_inst_pe_1_3_7_n61), .B2(
        npu_inst_pe_1_3_7_n60), .A(npu_inst_pe_1_3_7_n73), .ZN(
        npu_inst_pe_1_3_7_n96) );
  NAND2_X1 npu_inst_pe_1_3_7_U55 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_3_7_n56), .ZN(npu_inst_pe_1_3_7_n72) );
  OAI21_X1 npu_inst_pe_1_3_7_U54 ( .B1(npu_inst_pe_1_3_7_n63), .B2(
        npu_inst_pe_1_3_7_n56), .A(npu_inst_pe_1_3_7_n72), .ZN(
        npu_inst_pe_1_3_7_n95) );
  NAND2_X1 npu_inst_pe_1_3_7_U53 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_3_7_n56), .ZN(npu_inst_pe_1_3_7_n71) );
  OAI21_X1 npu_inst_pe_1_3_7_U52 ( .B1(npu_inst_pe_1_3_7_n61), .B2(
        npu_inst_pe_1_3_7_n56), .A(npu_inst_pe_1_3_7_n71), .ZN(
        npu_inst_pe_1_3_7_n94) );
  NAND2_X1 npu_inst_pe_1_3_7_U51 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_3_7_n52), .ZN(npu_inst_pe_1_3_7_n70) );
  OAI21_X1 npu_inst_pe_1_3_7_U50 ( .B1(npu_inst_pe_1_3_7_n63), .B2(
        npu_inst_pe_1_3_7_n52), .A(npu_inst_pe_1_3_7_n70), .ZN(
        npu_inst_pe_1_3_7_n93) );
  NAND2_X1 npu_inst_pe_1_3_7_U49 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_3_7_n52), .ZN(npu_inst_pe_1_3_7_n69) );
  OAI21_X1 npu_inst_pe_1_3_7_U48 ( .B1(npu_inst_pe_1_3_7_n61), .B2(
        npu_inst_pe_1_3_7_n52), .A(npu_inst_pe_1_3_7_n69), .ZN(
        npu_inst_pe_1_3_7_n92) );
  NAND2_X1 npu_inst_pe_1_3_7_U47 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_3_7_n48), .ZN(npu_inst_pe_1_3_7_n68) );
  OAI21_X1 npu_inst_pe_1_3_7_U46 ( .B1(npu_inst_pe_1_3_7_n63), .B2(
        npu_inst_pe_1_3_7_n48), .A(npu_inst_pe_1_3_7_n68), .ZN(
        npu_inst_pe_1_3_7_n91) );
  NAND2_X1 npu_inst_pe_1_3_7_U45 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_3_7_n48), .ZN(npu_inst_pe_1_3_7_n67) );
  OAI21_X1 npu_inst_pe_1_3_7_U44 ( .B1(npu_inst_pe_1_3_7_n61), .B2(
        npu_inst_pe_1_3_7_n48), .A(npu_inst_pe_1_3_7_n67), .ZN(
        npu_inst_pe_1_3_7_n90) );
  NAND2_X1 npu_inst_pe_1_3_7_U43 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_3_7_n44), .ZN(npu_inst_pe_1_3_7_n66) );
  OAI21_X1 npu_inst_pe_1_3_7_U42 ( .B1(npu_inst_pe_1_3_7_n63), .B2(
        npu_inst_pe_1_3_7_n44), .A(npu_inst_pe_1_3_7_n66), .ZN(
        npu_inst_pe_1_3_7_n89) );
  NAND2_X1 npu_inst_pe_1_3_7_U41 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_3_7_n44), .ZN(npu_inst_pe_1_3_7_n65) );
  OAI21_X1 npu_inst_pe_1_3_7_U40 ( .B1(npu_inst_pe_1_3_7_n61), .B2(
        npu_inst_pe_1_3_7_n44), .A(npu_inst_pe_1_3_7_n65), .ZN(
        npu_inst_pe_1_3_7_n88) );
  NAND2_X1 npu_inst_pe_1_3_7_U39 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_3_7_n40), .ZN(npu_inst_pe_1_3_7_n64) );
  OAI21_X1 npu_inst_pe_1_3_7_U38 ( .B1(npu_inst_pe_1_3_7_n63), .B2(
        npu_inst_pe_1_3_7_n40), .A(npu_inst_pe_1_3_7_n64), .ZN(
        npu_inst_pe_1_3_7_n87) );
  NAND2_X1 npu_inst_pe_1_3_7_U37 ( .A1(npu_inst_pe_1_3_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_3_7_n40), .ZN(npu_inst_pe_1_3_7_n62) );
  OAI21_X1 npu_inst_pe_1_3_7_U36 ( .B1(npu_inst_pe_1_3_7_n61), .B2(
        npu_inst_pe_1_3_7_n40), .A(npu_inst_pe_1_3_7_n62), .ZN(
        npu_inst_pe_1_3_7_n86) );
  NOR3_X1 npu_inst_pe_1_3_7_U35 ( .A1(npu_inst_pe_1_3_7_n26), .A2(npu_inst_n38), .A3(npu_inst_int_ckg[32]), .ZN(npu_inst_pe_1_3_7_n85) );
  OR2_X1 npu_inst_pe_1_3_7_U34 ( .A1(npu_inst_pe_1_3_7_n85), .A2(
        npu_inst_pe_1_3_7_n1), .ZN(npu_inst_pe_1_3_7_N84) );
  AOI222_X1 npu_inst_pe_1_3_7_U33 ( .A1(npu_inst_int_data_res_4__7__2_), .A2(
        npu_inst_pe_1_3_7_n1), .B1(npu_inst_pe_1_3_7_N75), .B2(
        npu_inst_pe_1_3_7_n76), .C1(npu_inst_pe_1_3_7_N67), .C2(
        npu_inst_pe_1_3_7_n77), .ZN(npu_inst_pe_1_3_7_n82) );
  INV_X1 npu_inst_pe_1_3_7_U32 ( .A(npu_inst_pe_1_3_7_n82), .ZN(
        npu_inst_pe_1_3_7_n98) );
  INV_X1 npu_inst_pe_1_3_7_U31 ( .A(npu_inst_pe_1_3_7_int_data_0_), .ZN(
        npu_inst_pe_1_3_7_n12) );
  INV_X1 npu_inst_pe_1_3_7_U30 ( .A(npu_inst_n51), .ZN(npu_inst_pe_1_3_7_n4)
         );
  AOI22_X1 npu_inst_pe_1_3_7_U29 ( .A1(npu_inst_n38), .A2(
        npu_inst_int_data_y_4__7__1_), .B1(npu_inst_pe_1_3_7_n2), .B2(
        int_i_data_h_npu[9]), .ZN(npu_inst_pe_1_3_7_n63) );
  AOI22_X1 npu_inst_pe_1_3_7_U28 ( .A1(npu_inst_n38), .A2(
        npu_inst_int_data_y_4__7__0_), .B1(npu_inst_pe_1_3_7_n2), .B2(
        int_i_data_h_npu[8]), .ZN(npu_inst_pe_1_3_7_n61) );
  OR3_X1 npu_inst_pe_1_3_7_U27 ( .A1(npu_inst_pe_1_3_7_n5), .A2(
        npu_inst_pe_1_3_7_n7), .A3(npu_inst_pe_1_3_7_n4), .ZN(
        npu_inst_pe_1_3_7_n56) );
  OR3_X1 npu_inst_pe_1_3_7_U26 ( .A1(npu_inst_pe_1_3_7_n4), .A2(
        npu_inst_pe_1_3_7_n7), .A3(npu_inst_pe_1_3_7_n6), .ZN(
        npu_inst_pe_1_3_7_n48) );
  INV_X1 npu_inst_pe_1_3_7_U25 ( .A(npu_inst_pe_1_3_7_n4), .ZN(
        npu_inst_pe_1_3_7_n3) );
  OR3_X1 npu_inst_pe_1_3_7_U24 ( .A1(npu_inst_pe_1_3_7_n3), .A2(
        npu_inst_pe_1_3_7_n7), .A3(npu_inst_pe_1_3_7_n6), .ZN(
        npu_inst_pe_1_3_7_n52) );
  OR3_X1 npu_inst_pe_1_3_7_U23 ( .A1(npu_inst_pe_1_3_7_n5), .A2(
        npu_inst_pe_1_3_7_n7), .A3(npu_inst_pe_1_3_7_n3), .ZN(
        npu_inst_pe_1_3_7_n60) );
  BUF_X1 npu_inst_pe_1_3_7_U22 ( .A(npu_inst_n21), .Z(npu_inst_pe_1_3_7_n1) );
  NOR2_X1 npu_inst_pe_1_3_7_U21 ( .A1(npu_inst_pe_1_3_7_n60), .A2(
        npu_inst_pe_1_3_7_n2), .ZN(npu_inst_pe_1_3_7_n58) );
  NOR2_X1 npu_inst_pe_1_3_7_U20 ( .A1(npu_inst_pe_1_3_7_n56), .A2(
        npu_inst_pe_1_3_7_n2), .ZN(npu_inst_pe_1_3_7_n54) );
  NOR2_X1 npu_inst_pe_1_3_7_U19 ( .A1(npu_inst_pe_1_3_7_n52), .A2(
        npu_inst_pe_1_3_7_n2), .ZN(npu_inst_pe_1_3_7_n50) );
  NOR2_X1 npu_inst_pe_1_3_7_U18 ( .A1(npu_inst_pe_1_3_7_n48), .A2(
        npu_inst_pe_1_3_7_n2), .ZN(npu_inst_pe_1_3_7_n46) );
  NOR2_X1 npu_inst_pe_1_3_7_U17 ( .A1(npu_inst_pe_1_3_7_n40), .A2(
        npu_inst_pe_1_3_7_n2), .ZN(npu_inst_pe_1_3_7_n38) );
  NOR2_X1 npu_inst_pe_1_3_7_U16 ( .A1(npu_inst_pe_1_3_7_n44), .A2(
        npu_inst_pe_1_3_7_n2), .ZN(npu_inst_pe_1_3_7_n42) );
  BUF_X1 npu_inst_pe_1_3_7_U15 ( .A(npu_inst_n82), .Z(npu_inst_pe_1_3_7_n7) );
  INV_X1 npu_inst_pe_1_3_7_U14 ( .A(npu_inst_n106), .ZN(npu_inst_pe_1_3_7_n11)
         );
  INV_X1 npu_inst_pe_1_3_7_U13 ( .A(npu_inst_pe_1_3_7_n38), .ZN(
        npu_inst_pe_1_3_7_n113) );
  INV_X1 npu_inst_pe_1_3_7_U12 ( .A(npu_inst_pe_1_3_7_n58), .ZN(
        npu_inst_pe_1_3_7_n118) );
  INV_X1 npu_inst_pe_1_3_7_U11 ( .A(npu_inst_pe_1_3_7_n54), .ZN(
        npu_inst_pe_1_3_7_n117) );
  INV_X1 npu_inst_pe_1_3_7_U10 ( .A(npu_inst_pe_1_3_7_n50), .ZN(
        npu_inst_pe_1_3_7_n116) );
  INV_X1 npu_inst_pe_1_3_7_U9 ( .A(npu_inst_pe_1_3_7_n46), .ZN(
        npu_inst_pe_1_3_7_n115) );
  INV_X1 npu_inst_pe_1_3_7_U8 ( .A(npu_inst_pe_1_3_7_n42), .ZN(
        npu_inst_pe_1_3_7_n114) );
  BUF_X1 npu_inst_pe_1_3_7_U7 ( .A(npu_inst_pe_1_3_7_n11), .Z(
        npu_inst_pe_1_3_7_n10) );
  BUF_X1 npu_inst_pe_1_3_7_U6 ( .A(npu_inst_pe_1_3_7_n11), .Z(
        npu_inst_pe_1_3_7_n9) );
  BUF_X1 npu_inst_pe_1_3_7_U5 ( .A(npu_inst_pe_1_3_7_n11), .Z(
        npu_inst_pe_1_3_7_n8) );
  NOR2_X1 npu_inst_pe_1_3_7_U4 ( .A1(npu_inst_pe_1_3_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_3_7_n1), .ZN(npu_inst_pe_1_3_7_n76) );
  NOR2_X1 npu_inst_pe_1_3_7_U3 ( .A1(npu_inst_pe_1_3_7_n27), .A2(
        npu_inst_pe_1_3_7_n1), .ZN(npu_inst_pe_1_3_7_n77) );
  FA_X1 npu_inst_pe_1_3_7_sub_77_U2_1 ( .A(npu_inst_int_data_res_3__7__1_), 
        .B(npu_inst_pe_1_3_7_n13), .CI(npu_inst_pe_1_3_7_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_3_7_sub_77_carry_2_), .S(npu_inst_pe_1_3_7_N66) );
  FA_X1 npu_inst_pe_1_3_7_add_79_U1_1 ( .A(npu_inst_int_data_res_3__7__1_), 
        .B(npu_inst_pe_1_3_7_int_data_1_), .CI(
        npu_inst_pe_1_3_7_add_79_carry_1_), .CO(
        npu_inst_pe_1_3_7_add_79_carry_2_), .S(npu_inst_pe_1_3_7_N74) );
  NAND3_X1 npu_inst_pe_1_3_7_U101 ( .A1(npu_inst_pe_1_3_7_n4), .A2(
        npu_inst_pe_1_3_7_n6), .A3(npu_inst_pe_1_3_7_n7), .ZN(
        npu_inst_pe_1_3_7_n44) );
  NAND3_X1 npu_inst_pe_1_3_7_U100 ( .A1(npu_inst_pe_1_3_7_n3), .A2(
        npu_inst_pe_1_3_7_n6), .A3(npu_inst_pe_1_3_7_n7), .ZN(
        npu_inst_pe_1_3_7_n40) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_3_7_n33), .CK(
        npu_inst_pe_1_3_7_net3765), .RN(npu_inst_pe_1_3_7_n8), .Q(
        npu_inst_int_data_res_3__7__6_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_3_7_n34), .CK(
        npu_inst_pe_1_3_7_net3765), .RN(npu_inst_pe_1_3_7_n8), .Q(
        npu_inst_int_data_res_3__7__5_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_3_7_n35), .CK(
        npu_inst_pe_1_3_7_net3765), .RN(npu_inst_pe_1_3_7_n8), .Q(
        npu_inst_int_data_res_3__7__4_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_3_7_n36), .CK(
        npu_inst_pe_1_3_7_net3765), .RN(npu_inst_pe_1_3_7_n8), .Q(
        npu_inst_int_data_res_3__7__3_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_3_7_n98), .CK(
        npu_inst_pe_1_3_7_net3765), .RN(npu_inst_pe_1_3_7_n8), .Q(
        npu_inst_int_data_res_3__7__2_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_3_7_n99), .CK(
        npu_inst_pe_1_3_7_net3765), .RN(npu_inst_pe_1_3_7_n8), .Q(
        npu_inst_int_data_res_3__7__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_3_7_n32), .CK(
        npu_inst_pe_1_3_7_net3765), .RN(npu_inst_pe_1_3_7_n8), .Q(
        npu_inst_int_data_res_3__7__7_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_3_7_n100), 
        .CK(npu_inst_pe_1_3_7_net3765), .RN(npu_inst_pe_1_3_7_n8), .Q(
        npu_inst_int_data_res_3__7__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_weight_reg_0_ ( .D(npu_inst_n92), .CK(
        npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n8), .Q(
        npu_inst_pe_1_3_7_int_q_weight_0_), .QN(npu_inst_pe_1_3_7_n27) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_weight_reg_1_ ( .D(npu_inst_n98), .CK(
        npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n8), .Q(
        npu_inst_pe_1_3_7_int_q_weight_1_), .QN(npu_inst_pe_1_3_7_n26) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_3_7_n112), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n8), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_3_7_n106), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n8), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_3_7_n111), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_3_7_n105), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_3_7_n110), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_3_7_n104), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_3_7_n109), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_3_7_n103), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_3_7_n108), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_3_7_n102), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_3_7_n107), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_3_7_n101), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_3_7_n86), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_3_7_n87), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n9), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_3_7_n88), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_3_7_n89), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_3_7_n90), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_3_7_n91), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_3_7_n92), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_3_7_n93), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_3_7_n94), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_3_7_n95), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_3_7_n96), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_3_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_3_7_n97), 
        .CK(npu_inst_pe_1_3_7_net3771), .RN(npu_inst_pe_1_3_7_n10), .Q(
        npu_inst_pe_1_3_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_3_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_3_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_3_7_net3765) );
  CLKGATETST_X1 npu_inst_pe_1_3_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n45), .SE(1'b0), .GCK(npu_inst_pe_1_3_7_net3771) );
  MUX2_X1 npu_inst_pe_1_4_0_U153 ( .A(npu_inst_pe_1_4_0_n31), .B(
        npu_inst_pe_1_4_0_n28), .S(npu_inst_pe_1_4_0_n7), .Z(
        npu_inst_pe_1_4_0_N93) );
  MUX2_X1 npu_inst_pe_1_4_0_U152 ( .A(npu_inst_pe_1_4_0_n30), .B(
        npu_inst_pe_1_4_0_n29), .S(npu_inst_pe_1_4_0_n5), .Z(
        npu_inst_pe_1_4_0_n31) );
  MUX2_X1 npu_inst_pe_1_4_0_U151 ( .A(npu_inst_pe_1_4_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_0_n3), .Z(
        npu_inst_pe_1_4_0_n30) );
  MUX2_X1 npu_inst_pe_1_4_0_U150 ( .A(npu_inst_pe_1_4_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_0_n3), .Z(
        npu_inst_pe_1_4_0_n29) );
  MUX2_X1 npu_inst_pe_1_4_0_U149 ( .A(npu_inst_pe_1_4_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_0_n3), .Z(
        npu_inst_pe_1_4_0_n28) );
  MUX2_X1 npu_inst_pe_1_4_0_U148 ( .A(npu_inst_pe_1_4_0_n25), .B(
        npu_inst_pe_1_4_0_n22), .S(npu_inst_pe_1_4_0_n7), .Z(
        npu_inst_pe_1_4_0_N94) );
  MUX2_X1 npu_inst_pe_1_4_0_U147 ( .A(npu_inst_pe_1_4_0_n24), .B(
        npu_inst_pe_1_4_0_n23), .S(npu_inst_pe_1_4_0_n5), .Z(
        npu_inst_pe_1_4_0_n25) );
  MUX2_X1 npu_inst_pe_1_4_0_U146 ( .A(npu_inst_pe_1_4_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_0_n3), .Z(
        npu_inst_pe_1_4_0_n24) );
  MUX2_X1 npu_inst_pe_1_4_0_U145 ( .A(npu_inst_pe_1_4_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_0_n3), .Z(
        npu_inst_pe_1_4_0_n23) );
  MUX2_X1 npu_inst_pe_1_4_0_U144 ( .A(npu_inst_pe_1_4_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_0_n3), .Z(
        npu_inst_pe_1_4_0_n22) );
  MUX2_X1 npu_inst_pe_1_4_0_U143 ( .A(npu_inst_pe_1_4_0_n21), .B(
        npu_inst_pe_1_4_0_n18), .S(npu_inst_pe_1_4_0_n7), .Z(
        npu_inst_pe_1_4_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_4_0_U142 ( .A(npu_inst_pe_1_4_0_n20), .B(
        npu_inst_pe_1_4_0_n19), .S(npu_inst_pe_1_4_0_n5), .Z(
        npu_inst_pe_1_4_0_n21) );
  MUX2_X1 npu_inst_pe_1_4_0_U141 ( .A(npu_inst_pe_1_4_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_0_n3), .Z(
        npu_inst_pe_1_4_0_n20) );
  MUX2_X1 npu_inst_pe_1_4_0_U140 ( .A(npu_inst_pe_1_4_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_0_n3), .Z(
        npu_inst_pe_1_4_0_n19) );
  MUX2_X1 npu_inst_pe_1_4_0_U139 ( .A(npu_inst_pe_1_4_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_0_n3), .Z(
        npu_inst_pe_1_4_0_n18) );
  MUX2_X1 npu_inst_pe_1_4_0_U138 ( .A(npu_inst_pe_1_4_0_n17), .B(
        npu_inst_pe_1_4_0_n14), .S(npu_inst_pe_1_4_0_n7), .Z(
        npu_inst_pe_1_4_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_4_0_U137 ( .A(npu_inst_pe_1_4_0_n16), .B(
        npu_inst_pe_1_4_0_n15), .S(npu_inst_pe_1_4_0_n5), .Z(
        npu_inst_pe_1_4_0_n17) );
  MUX2_X1 npu_inst_pe_1_4_0_U136 ( .A(npu_inst_pe_1_4_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_0_n3), .Z(
        npu_inst_pe_1_4_0_n16) );
  MUX2_X1 npu_inst_pe_1_4_0_U135 ( .A(npu_inst_pe_1_4_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_0_n3), .Z(
        npu_inst_pe_1_4_0_n15) );
  MUX2_X1 npu_inst_pe_1_4_0_U134 ( .A(npu_inst_pe_1_4_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_0_n3), .Z(
        npu_inst_pe_1_4_0_n14) );
  XOR2_X1 npu_inst_pe_1_4_0_U133 ( .A(npu_inst_pe_1_4_0_int_data_0_), .B(
        npu_inst_int_data_res_4__0__0_), .Z(npu_inst_pe_1_4_0_N73) );
  AND2_X1 npu_inst_pe_1_4_0_U132 ( .A1(npu_inst_int_data_res_4__0__0_), .A2(
        npu_inst_pe_1_4_0_int_data_0_), .ZN(npu_inst_pe_1_4_0_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_0_U131 ( .A(npu_inst_int_data_res_4__0__0_), .B(
        npu_inst_pe_1_4_0_n12), .ZN(npu_inst_pe_1_4_0_N65) );
  OR2_X1 npu_inst_pe_1_4_0_U130 ( .A1(npu_inst_pe_1_4_0_n12), .A2(
        npu_inst_int_data_res_4__0__0_), .ZN(npu_inst_pe_1_4_0_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_0_U129 ( .A(npu_inst_int_data_res_4__0__2_), .B(
        npu_inst_pe_1_4_0_add_79_carry_2_), .Z(npu_inst_pe_1_4_0_N75) );
  AND2_X1 npu_inst_pe_1_4_0_U128 ( .A1(npu_inst_pe_1_4_0_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_4__0__2_), .ZN(
        npu_inst_pe_1_4_0_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_0_U127 ( .A(npu_inst_int_data_res_4__0__3_), .B(
        npu_inst_pe_1_4_0_add_79_carry_3_), .Z(npu_inst_pe_1_4_0_N76) );
  AND2_X1 npu_inst_pe_1_4_0_U126 ( .A1(npu_inst_pe_1_4_0_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_4__0__3_), .ZN(
        npu_inst_pe_1_4_0_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_0_U125 ( .A(npu_inst_int_data_res_4__0__4_), .B(
        npu_inst_pe_1_4_0_add_79_carry_4_), .Z(npu_inst_pe_1_4_0_N77) );
  AND2_X1 npu_inst_pe_1_4_0_U124 ( .A1(npu_inst_pe_1_4_0_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_4__0__4_), .ZN(
        npu_inst_pe_1_4_0_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_0_U123 ( .A(npu_inst_int_data_res_4__0__5_), .B(
        npu_inst_pe_1_4_0_add_79_carry_5_), .Z(npu_inst_pe_1_4_0_N78) );
  AND2_X1 npu_inst_pe_1_4_0_U122 ( .A1(npu_inst_pe_1_4_0_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_4__0__5_), .ZN(
        npu_inst_pe_1_4_0_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_0_U121 ( .A(npu_inst_int_data_res_4__0__6_), .B(
        npu_inst_pe_1_4_0_add_79_carry_6_), .Z(npu_inst_pe_1_4_0_N79) );
  AND2_X1 npu_inst_pe_1_4_0_U120 ( .A1(npu_inst_pe_1_4_0_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_4__0__6_), .ZN(
        npu_inst_pe_1_4_0_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_0_U119 ( .A(npu_inst_int_data_res_4__0__7_), .B(
        npu_inst_pe_1_4_0_add_79_carry_7_), .Z(npu_inst_pe_1_4_0_N80) );
  XNOR2_X1 npu_inst_pe_1_4_0_U118 ( .A(npu_inst_pe_1_4_0_sub_77_carry_2_), .B(
        npu_inst_int_data_res_4__0__2_), .ZN(npu_inst_pe_1_4_0_N67) );
  OR2_X1 npu_inst_pe_1_4_0_U117 ( .A1(npu_inst_int_data_res_4__0__2_), .A2(
        npu_inst_pe_1_4_0_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_4_0_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_0_U116 ( .A(npu_inst_pe_1_4_0_sub_77_carry_3_), .B(
        npu_inst_int_data_res_4__0__3_), .ZN(npu_inst_pe_1_4_0_N68) );
  OR2_X1 npu_inst_pe_1_4_0_U115 ( .A1(npu_inst_int_data_res_4__0__3_), .A2(
        npu_inst_pe_1_4_0_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_4_0_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_0_U114 ( .A(npu_inst_pe_1_4_0_sub_77_carry_4_), .B(
        npu_inst_int_data_res_4__0__4_), .ZN(npu_inst_pe_1_4_0_N69) );
  OR2_X1 npu_inst_pe_1_4_0_U113 ( .A1(npu_inst_int_data_res_4__0__4_), .A2(
        npu_inst_pe_1_4_0_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_4_0_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_0_U112 ( .A(npu_inst_pe_1_4_0_sub_77_carry_5_), .B(
        npu_inst_int_data_res_4__0__5_), .ZN(npu_inst_pe_1_4_0_N70) );
  OR2_X1 npu_inst_pe_1_4_0_U111 ( .A1(npu_inst_int_data_res_4__0__5_), .A2(
        npu_inst_pe_1_4_0_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_4_0_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_0_U110 ( .A(npu_inst_pe_1_4_0_sub_77_carry_6_), .B(
        npu_inst_int_data_res_4__0__6_), .ZN(npu_inst_pe_1_4_0_N71) );
  OR2_X1 npu_inst_pe_1_4_0_U109 ( .A1(npu_inst_int_data_res_4__0__6_), .A2(
        npu_inst_pe_1_4_0_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_4_0_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_0_U108 ( .A(npu_inst_int_data_res_4__0__7_), .B(
        npu_inst_pe_1_4_0_sub_77_carry_7_), .ZN(npu_inst_pe_1_4_0_N72) );
  INV_X1 npu_inst_pe_1_4_0_U107 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_4_0_n6)
         );
  INV_X1 npu_inst_pe_1_4_0_U106 ( .A(npu_inst_pe_1_4_0_n6), .ZN(
        npu_inst_pe_1_4_0_n5) );
  INV_X1 npu_inst_pe_1_4_0_U105 ( .A(npu_inst_n38), .ZN(npu_inst_pe_1_4_0_n2)
         );
  AOI22_X1 npu_inst_pe_1_4_0_U104 ( .A1(npu_inst_int_data_y_5__0__0_), .A2(
        npu_inst_pe_1_4_0_n58), .B1(npu_inst_pe_1_4_0_n118), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_0_n57) );
  INV_X1 npu_inst_pe_1_4_0_U103 ( .A(npu_inst_pe_1_4_0_n57), .ZN(
        npu_inst_pe_1_4_0_n107) );
  AOI22_X1 npu_inst_pe_1_4_0_U102 ( .A1(npu_inst_int_data_y_5__0__0_), .A2(
        npu_inst_pe_1_4_0_n54), .B1(npu_inst_pe_1_4_0_n117), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_0_n53) );
  INV_X1 npu_inst_pe_1_4_0_U99 ( .A(npu_inst_pe_1_4_0_n53), .ZN(
        npu_inst_pe_1_4_0_n108) );
  AOI22_X1 npu_inst_pe_1_4_0_U98 ( .A1(npu_inst_int_data_y_5__0__0_), .A2(
        npu_inst_pe_1_4_0_n50), .B1(npu_inst_pe_1_4_0_n116), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_0_n49) );
  INV_X1 npu_inst_pe_1_4_0_U97 ( .A(npu_inst_pe_1_4_0_n49), .ZN(
        npu_inst_pe_1_4_0_n109) );
  AOI22_X1 npu_inst_pe_1_4_0_U96 ( .A1(npu_inst_int_data_y_5__0__0_), .A2(
        npu_inst_pe_1_4_0_n46), .B1(npu_inst_pe_1_4_0_n115), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_0_n45) );
  INV_X1 npu_inst_pe_1_4_0_U95 ( .A(npu_inst_pe_1_4_0_n45), .ZN(
        npu_inst_pe_1_4_0_n110) );
  AOI22_X1 npu_inst_pe_1_4_0_U94 ( .A1(npu_inst_int_data_y_5__0__0_), .A2(
        npu_inst_pe_1_4_0_n42), .B1(npu_inst_pe_1_4_0_n114), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_0_n41) );
  INV_X1 npu_inst_pe_1_4_0_U93 ( .A(npu_inst_pe_1_4_0_n41), .ZN(
        npu_inst_pe_1_4_0_n111) );
  AOI22_X1 npu_inst_pe_1_4_0_U92 ( .A1(npu_inst_int_data_y_5__0__1_), .A2(
        npu_inst_pe_1_4_0_n58), .B1(npu_inst_pe_1_4_0_n118), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_0_n59) );
  INV_X1 npu_inst_pe_1_4_0_U91 ( .A(npu_inst_pe_1_4_0_n59), .ZN(
        npu_inst_pe_1_4_0_n101) );
  AOI22_X1 npu_inst_pe_1_4_0_U90 ( .A1(npu_inst_int_data_y_5__0__1_), .A2(
        npu_inst_pe_1_4_0_n54), .B1(npu_inst_pe_1_4_0_n117), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_0_n55) );
  INV_X1 npu_inst_pe_1_4_0_U89 ( .A(npu_inst_pe_1_4_0_n55), .ZN(
        npu_inst_pe_1_4_0_n102) );
  AOI22_X1 npu_inst_pe_1_4_0_U88 ( .A1(npu_inst_int_data_y_5__0__1_), .A2(
        npu_inst_pe_1_4_0_n50), .B1(npu_inst_pe_1_4_0_n116), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_0_n51) );
  INV_X1 npu_inst_pe_1_4_0_U87 ( .A(npu_inst_pe_1_4_0_n51), .ZN(
        npu_inst_pe_1_4_0_n103) );
  AOI22_X1 npu_inst_pe_1_4_0_U86 ( .A1(npu_inst_int_data_y_5__0__1_), .A2(
        npu_inst_pe_1_4_0_n46), .B1(npu_inst_pe_1_4_0_n115), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_0_n47) );
  INV_X1 npu_inst_pe_1_4_0_U85 ( .A(npu_inst_pe_1_4_0_n47), .ZN(
        npu_inst_pe_1_4_0_n104) );
  AOI22_X1 npu_inst_pe_1_4_0_U84 ( .A1(npu_inst_int_data_y_5__0__1_), .A2(
        npu_inst_pe_1_4_0_n42), .B1(npu_inst_pe_1_4_0_n114), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_0_n43) );
  INV_X1 npu_inst_pe_1_4_0_U83 ( .A(npu_inst_pe_1_4_0_n43), .ZN(
        npu_inst_pe_1_4_0_n105) );
  AOI22_X1 npu_inst_pe_1_4_0_U82 ( .A1(npu_inst_pe_1_4_0_n38), .A2(
        npu_inst_int_data_y_5__0__1_), .B1(npu_inst_pe_1_4_0_n113), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_0_n39) );
  INV_X1 npu_inst_pe_1_4_0_U81 ( .A(npu_inst_pe_1_4_0_n39), .ZN(
        npu_inst_pe_1_4_0_n106) );
  AND2_X1 npu_inst_pe_1_4_0_U80 ( .A1(npu_inst_pe_1_4_0_N93), .A2(npu_inst_n38), .ZN(npu_inst_int_data_y_4__0__0_) );
  NAND2_X1 npu_inst_pe_1_4_0_U79 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_0_n60), .ZN(npu_inst_pe_1_4_0_n74) );
  OAI21_X1 npu_inst_pe_1_4_0_U78 ( .B1(npu_inst_pe_1_4_0_n63), .B2(
        npu_inst_pe_1_4_0_n60), .A(npu_inst_pe_1_4_0_n74), .ZN(
        npu_inst_pe_1_4_0_n97) );
  NAND2_X1 npu_inst_pe_1_4_0_U77 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_0_n60), .ZN(npu_inst_pe_1_4_0_n73) );
  OAI21_X1 npu_inst_pe_1_4_0_U76 ( .B1(npu_inst_pe_1_4_0_n61), .B2(
        npu_inst_pe_1_4_0_n60), .A(npu_inst_pe_1_4_0_n73), .ZN(
        npu_inst_pe_1_4_0_n96) );
  NAND2_X1 npu_inst_pe_1_4_0_U75 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_0_n56), .ZN(npu_inst_pe_1_4_0_n72) );
  OAI21_X1 npu_inst_pe_1_4_0_U74 ( .B1(npu_inst_pe_1_4_0_n63), .B2(
        npu_inst_pe_1_4_0_n56), .A(npu_inst_pe_1_4_0_n72), .ZN(
        npu_inst_pe_1_4_0_n95) );
  NAND2_X1 npu_inst_pe_1_4_0_U73 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_0_n56), .ZN(npu_inst_pe_1_4_0_n71) );
  OAI21_X1 npu_inst_pe_1_4_0_U72 ( .B1(npu_inst_pe_1_4_0_n61), .B2(
        npu_inst_pe_1_4_0_n56), .A(npu_inst_pe_1_4_0_n71), .ZN(
        npu_inst_pe_1_4_0_n94) );
  NAND2_X1 npu_inst_pe_1_4_0_U71 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_0_n52), .ZN(npu_inst_pe_1_4_0_n70) );
  OAI21_X1 npu_inst_pe_1_4_0_U70 ( .B1(npu_inst_pe_1_4_0_n63), .B2(
        npu_inst_pe_1_4_0_n52), .A(npu_inst_pe_1_4_0_n70), .ZN(
        npu_inst_pe_1_4_0_n93) );
  NAND2_X1 npu_inst_pe_1_4_0_U69 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_0_n52), .ZN(npu_inst_pe_1_4_0_n69) );
  OAI21_X1 npu_inst_pe_1_4_0_U68 ( .B1(npu_inst_pe_1_4_0_n61), .B2(
        npu_inst_pe_1_4_0_n52), .A(npu_inst_pe_1_4_0_n69), .ZN(
        npu_inst_pe_1_4_0_n92) );
  NAND2_X1 npu_inst_pe_1_4_0_U67 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_0_n48), .ZN(npu_inst_pe_1_4_0_n68) );
  OAI21_X1 npu_inst_pe_1_4_0_U66 ( .B1(npu_inst_pe_1_4_0_n63), .B2(
        npu_inst_pe_1_4_0_n48), .A(npu_inst_pe_1_4_0_n68), .ZN(
        npu_inst_pe_1_4_0_n91) );
  NAND2_X1 npu_inst_pe_1_4_0_U65 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_0_n48), .ZN(npu_inst_pe_1_4_0_n67) );
  OAI21_X1 npu_inst_pe_1_4_0_U64 ( .B1(npu_inst_pe_1_4_0_n61), .B2(
        npu_inst_pe_1_4_0_n48), .A(npu_inst_pe_1_4_0_n67), .ZN(
        npu_inst_pe_1_4_0_n90) );
  NAND2_X1 npu_inst_pe_1_4_0_U63 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_0_n44), .ZN(npu_inst_pe_1_4_0_n66) );
  OAI21_X1 npu_inst_pe_1_4_0_U62 ( .B1(npu_inst_pe_1_4_0_n63), .B2(
        npu_inst_pe_1_4_0_n44), .A(npu_inst_pe_1_4_0_n66), .ZN(
        npu_inst_pe_1_4_0_n89) );
  NAND2_X1 npu_inst_pe_1_4_0_U61 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_0_n44), .ZN(npu_inst_pe_1_4_0_n65) );
  OAI21_X1 npu_inst_pe_1_4_0_U60 ( .B1(npu_inst_pe_1_4_0_n61), .B2(
        npu_inst_pe_1_4_0_n44), .A(npu_inst_pe_1_4_0_n65), .ZN(
        npu_inst_pe_1_4_0_n88) );
  NAND2_X1 npu_inst_pe_1_4_0_U59 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_0_n40), .ZN(npu_inst_pe_1_4_0_n64) );
  OAI21_X1 npu_inst_pe_1_4_0_U58 ( .B1(npu_inst_pe_1_4_0_n63), .B2(
        npu_inst_pe_1_4_0_n40), .A(npu_inst_pe_1_4_0_n64), .ZN(
        npu_inst_pe_1_4_0_n87) );
  NAND2_X1 npu_inst_pe_1_4_0_U57 ( .A1(npu_inst_pe_1_4_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_0_n40), .ZN(npu_inst_pe_1_4_0_n62) );
  OAI21_X1 npu_inst_pe_1_4_0_U56 ( .B1(npu_inst_pe_1_4_0_n61), .B2(
        npu_inst_pe_1_4_0_n40), .A(npu_inst_pe_1_4_0_n62), .ZN(
        npu_inst_pe_1_4_0_n86) );
  AOI22_X1 npu_inst_pe_1_4_0_U55 ( .A1(npu_inst_pe_1_4_0_n38), .A2(
        npu_inst_int_data_y_5__0__0_), .B1(npu_inst_pe_1_4_0_n113), .B2(
        npu_inst_pe_1_4_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_0_n37) );
  INV_X1 npu_inst_pe_1_4_0_U54 ( .A(npu_inst_pe_1_4_0_n37), .ZN(
        npu_inst_pe_1_4_0_n112) );
  NOR3_X1 npu_inst_pe_1_4_0_U53 ( .A1(npu_inst_pe_1_4_0_n26), .A2(npu_inst_n38), .A3(npu_inst_int_ckg[31]), .ZN(npu_inst_pe_1_4_0_n85) );
  OR2_X1 npu_inst_pe_1_4_0_U52 ( .A1(npu_inst_pe_1_4_0_n85), .A2(
        npu_inst_pe_1_4_0_n1), .ZN(npu_inst_pe_1_4_0_N84) );
  AND2_X1 npu_inst_pe_1_4_0_U51 ( .A1(npu_inst_n38), .A2(npu_inst_pe_1_4_0_N94), .ZN(npu_inst_int_data_y_4__0__1_) );
  AOI222_X1 npu_inst_pe_1_4_0_U50 ( .A1(npu_inst_int_data_res_5__0__0_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N73), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N65), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n84) );
  INV_X1 npu_inst_pe_1_4_0_U49 ( .A(npu_inst_pe_1_4_0_n84), .ZN(
        npu_inst_pe_1_4_0_n100) );
  AOI222_X1 npu_inst_pe_1_4_0_U48 ( .A1(npu_inst_pe_1_4_0_n1), .A2(
        npu_inst_int_data_res_5__0__7_), .B1(npu_inst_pe_1_4_0_N80), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N72), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n75) );
  INV_X1 npu_inst_pe_1_4_0_U47 ( .A(npu_inst_pe_1_4_0_n75), .ZN(
        npu_inst_pe_1_4_0_n32) );
  AOI222_X1 npu_inst_pe_1_4_0_U46 ( .A1(npu_inst_int_data_res_5__0__1_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N74), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N66), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n83) );
  INV_X1 npu_inst_pe_1_4_0_U45 ( .A(npu_inst_pe_1_4_0_n83), .ZN(
        npu_inst_pe_1_4_0_n99) );
  AOI222_X1 npu_inst_pe_1_4_0_U44 ( .A1(npu_inst_int_data_res_5__0__3_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N76), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N68), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n81) );
  INV_X1 npu_inst_pe_1_4_0_U43 ( .A(npu_inst_pe_1_4_0_n81), .ZN(
        npu_inst_pe_1_4_0_n36) );
  AOI222_X1 npu_inst_pe_1_4_0_U42 ( .A1(npu_inst_int_data_res_5__0__4_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N77), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N69), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n80) );
  INV_X1 npu_inst_pe_1_4_0_U41 ( .A(npu_inst_pe_1_4_0_n80), .ZN(
        npu_inst_pe_1_4_0_n35) );
  AOI222_X1 npu_inst_pe_1_4_0_U40 ( .A1(npu_inst_int_data_res_5__0__5_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N78), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N70), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n79) );
  INV_X1 npu_inst_pe_1_4_0_U39 ( .A(npu_inst_pe_1_4_0_n79), .ZN(
        npu_inst_pe_1_4_0_n34) );
  AOI222_X1 npu_inst_pe_1_4_0_U38 ( .A1(npu_inst_int_data_res_5__0__6_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N79), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N71), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n78) );
  INV_X1 npu_inst_pe_1_4_0_U37 ( .A(npu_inst_pe_1_4_0_n78), .ZN(
        npu_inst_pe_1_4_0_n33) );
  AND2_X1 npu_inst_pe_1_4_0_U36 ( .A1(npu_inst_pe_1_4_0_o_data_h_1_), .A2(
        npu_inst_pe_1_4_0_int_q_weight_1_), .ZN(npu_inst_pe_1_4_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_0_U35 ( .A1(npu_inst_pe_1_4_0_o_data_h_0_), .A2(
        npu_inst_pe_1_4_0_int_q_weight_1_), .ZN(npu_inst_pe_1_4_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_4_0_U34 ( .A(npu_inst_pe_1_4_0_int_data_1_), .ZN(
        npu_inst_pe_1_4_0_n13) );
  AOI222_X1 npu_inst_pe_1_4_0_U33 ( .A1(npu_inst_int_data_res_5__0__2_), .A2(
        npu_inst_pe_1_4_0_n1), .B1(npu_inst_pe_1_4_0_N75), .B2(
        npu_inst_pe_1_4_0_n76), .C1(npu_inst_pe_1_4_0_N67), .C2(
        npu_inst_pe_1_4_0_n77), .ZN(npu_inst_pe_1_4_0_n82) );
  INV_X1 npu_inst_pe_1_4_0_U32 ( .A(npu_inst_pe_1_4_0_n82), .ZN(
        npu_inst_pe_1_4_0_n98) );
  AOI22_X1 npu_inst_pe_1_4_0_U31 ( .A1(npu_inst_n38), .A2(
        npu_inst_int_data_y_5__0__1_), .B1(npu_inst_pe_1_4_0_n2), .B2(
        npu_inst_int_data_x_4__1__1_), .ZN(npu_inst_pe_1_4_0_n63) );
  AOI22_X1 npu_inst_pe_1_4_0_U30 ( .A1(npu_inst_n38), .A2(
        npu_inst_int_data_y_5__0__0_), .B1(npu_inst_pe_1_4_0_n2), .B2(
        npu_inst_int_data_x_4__1__0_), .ZN(npu_inst_pe_1_4_0_n61) );
  INV_X1 npu_inst_pe_1_4_0_U29 ( .A(npu_inst_pe_1_4_0_int_data_0_), .ZN(
        npu_inst_pe_1_4_0_n12) );
  INV_X1 npu_inst_pe_1_4_0_U28 ( .A(npu_inst_n51), .ZN(npu_inst_pe_1_4_0_n4)
         );
  OR3_X1 npu_inst_pe_1_4_0_U27 ( .A1(npu_inst_pe_1_4_0_n5), .A2(
        npu_inst_pe_1_4_0_n7), .A3(npu_inst_pe_1_4_0_n4), .ZN(
        npu_inst_pe_1_4_0_n56) );
  OR3_X1 npu_inst_pe_1_4_0_U26 ( .A1(npu_inst_pe_1_4_0_n4), .A2(
        npu_inst_pe_1_4_0_n7), .A3(npu_inst_pe_1_4_0_n6), .ZN(
        npu_inst_pe_1_4_0_n48) );
  INV_X1 npu_inst_pe_1_4_0_U25 ( .A(npu_inst_pe_1_4_0_n4), .ZN(
        npu_inst_pe_1_4_0_n3) );
  OR3_X1 npu_inst_pe_1_4_0_U24 ( .A1(npu_inst_pe_1_4_0_n3), .A2(
        npu_inst_pe_1_4_0_n7), .A3(npu_inst_pe_1_4_0_n6), .ZN(
        npu_inst_pe_1_4_0_n52) );
  OR3_X1 npu_inst_pe_1_4_0_U23 ( .A1(npu_inst_pe_1_4_0_n5), .A2(
        npu_inst_pe_1_4_0_n7), .A3(npu_inst_pe_1_4_0_n3), .ZN(
        npu_inst_pe_1_4_0_n60) );
  BUF_X1 npu_inst_pe_1_4_0_U22 ( .A(npu_inst_n21), .Z(npu_inst_pe_1_4_0_n1) );
  NOR2_X1 npu_inst_pe_1_4_0_U21 ( .A1(npu_inst_pe_1_4_0_n60), .A2(
        npu_inst_pe_1_4_0_n2), .ZN(npu_inst_pe_1_4_0_n58) );
  NOR2_X1 npu_inst_pe_1_4_0_U20 ( .A1(npu_inst_pe_1_4_0_n56), .A2(
        npu_inst_pe_1_4_0_n2), .ZN(npu_inst_pe_1_4_0_n54) );
  NOR2_X1 npu_inst_pe_1_4_0_U19 ( .A1(npu_inst_pe_1_4_0_n52), .A2(
        npu_inst_pe_1_4_0_n2), .ZN(npu_inst_pe_1_4_0_n50) );
  NOR2_X1 npu_inst_pe_1_4_0_U18 ( .A1(npu_inst_pe_1_4_0_n48), .A2(
        npu_inst_pe_1_4_0_n2), .ZN(npu_inst_pe_1_4_0_n46) );
  NOR2_X1 npu_inst_pe_1_4_0_U17 ( .A1(npu_inst_pe_1_4_0_n40), .A2(
        npu_inst_pe_1_4_0_n2), .ZN(npu_inst_pe_1_4_0_n38) );
  NOR2_X1 npu_inst_pe_1_4_0_U16 ( .A1(npu_inst_pe_1_4_0_n44), .A2(
        npu_inst_pe_1_4_0_n2), .ZN(npu_inst_pe_1_4_0_n42) );
  BUF_X1 npu_inst_pe_1_4_0_U15 ( .A(npu_inst_n81), .Z(npu_inst_pe_1_4_0_n7) );
  INV_X1 npu_inst_pe_1_4_0_U14 ( .A(npu_inst_n106), .ZN(npu_inst_pe_1_4_0_n11)
         );
  INV_X1 npu_inst_pe_1_4_0_U13 ( .A(npu_inst_pe_1_4_0_n38), .ZN(
        npu_inst_pe_1_4_0_n113) );
  INV_X1 npu_inst_pe_1_4_0_U12 ( .A(npu_inst_pe_1_4_0_n58), .ZN(
        npu_inst_pe_1_4_0_n118) );
  INV_X1 npu_inst_pe_1_4_0_U11 ( .A(npu_inst_pe_1_4_0_n54), .ZN(
        npu_inst_pe_1_4_0_n117) );
  INV_X1 npu_inst_pe_1_4_0_U10 ( .A(npu_inst_pe_1_4_0_n50), .ZN(
        npu_inst_pe_1_4_0_n116) );
  INV_X1 npu_inst_pe_1_4_0_U9 ( .A(npu_inst_pe_1_4_0_n46), .ZN(
        npu_inst_pe_1_4_0_n115) );
  INV_X1 npu_inst_pe_1_4_0_U8 ( .A(npu_inst_pe_1_4_0_n42), .ZN(
        npu_inst_pe_1_4_0_n114) );
  BUF_X1 npu_inst_pe_1_4_0_U7 ( .A(npu_inst_pe_1_4_0_n11), .Z(
        npu_inst_pe_1_4_0_n10) );
  BUF_X1 npu_inst_pe_1_4_0_U6 ( .A(npu_inst_pe_1_4_0_n11), .Z(
        npu_inst_pe_1_4_0_n9) );
  BUF_X1 npu_inst_pe_1_4_0_U5 ( .A(npu_inst_pe_1_4_0_n11), .Z(
        npu_inst_pe_1_4_0_n8) );
  NOR2_X1 npu_inst_pe_1_4_0_U4 ( .A1(npu_inst_pe_1_4_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_0_n1), .ZN(npu_inst_pe_1_4_0_n76) );
  NOR2_X1 npu_inst_pe_1_4_0_U3 ( .A1(npu_inst_pe_1_4_0_n27), .A2(
        npu_inst_pe_1_4_0_n1), .ZN(npu_inst_pe_1_4_0_n77) );
  FA_X1 npu_inst_pe_1_4_0_sub_77_U2_1 ( .A(npu_inst_int_data_res_4__0__1_), 
        .B(npu_inst_pe_1_4_0_n13), .CI(npu_inst_pe_1_4_0_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_4_0_sub_77_carry_2_), .S(npu_inst_pe_1_4_0_N66) );
  FA_X1 npu_inst_pe_1_4_0_add_79_U1_1 ( .A(npu_inst_int_data_res_4__0__1_), 
        .B(npu_inst_pe_1_4_0_int_data_1_), .CI(
        npu_inst_pe_1_4_0_add_79_carry_1_), .CO(
        npu_inst_pe_1_4_0_add_79_carry_2_), .S(npu_inst_pe_1_4_0_N74) );
  NAND3_X1 npu_inst_pe_1_4_0_U101 ( .A1(npu_inst_pe_1_4_0_n4), .A2(
        npu_inst_pe_1_4_0_n6), .A3(npu_inst_pe_1_4_0_n7), .ZN(
        npu_inst_pe_1_4_0_n44) );
  NAND3_X1 npu_inst_pe_1_4_0_U100 ( .A1(npu_inst_pe_1_4_0_n3), .A2(
        npu_inst_pe_1_4_0_n6), .A3(npu_inst_pe_1_4_0_n7), .ZN(
        npu_inst_pe_1_4_0_n40) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_0_n33), .CK(
        npu_inst_pe_1_4_0_net3742), .RN(npu_inst_pe_1_4_0_n8), .Q(
        npu_inst_int_data_res_4__0__6_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_0_n34), .CK(
        npu_inst_pe_1_4_0_net3742), .RN(npu_inst_pe_1_4_0_n8), .Q(
        npu_inst_int_data_res_4__0__5_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_0_n35), .CK(
        npu_inst_pe_1_4_0_net3742), .RN(npu_inst_pe_1_4_0_n8), .Q(
        npu_inst_int_data_res_4__0__4_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_0_n36), .CK(
        npu_inst_pe_1_4_0_net3742), .RN(npu_inst_pe_1_4_0_n8), .Q(
        npu_inst_int_data_res_4__0__3_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_0_n98), .CK(
        npu_inst_pe_1_4_0_net3742), .RN(npu_inst_pe_1_4_0_n8), .Q(
        npu_inst_int_data_res_4__0__2_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_0_n99), .CK(
        npu_inst_pe_1_4_0_net3742), .RN(npu_inst_pe_1_4_0_n8), .Q(
        npu_inst_int_data_res_4__0__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_0_n32), .CK(
        npu_inst_pe_1_4_0_net3742), .RN(npu_inst_pe_1_4_0_n8), .Q(
        npu_inst_int_data_res_4__0__7_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_0_n100), 
        .CK(npu_inst_pe_1_4_0_net3742), .RN(npu_inst_pe_1_4_0_n8), .Q(
        npu_inst_int_data_res_4__0__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_weight_reg_0_ ( .D(npu_inst_n92), .CK(
        npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n8), .Q(
        npu_inst_pe_1_4_0_int_q_weight_0_), .QN(npu_inst_pe_1_4_0_n27) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_weight_reg_1_ ( .D(npu_inst_n98), .CK(
        npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n8), .Q(
        npu_inst_pe_1_4_0_int_q_weight_1_), .QN(npu_inst_pe_1_4_0_n26) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_0_n112), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n8), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_0_n106), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n8), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_0_n111), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_0_n105), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_0_n110), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_0_n104), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_0_n109), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_0_n103), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_0_n108), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_0_n102), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_0_n107), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_0_n101), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_0_n86), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_0_n87), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n9), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_0_n88), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_0_n89), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_0_n90), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_0_n91), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_0_n92), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_0_n93), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_0_n94), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_0_n95), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_0_n96), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_0_n97), 
        .CK(npu_inst_pe_1_4_0_net3748), .RN(npu_inst_pe_1_4_0_n10), .Q(
        npu_inst_pe_1_4_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_0_net3742) );
  CLKGATETST_X1 npu_inst_pe_1_4_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n45), .SE(1'b0), .GCK(npu_inst_pe_1_4_0_net3748) );
  MUX2_X1 npu_inst_pe_1_4_1_U153 ( .A(npu_inst_pe_1_4_1_n31), .B(
        npu_inst_pe_1_4_1_n28), .S(npu_inst_pe_1_4_1_n7), .Z(
        npu_inst_pe_1_4_1_N93) );
  MUX2_X1 npu_inst_pe_1_4_1_U152 ( .A(npu_inst_pe_1_4_1_n30), .B(
        npu_inst_pe_1_4_1_n29), .S(npu_inst_pe_1_4_1_n5), .Z(
        npu_inst_pe_1_4_1_n31) );
  MUX2_X1 npu_inst_pe_1_4_1_U151 ( .A(npu_inst_pe_1_4_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_1_n3), .Z(
        npu_inst_pe_1_4_1_n30) );
  MUX2_X1 npu_inst_pe_1_4_1_U150 ( .A(npu_inst_pe_1_4_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_1_n3), .Z(
        npu_inst_pe_1_4_1_n29) );
  MUX2_X1 npu_inst_pe_1_4_1_U149 ( .A(npu_inst_pe_1_4_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_1_n3), .Z(
        npu_inst_pe_1_4_1_n28) );
  MUX2_X1 npu_inst_pe_1_4_1_U148 ( .A(npu_inst_pe_1_4_1_n25), .B(
        npu_inst_pe_1_4_1_n22), .S(npu_inst_pe_1_4_1_n7), .Z(
        npu_inst_pe_1_4_1_N94) );
  MUX2_X1 npu_inst_pe_1_4_1_U147 ( .A(npu_inst_pe_1_4_1_n24), .B(
        npu_inst_pe_1_4_1_n23), .S(npu_inst_pe_1_4_1_n5), .Z(
        npu_inst_pe_1_4_1_n25) );
  MUX2_X1 npu_inst_pe_1_4_1_U146 ( .A(npu_inst_pe_1_4_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_1_n3), .Z(
        npu_inst_pe_1_4_1_n24) );
  MUX2_X1 npu_inst_pe_1_4_1_U145 ( .A(npu_inst_pe_1_4_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_1_n3), .Z(
        npu_inst_pe_1_4_1_n23) );
  MUX2_X1 npu_inst_pe_1_4_1_U144 ( .A(npu_inst_pe_1_4_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_1_n3), .Z(
        npu_inst_pe_1_4_1_n22) );
  MUX2_X1 npu_inst_pe_1_4_1_U143 ( .A(npu_inst_pe_1_4_1_n21), .B(
        npu_inst_pe_1_4_1_n18), .S(npu_inst_pe_1_4_1_n7), .Z(
        npu_inst_int_data_x_4__1__1_) );
  MUX2_X1 npu_inst_pe_1_4_1_U142 ( .A(npu_inst_pe_1_4_1_n20), .B(
        npu_inst_pe_1_4_1_n19), .S(npu_inst_pe_1_4_1_n5), .Z(
        npu_inst_pe_1_4_1_n21) );
  MUX2_X1 npu_inst_pe_1_4_1_U141 ( .A(npu_inst_pe_1_4_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_1_n3), .Z(
        npu_inst_pe_1_4_1_n20) );
  MUX2_X1 npu_inst_pe_1_4_1_U140 ( .A(npu_inst_pe_1_4_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_1_n3), .Z(
        npu_inst_pe_1_4_1_n19) );
  MUX2_X1 npu_inst_pe_1_4_1_U139 ( .A(npu_inst_pe_1_4_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_1_n3), .Z(
        npu_inst_pe_1_4_1_n18) );
  MUX2_X1 npu_inst_pe_1_4_1_U138 ( .A(npu_inst_pe_1_4_1_n17), .B(
        npu_inst_pe_1_4_1_n14), .S(npu_inst_pe_1_4_1_n7), .Z(
        npu_inst_int_data_x_4__1__0_) );
  MUX2_X1 npu_inst_pe_1_4_1_U137 ( .A(npu_inst_pe_1_4_1_n16), .B(
        npu_inst_pe_1_4_1_n15), .S(npu_inst_pe_1_4_1_n5), .Z(
        npu_inst_pe_1_4_1_n17) );
  MUX2_X1 npu_inst_pe_1_4_1_U136 ( .A(npu_inst_pe_1_4_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_1_n3), .Z(
        npu_inst_pe_1_4_1_n16) );
  MUX2_X1 npu_inst_pe_1_4_1_U135 ( .A(npu_inst_pe_1_4_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_1_n3), .Z(
        npu_inst_pe_1_4_1_n15) );
  MUX2_X1 npu_inst_pe_1_4_1_U134 ( .A(npu_inst_pe_1_4_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_1_n3), .Z(
        npu_inst_pe_1_4_1_n14) );
  XOR2_X1 npu_inst_pe_1_4_1_U133 ( .A(npu_inst_pe_1_4_1_int_data_0_), .B(
        npu_inst_int_data_res_4__1__0_), .Z(npu_inst_pe_1_4_1_N73) );
  AND2_X1 npu_inst_pe_1_4_1_U132 ( .A1(npu_inst_int_data_res_4__1__0_), .A2(
        npu_inst_pe_1_4_1_int_data_0_), .ZN(npu_inst_pe_1_4_1_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_1_U131 ( .A(npu_inst_int_data_res_4__1__0_), .B(
        npu_inst_pe_1_4_1_n12), .ZN(npu_inst_pe_1_4_1_N65) );
  OR2_X1 npu_inst_pe_1_4_1_U130 ( .A1(npu_inst_pe_1_4_1_n12), .A2(
        npu_inst_int_data_res_4__1__0_), .ZN(npu_inst_pe_1_4_1_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_1_U129 ( .A(npu_inst_int_data_res_4__1__2_), .B(
        npu_inst_pe_1_4_1_add_79_carry_2_), .Z(npu_inst_pe_1_4_1_N75) );
  AND2_X1 npu_inst_pe_1_4_1_U128 ( .A1(npu_inst_pe_1_4_1_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_4__1__2_), .ZN(
        npu_inst_pe_1_4_1_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_1_U127 ( .A(npu_inst_int_data_res_4__1__3_), .B(
        npu_inst_pe_1_4_1_add_79_carry_3_), .Z(npu_inst_pe_1_4_1_N76) );
  AND2_X1 npu_inst_pe_1_4_1_U126 ( .A1(npu_inst_pe_1_4_1_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_4__1__3_), .ZN(
        npu_inst_pe_1_4_1_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_1_U125 ( .A(npu_inst_int_data_res_4__1__4_), .B(
        npu_inst_pe_1_4_1_add_79_carry_4_), .Z(npu_inst_pe_1_4_1_N77) );
  AND2_X1 npu_inst_pe_1_4_1_U124 ( .A1(npu_inst_pe_1_4_1_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_4__1__4_), .ZN(
        npu_inst_pe_1_4_1_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_1_U123 ( .A(npu_inst_int_data_res_4__1__5_), .B(
        npu_inst_pe_1_4_1_add_79_carry_5_), .Z(npu_inst_pe_1_4_1_N78) );
  AND2_X1 npu_inst_pe_1_4_1_U122 ( .A1(npu_inst_pe_1_4_1_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_4__1__5_), .ZN(
        npu_inst_pe_1_4_1_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_1_U121 ( .A(npu_inst_int_data_res_4__1__6_), .B(
        npu_inst_pe_1_4_1_add_79_carry_6_), .Z(npu_inst_pe_1_4_1_N79) );
  AND2_X1 npu_inst_pe_1_4_1_U120 ( .A1(npu_inst_pe_1_4_1_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_4__1__6_), .ZN(
        npu_inst_pe_1_4_1_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_1_U119 ( .A(npu_inst_int_data_res_4__1__7_), .B(
        npu_inst_pe_1_4_1_add_79_carry_7_), .Z(npu_inst_pe_1_4_1_N80) );
  XNOR2_X1 npu_inst_pe_1_4_1_U118 ( .A(npu_inst_pe_1_4_1_sub_77_carry_2_), .B(
        npu_inst_int_data_res_4__1__2_), .ZN(npu_inst_pe_1_4_1_N67) );
  OR2_X1 npu_inst_pe_1_4_1_U117 ( .A1(npu_inst_int_data_res_4__1__2_), .A2(
        npu_inst_pe_1_4_1_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_4_1_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_1_U116 ( .A(npu_inst_pe_1_4_1_sub_77_carry_3_), .B(
        npu_inst_int_data_res_4__1__3_), .ZN(npu_inst_pe_1_4_1_N68) );
  OR2_X1 npu_inst_pe_1_4_1_U115 ( .A1(npu_inst_int_data_res_4__1__3_), .A2(
        npu_inst_pe_1_4_1_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_4_1_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_1_U114 ( .A(npu_inst_pe_1_4_1_sub_77_carry_4_), .B(
        npu_inst_int_data_res_4__1__4_), .ZN(npu_inst_pe_1_4_1_N69) );
  OR2_X1 npu_inst_pe_1_4_1_U113 ( .A1(npu_inst_int_data_res_4__1__4_), .A2(
        npu_inst_pe_1_4_1_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_4_1_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_1_U112 ( .A(npu_inst_pe_1_4_1_sub_77_carry_5_), .B(
        npu_inst_int_data_res_4__1__5_), .ZN(npu_inst_pe_1_4_1_N70) );
  OR2_X1 npu_inst_pe_1_4_1_U111 ( .A1(npu_inst_int_data_res_4__1__5_), .A2(
        npu_inst_pe_1_4_1_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_4_1_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_1_U110 ( .A(npu_inst_pe_1_4_1_sub_77_carry_6_), .B(
        npu_inst_int_data_res_4__1__6_), .ZN(npu_inst_pe_1_4_1_N71) );
  OR2_X1 npu_inst_pe_1_4_1_U109 ( .A1(npu_inst_int_data_res_4__1__6_), .A2(
        npu_inst_pe_1_4_1_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_4_1_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_1_U108 ( .A(npu_inst_int_data_res_4__1__7_), .B(
        npu_inst_pe_1_4_1_sub_77_carry_7_), .ZN(npu_inst_pe_1_4_1_N72) );
  INV_X1 npu_inst_pe_1_4_1_U107 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_4_1_n6)
         );
  INV_X1 npu_inst_pe_1_4_1_U106 ( .A(npu_inst_pe_1_4_1_n6), .ZN(
        npu_inst_pe_1_4_1_n5) );
  INV_X1 npu_inst_pe_1_4_1_U105 ( .A(npu_inst_n38), .ZN(npu_inst_pe_1_4_1_n2)
         );
  AOI22_X1 npu_inst_pe_1_4_1_U104 ( .A1(npu_inst_int_data_y_5__1__0_), .A2(
        npu_inst_pe_1_4_1_n58), .B1(npu_inst_pe_1_4_1_n118), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_1_n57) );
  INV_X1 npu_inst_pe_1_4_1_U103 ( .A(npu_inst_pe_1_4_1_n57), .ZN(
        npu_inst_pe_1_4_1_n107) );
  AOI22_X1 npu_inst_pe_1_4_1_U102 ( .A1(npu_inst_int_data_y_5__1__0_), .A2(
        npu_inst_pe_1_4_1_n54), .B1(npu_inst_pe_1_4_1_n117), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_1_n53) );
  INV_X1 npu_inst_pe_1_4_1_U99 ( .A(npu_inst_pe_1_4_1_n53), .ZN(
        npu_inst_pe_1_4_1_n108) );
  AOI22_X1 npu_inst_pe_1_4_1_U98 ( .A1(npu_inst_int_data_y_5__1__0_), .A2(
        npu_inst_pe_1_4_1_n50), .B1(npu_inst_pe_1_4_1_n116), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_1_n49) );
  INV_X1 npu_inst_pe_1_4_1_U97 ( .A(npu_inst_pe_1_4_1_n49), .ZN(
        npu_inst_pe_1_4_1_n109) );
  AOI22_X1 npu_inst_pe_1_4_1_U96 ( .A1(npu_inst_int_data_y_5__1__0_), .A2(
        npu_inst_pe_1_4_1_n46), .B1(npu_inst_pe_1_4_1_n115), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_1_n45) );
  INV_X1 npu_inst_pe_1_4_1_U95 ( .A(npu_inst_pe_1_4_1_n45), .ZN(
        npu_inst_pe_1_4_1_n110) );
  AOI22_X1 npu_inst_pe_1_4_1_U94 ( .A1(npu_inst_int_data_y_5__1__0_), .A2(
        npu_inst_pe_1_4_1_n42), .B1(npu_inst_pe_1_4_1_n114), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_1_n41) );
  INV_X1 npu_inst_pe_1_4_1_U93 ( .A(npu_inst_pe_1_4_1_n41), .ZN(
        npu_inst_pe_1_4_1_n111) );
  AOI22_X1 npu_inst_pe_1_4_1_U92 ( .A1(npu_inst_int_data_y_5__1__1_), .A2(
        npu_inst_pe_1_4_1_n58), .B1(npu_inst_pe_1_4_1_n118), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_1_n59) );
  INV_X1 npu_inst_pe_1_4_1_U91 ( .A(npu_inst_pe_1_4_1_n59), .ZN(
        npu_inst_pe_1_4_1_n101) );
  AOI22_X1 npu_inst_pe_1_4_1_U90 ( .A1(npu_inst_int_data_y_5__1__1_), .A2(
        npu_inst_pe_1_4_1_n54), .B1(npu_inst_pe_1_4_1_n117), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_1_n55) );
  INV_X1 npu_inst_pe_1_4_1_U89 ( .A(npu_inst_pe_1_4_1_n55), .ZN(
        npu_inst_pe_1_4_1_n102) );
  AOI22_X1 npu_inst_pe_1_4_1_U88 ( .A1(npu_inst_int_data_y_5__1__1_), .A2(
        npu_inst_pe_1_4_1_n50), .B1(npu_inst_pe_1_4_1_n116), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_1_n51) );
  INV_X1 npu_inst_pe_1_4_1_U87 ( .A(npu_inst_pe_1_4_1_n51), .ZN(
        npu_inst_pe_1_4_1_n103) );
  AOI22_X1 npu_inst_pe_1_4_1_U86 ( .A1(npu_inst_int_data_y_5__1__1_), .A2(
        npu_inst_pe_1_4_1_n46), .B1(npu_inst_pe_1_4_1_n115), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_1_n47) );
  INV_X1 npu_inst_pe_1_4_1_U85 ( .A(npu_inst_pe_1_4_1_n47), .ZN(
        npu_inst_pe_1_4_1_n104) );
  AOI22_X1 npu_inst_pe_1_4_1_U84 ( .A1(npu_inst_int_data_y_5__1__1_), .A2(
        npu_inst_pe_1_4_1_n42), .B1(npu_inst_pe_1_4_1_n114), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_1_n43) );
  INV_X1 npu_inst_pe_1_4_1_U83 ( .A(npu_inst_pe_1_4_1_n43), .ZN(
        npu_inst_pe_1_4_1_n105) );
  AOI22_X1 npu_inst_pe_1_4_1_U82 ( .A1(npu_inst_pe_1_4_1_n38), .A2(
        npu_inst_int_data_y_5__1__1_), .B1(npu_inst_pe_1_4_1_n113), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_1_n39) );
  INV_X1 npu_inst_pe_1_4_1_U81 ( .A(npu_inst_pe_1_4_1_n39), .ZN(
        npu_inst_pe_1_4_1_n106) );
  AND2_X1 npu_inst_pe_1_4_1_U80 ( .A1(npu_inst_pe_1_4_1_N93), .A2(npu_inst_n38), .ZN(npu_inst_int_data_y_4__1__0_) );
  NAND2_X1 npu_inst_pe_1_4_1_U79 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_1_n60), .ZN(npu_inst_pe_1_4_1_n74) );
  OAI21_X1 npu_inst_pe_1_4_1_U78 ( .B1(npu_inst_pe_1_4_1_n63), .B2(
        npu_inst_pe_1_4_1_n60), .A(npu_inst_pe_1_4_1_n74), .ZN(
        npu_inst_pe_1_4_1_n97) );
  NAND2_X1 npu_inst_pe_1_4_1_U77 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_1_n60), .ZN(npu_inst_pe_1_4_1_n73) );
  OAI21_X1 npu_inst_pe_1_4_1_U76 ( .B1(npu_inst_pe_1_4_1_n61), .B2(
        npu_inst_pe_1_4_1_n60), .A(npu_inst_pe_1_4_1_n73), .ZN(
        npu_inst_pe_1_4_1_n96) );
  NAND2_X1 npu_inst_pe_1_4_1_U75 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_1_n56), .ZN(npu_inst_pe_1_4_1_n72) );
  OAI21_X1 npu_inst_pe_1_4_1_U74 ( .B1(npu_inst_pe_1_4_1_n63), .B2(
        npu_inst_pe_1_4_1_n56), .A(npu_inst_pe_1_4_1_n72), .ZN(
        npu_inst_pe_1_4_1_n95) );
  NAND2_X1 npu_inst_pe_1_4_1_U73 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_1_n56), .ZN(npu_inst_pe_1_4_1_n71) );
  OAI21_X1 npu_inst_pe_1_4_1_U72 ( .B1(npu_inst_pe_1_4_1_n61), .B2(
        npu_inst_pe_1_4_1_n56), .A(npu_inst_pe_1_4_1_n71), .ZN(
        npu_inst_pe_1_4_1_n94) );
  NAND2_X1 npu_inst_pe_1_4_1_U71 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_1_n52), .ZN(npu_inst_pe_1_4_1_n70) );
  OAI21_X1 npu_inst_pe_1_4_1_U70 ( .B1(npu_inst_pe_1_4_1_n63), .B2(
        npu_inst_pe_1_4_1_n52), .A(npu_inst_pe_1_4_1_n70), .ZN(
        npu_inst_pe_1_4_1_n93) );
  NAND2_X1 npu_inst_pe_1_4_1_U69 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_1_n52), .ZN(npu_inst_pe_1_4_1_n69) );
  OAI21_X1 npu_inst_pe_1_4_1_U68 ( .B1(npu_inst_pe_1_4_1_n61), .B2(
        npu_inst_pe_1_4_1_n52), .A(npu_inst_pe_1_4_1_n69), .ZN(
        npu_inst_pe_1_4_1_n92) );
  NAND2_X1 npu_inst_pe_1_4_1_U67 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_1_n48), .ZN(npu_inst_pe_1_4_1_n68) );
  OAI21_X1 npu_inst_pe_1_4_1_U66 ( .B1(npu_inst_pe_1_4_1_n63), .B2(
        npu_inst_pe_1_4_1_n48), .A(npu_inst_pe_1_4_1_n68), .ZN(
        npu_inst_pe_1_4_1_n91) );
  NAND2_X1 npu_inst_pe_1_4_1_U65 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_1_n48), .ZN(npu_inst_pe_1_4_1_n67) );
  OAI21_X1 npu_inst_pe_1_4_1_U64 ( .B1(npu_inst_pe_1_4_1_n61), .B2(
        npu_inst_pe_1_4_1_n48), .A(npu_inst_pe_1_4_1_n67), .ZN(
        npu_inst_pe_1_4_1_n90) );
  NAND2_X1 npu_inst_pe_1_4_1_U63 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_1_n44), .ZN(npu_inst_pe_1_4_1_n66) );
  OAI21_X1 npu_inst_pe_1_4_1_U62 ( .B1(npu_inst_pe_1_4_1_n63), .B2(
        npu_inst_pe_1_4_1_n44), .A(npu_inst_pe_1_4_1_n66), .ZN(
        npu_inst_pe_1_4_1_n89) );
  NAND2_X1 npu_inst_pe_1_4_1_U61 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_1_n44), .ZN(npu_inst_pe_1_4_1_n65) );
  OAI21_X1 npu_inst_pe_1_4_1_U60 ( .B1(npu_inst_pe_1_4_1_n61), .B2(
        npu_inst_pe_1_4_1_n44), .A(npu_inst_pe_1_4_1_n65), .ZN(
        npu_inst_pe_1_4_1_n88) );
  NAND2_X1 npu_inst_pe_1_4_1_U59 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_1_n40), .ZN(npu_inst_pe_1_4_1_n64) );
  OAI21_X1 npu_inst_pe_1_4_1_U58 ( .B1(npu_inst_pe_1_4_1_n63), .B2(
        npu_inst_pe_1_4_1_n40), .A(npu_inst_pe_1_4_1_n64), .ZN(
        npu_inst_pe_1_4_1_n87) );
  NAND2_X1 npu_inst_pe_1_4_1_U57 ( .A1(npu_inst_pe_1_4_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_1_n40), .ZN(npu_inst_pe_1_4_1_n62) );
  OAI21_X1 npu_inst_pe_1_4_1_U56 ( .B1(npu_inst_pe_1_4_1_n61), .B2(
        npu_inst_pe_1_4_1_n40), .A(npu_inst_pe_1_4_1_n62), .ZN(
        npu_inst_pe_1_4_1_n86) );
  AOI22_X1 npu_inst_pe_1_4_1_U55 ( .A1(npu_inst_pe_1_4_1_n38), .A2(
        npu_inst_int_data_y_5__1__0_), .B1(npu_inst_pe_1_4_1_n113), .B2(
        npu_inst_pe_1_4_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_1_n37) );
  INV_X1 npu_inst_pe_1_4_1_U54 ( .A(npu_inst_pe_1_4_1_n37), .ZN(
        npu_inst_pe_1_4_1_n112) );
  AND2_X1 npu_inst_pe_1_4_1_U53 ( .A1(npu_inst_n38), .A2(npu_inst_pe_1_4_1_N94), .ZN(npu_inst_int_data_y_4__1__1_) );
  AOI222_X1 npu_inst_pe_1_4_1_U52 ( .A1(npu_inst_int_data_res_5__1__0_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N73), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N65), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n84) );
  INV_X1 npu_inst_pe_1_4_1_U51 ( .A(npu_inst_pe_1_4_1_n84), .ZN(
        npu_inst_pe_1_4_1_n100) );
  AOI222_X1 npu_inst_pe_1_4_1_U50 ( .A1(npu_inst_pe_1_4_1_n1), .A2(
        npu_inst_int_data_res_5__1__7_), .B1(npu_inst_pe_1_4_1_N80), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N72), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n75) );
  INV_X1 npu_inst_pe_1_4_1_U49 ( .A(npu_inst_pe_1_4_1_n75), .ZN(
        npu_inst_pe_1_4_1_n32) );
  AOI222_X1 npu_inst_pe_1_4_1_U48 ( .A1(npu_inst_int_data_res_5__1__1_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N74), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N66), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n83) );
  INV_X1 npu_inst_pe_1_4_1_U47 ( .A(npu_inst_pe_1_4_1_n83), .ZN(
        npu_inst_pe_1_4_1_n99) );
  AOI222_X1 npu_inst_pe_1_4_1_U46 ( .A1(npu_inst_int_data_res_5__1__3_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N76), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N68), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n81) );
  INV_X1 npu_inst_pe_1_4_1_U45 ( .A(npu_inst_pe_1_4_1_n81), .ZN(
        npu_inst_pe_1_4_1_n36) );
  AOI222_X1 npu_inst_pe_1_4_1_U44 ( .A1(npu_inst_int_data_res_5__1__4_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N77), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N69), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n80) );
  INV_X1 npu_inst_pe_1_4_1_U43 ( .A(npu_inst_pe_1_4_1_n80), .ZN(
        npu_inst_pe_1_4_1_n35) );
  AOI222_X1 npu_inst_pe_1_4_1_U42 ( .A1(npu_inst_int_data_res_5__1__5_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N78), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N70), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n79) );
  INV_X1 npu_inst_pe_1_4_1_U41 ( .A(npu_inst_pe_1_4_1_n79), .ZN(
        npu_inst_pe_1_4_1_n34) );
  AOI222_X1 npu_inst_pe_1_4_1_U40 ( .A1(npu_inst_int_data_res_5__1__6_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N79), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N71), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n78) );
  INV_X1 npu_inst_pe_1_4_1_U39 ( .A(npu_inst_pe_1_4_1_n78), .ZN(
        npu_inst_pe_1_4_1_n33) );
  AND2_X1 npu_inst_pe_1_4_1_U38 ( .A1(npu_inst_int_data_x_4__1__1_), .A2(
        npu_inst_pe_1_4_1_int_q_weight_1_), .ZN(npu_inst_pe_1_4_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_1_U37 ( .A1(npu_inst_int_data_x_4__1__0_), .A2(
        npu_inst_pe_1_4_1_int_q_weight_1_), .ZN(npu_inst_pe_1_4_1_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_4_1_U36 ( .A(npu_inst_pe_1_4_1_int_data_1_), .ZN(
        npu_inst_pe_1_4_1_n13) );
  NOR3_X1 npu_inst_pe_1_4_1_U35 ( .A1(npu_inst_pe_1_4_1_n26), .A2(npu_inst_n38), .A3(npu_inst_int_ckg[30]), .ZN(npu_inst_pe_1_4_1_n85) );
  OR2_X1 npu_inst_pe_1_4_1_U34 ( .A1(npu_inst_pe_1_4_1_n85), .A2(
        npu_inst_pe_1_4_1_n1), .ZN(npu_inst_pe_1_4_1_N84) );
  AOI222_X1 npu_inst_pe_1_4_1_U33 ( .A1(npu_inst_int_data_res_5__1__2_), .A2(
        npu_inst_pe_1_4_1_n1), .B1(npu_inst_pe_1_4_1_N75), .B2(
        npu_inst_pe_1_4_1_n76), .C1(npu_inst_pe_1_4_1_N67), .C2(
        npu_inst_pe_1_4_1_n77), .ZN(npu_inst_pe_1_4_1_n82) );
  INV_X1 npu_inst_pe_1_4_1_U32 ( .A(npu_inst_pe_1_4_1_n82), .ZN(
        npu_inst_pe_1_4_1_n98) );
  AOI22_X1 npu_inst_pe_1_4_1_U31 ( .A1(npu_inst_n38), .A2(
        npu_inst_int_data_y_5__1__1_), .B1(npu_inst_pe_1_4_1_n2), .B2(
        npu_inst_int_data_x_4__2__1_), .ZN(npu_inst_pe_1_4_1_n63) );
  AOI22_X1 npu_inst_pe_1_4_1_U30 ( .A1(npu_inst_n38), .A2(
        npu_inst_int_data_y_5__1__0_), .B1(npu_inst_pe_1_4_1_n2), .B2(
        npu_inst_int_data_x_4__2__0_), .ZN(npu_inst_pe_1_4_1_n61) );
  INV_X1 npu_inst_pe_1_4_1_U29 ( .A(npu_inst_pe_1_4_1_int_data_0_), .ZN(
        npu_inst_pe_1_4_1_n12) );
  INV_X1 npu_inst_pe_1_4_1_U28 ( .A(npu_inst_n51), .ZN(npu_inst_pe_1_4_1_n4)
         );
  OR3_X1 npu_inst_pe_1_4_1_U27 ( .A1(npu_inst_pe_1_4_1_n5), .A2(
        npu_inst_pe_1_4_1_n7), .A3(npu_inst_pe_1_4_1_n4), .ZN(
        npu_inst_pe_1_4_1_n56) );
  OR3_X1 npu_inst_pe_1_4_1_U26 ( .A1(npu_inst_pe_1_4_1_n4), .A2(
        npu_inst_pe_1_4_1_n7), .A3(npu_inst_pe_1_4_1_n6), .ZN(
        npu_inst_pe_1_4_1_n48) );
  INV_X1 npu_inst_pe_1_4_1_U25 ( .A(npu_inst_pe_1_4_1_n4), .ZN(
        npu_inst_pe_1_4_1_n3) );
  OR3_X1 npu_inst_pe_1_4_1_U24 ( .A1(npu_inst_pe_1_4_1_n3), .A2(
        npu_inst_pe_1_4_1_n7), .A3(npu_inst_pe_1_4_1_n6), .ZN(
        npu_inst_pe_1_4_1_n52) );
  OR3_X1 npu_inst_pe_1_4_1_U23 ( .A1(npu_inst_pe_1_4_1_n5), .A2(
        npu_inst_pe_1_4_1_n7), .A3(npu_inst_pe_1_4_1_n3), .ZN(
        npu_inst_pe_1_4_1_n60) );
  BUF_X1 npu_inst_pe_1_4_1_U22 ( .A(npu_inst_n21), .Z(npu_inst_pe_1_4_1_n1) );
  NOR2_X1 npu_inst_pe_1_4_1_U21 ( .A1(npu_inst_pe_1_4_1_n60), .A2(
        npu_inst_pe_1_4_1_n2), .ZN(npu_inst_pe_1_4_1_n58) );
  NOR2_X1 npu_inst_pe_1_4_1_U20 ( .A1(npu_inst_pe_1_4_1_n56), .A2(
        npu_inst_pe_1_4_1_n2), .ZN(npu_inst_pe_1_4_1_n54) );
  NOR2_X1 npu_inst_pe_1_4_1_U19 ( .A1(npu_inst_pe_1_4_1_n52), .A2(
        npu_inst_pe_1_4_1_n2), .ZN(npu_inst_pe_1_4_1_n50) );
  NOR2_X1 npu_inst_pe_1_4_1_U18 ( .A1(npu_inst_pe_1_4_1_n48), .A2(
        npu_inst_pe_1_4_1_n2), .ZN(npu_inst_pe_1_4_1_n46) );
  NOR2_X1 npu_inst_pe_1_4_1_U17 ( .A1(npu_inst_pe_1_4_1_n40), .A2(
        npu_inst_pe_1_4_1_n2), .ZN(npu_inst_pe_1_4_1_n38) );
  NOR2_X1 npu_inst_pe_1_4_1_U16 ( .A1(npu_inst_pe_1_4_1_n44), .A2(
        npu_inst_pe_1_4_1_n2), .ZN(npu_inst_pe_1_4_1_n42) );
  BUF_X1 npu_inst_pe_1_4_1_U15 ( .A(npu_inst_n81), .Z(npu_inst_pe_1_4_1_n7) );
  INV_X1 npu_inst_pe_1_4_1_U14 ( .A(npu_inst_n106), .ZN(npu_inst_pe_1_4_1_n11)
         );
  INV_X1 npu_inst_pe_1_4_1_U13 ( .A(npu_inst_pe_1_4_1_n38), .ZN(
        npu_inst_pe_1_4_1_n113) );
  INV_X1 npu_inst_pe_1_4_1_U12 ( .A(npu_inst_pe_1_4_1_n58), .ZN(
        npu_inst_pe_1_4_1_n118) );
  INV_X1 npu_inst_pe_1_4_1_U11 ( .A(npu_inst_pe_1_4_1_n54), .ZN(
        npu_inst_pe_1_4_1_n117) );
  INV_X1 npu_inst_pe_1_4_1_U10 ( .A(npu_inst_pe_1_4_1_n50), .ZN(
        npu_inst_pe_1_4_1_n116) );
  INV_X1 npu_inst_pe_1_4_1_U9 ( .A(npu_inst_pe_1_4_1_n46), .ZN(
        npu_inst_pe_1_4_1_n115) );
  INV_X1 npu_inst_pe_1_4_1_U8 ( .A(npu_inst_pe_1_4_1_n42), .ZN(
        npu_inst_pe_1_4_1_n114) );
  BUF_X1 npu_inst_pe_1_4_1_U7 ( .A(npu_inst_pe_1_4_1_n11), .Z(
        npu_inst_pe_1_4_1_n10) );
  BUF_X1 npu_inst_pe_1_4_1_U6 ( .A(npu_inst_pe_1_4_1_n11), .Z(
        npu_inst_pe_1_4_1_n9) );
  BUF_X1 npu_inst_pe_1_4_1_U5 ( .A(npu_inst_pe_1_4_1_n11), .Z(
        npu_inst_pe_1_4_1_n8) );
  NOR2_X1 npu_inst_pe_1_4_1_U4 ( .A1(npu_inst_pe_1_4_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_1_n1), .ZN(npu_inst_pe_1_4_1_n76) );
  NOR2_X1 npu_inst_pe_1_4_1_U3 ( .A1(npu_inst_pe_1_4_1_n27), .A2(
        npu_inst_pe_1_4_1_n1), .ZN(npu_inst_pe_1_4_1_n77) );
  FA_X1 npu_inst_pe_1_4_1_sub_77_U2_1 ( .A(npu_inst_int_data_res_4__1__1_), 
        .B(npu_inst_pe_1_4_1_n13), .CI(npu_inst_pe_1_4_1_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_4_1_sub_77_carry_2_), .S(npu_inst_pe_1_4_1_N66) );
  FA_X1 npu_inst_pe_1_4_1_add_79_U1_1 ( .A(npu_inst_int_data_res_4__1__1_), 
        .B(npu_inst_pe_1_4_1_int_data_1_), .CI(
        npu_inst_pe_1_4_1_add_79_carry_1_), .CO(
        npu_inst_pe_1_4_1_add_79_carry_2_), .S(npu_inst_pe_1_4_1_N74) );
  NAND3_X1 npu_inst_pe_1_4_1_U101 ( .A1(npu_inst_pe_1_4_1_n4), .A2(
        npu_inst_pe_1_4_1_n6), .A3(npu_inst_pe_1_4_1_n7), .ZN(
        npu_inst_pe_1_4_1_n44) );
  NAND3_X1 npu_inst_pe_1_4_1_U100 ( .A1(npu_inst_pe_1_4_1_n3), .A2(
        npu_inst_pe_1_4_1_n6), .A3(npu_inst_pe_1_4_1_n7), .ZN(
        npu_inst_pe_1_4_1_n40) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_1_n33), .CK(
        npu_inst_pe_1_4_1_net3719), .RN(npu_inst_pe_1_4_1_n8), .Q(
        npu_inst_int_data_res_4__1__6_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_1_n34), .CK(
        npu_inst_pe_1_4_1_net3719), .RN(npu_inst_pe_1_4_1_n8), .Q(
        npu_inst_int_data_res_4__1__5_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_1_n35), .CK(
        npu_inst_pe_1_4_1_net3719), .RN(npu_inst_pe_1_4_1_n8), .Q(
        npu_inst_int_data_res_4__1__4_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_1_n36), .CK(
        npu_inst_pe_1_4_1_net3719), .RN(npu_inst_pe_1_4_1_n8), .Q(
        npu_inst_int_data_res_4__1__3_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_1_n98), .CK(
        npu_inst_pe_1_4_1_net3719), .RN(npu_inst_pe_1_4_1_n8), .Q(
        npu_inst_int_data_res_4__1__2_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_1_n99), .CK(
        npu_inst_pe_1_4_1_net3719), .RN(npu_inst_pe_1_4_1_n8), .Q(
        npu_inst_int_data_res_4__1__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_1_n32), .CK(
        npu_inst_pe_1_4_1_net3719), .RN(npu_inst_pe_1_4_1_n8), .Q(
        npu_inst_int_data_res_4__1__7_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_1_n100), 
        .CK(npu_inst_pe_1_4_1_net3719), .RN(npu_inst_pe_1_4_1_n8), .Q(
        npu_inst_int_data_res_4__1__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_weight_reg_0_ ( .D(npu_inst_n92), .CK(
        npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n8), .Q(
        npu_inst_pe_1_4_1_int_q_weight_0_), .QN(npu_inst_pe_1_4_1_n27) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_weight_reg_1_ ( .D(npu_inst_n98), .CK(
        npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n8), .Q(
        npu_inst_pe_1_4_1_int_q_weight_1_), .QN(npu_inst_pe_1_4_1_n26) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_1_n112), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n8), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_1_n106), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n8), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_1_n111), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_1_n105), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_1_n110), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_1_n104), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_1_n109), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_1_n103), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_1_n108), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_1_n102), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_1_n107), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_1_n101), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_1_n86), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_1_n87), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n9), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_1_n88), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_1_n89), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_1_n90), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_1_n91), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_1_n92), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_1_n93), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_1_n94), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_1_n95), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_1_n96), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_1_n97), 
        .CK(npu_inst_pe_1_4_1_net3725), .RN(npu_inst_pe_1_4_1_n10), .Q(
        npu_inst_pe_1_4_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_1_net3719) );
  CLKGATETST_X1 npu_inst_pe_1_4_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n45), .SE(1'b0), .GCK(npu_inst_pe_1_4_1_net3725) );
  MUX2_X1 npu_inst_pe_1_4_2_U153 ( .A(npu_inst_pe_1_4_2_n31), .B(
        npu_inst_pe_1_4_2_n28), .S(npu_inst_pe_1_4_2_n7), .Z(
        npu_inst_pe_1_4_2_N93) );
  MUX2_X1 npu_inst_pe_1_4_2_U152 ( .A(npu_inst_pe_1_4_2_n30), .B(
        npu_inst_pe_1_4_2_n29), .S(npu_inst_pe_1_4_2_n5), .Z(
        npu_inst_pe_1_4_2_n31) );
  MUX2_X1 npu_inst_pe_1_4_2_U151 ( .A(npu_inst_pe_1_4_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_2_n3), .Z(
        npu_inst_pe_1_4_2_n30) );
  MUX2_X1 npu_inst_pe_1_4_2_U150 ( .A(npu_inst_pe_1_4_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_2_n3), .Z(
        npu_inst_pe_1_4_2_n29) );
  MUX2_X1 npu_inst_pe_1_4_2_U149 ( .A(npu_inst_pe_1_4_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_2_n3), .Z(
        npu_inst_pe_1_4_2_n28) );
  MUX2_X1 npu_inst_pe_1_4_2_U148 ( .A(npu_inst_pe_1_4_2_n25), .B(
        npu_inst_pe_1_4_2_n22), .S(npu_inst_pe_1_4_2_n7), .Z(
        npu_inst_pe_1_4_2_N94) );
  MUX2_X1 npu_inst_pe_1_4_2_U147 ( .A(npu_inst_pe_1_4_2_n24), .B(
        npu_inst_pe_1_4_2_n23), .S(npu_inst_pe_1_4_2_n5), .Z(
        npu_inst_pe_1_4_2_n25) );
  MUX2_X1 npu_inst_pe_1_4_2_U146 ( .A(npu_inst_pe_1_4_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_2_n3), .Z(
        npu_inst_pe_1_4_2_n24) );
  MUX2_X1 npu_inst_pe_1_4_2_U145 ( .A(npu_inst_pe_1_4_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_2_n3), .Z(
        npu_inst_pe_1_4_2_n23) );
  MUX2_X1 npu_inst_pe_1_4_2_U144 ( .A(npu_inst_pe_1_4_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_2_n3), .Z(
        npu_inst_pe_1_4_2_n22) );
  MUX2_X1 npu_inst_pe_1_4_2_U143 ( .A(npu_inst_pe_1_4_2_n21), .B(
        npu_inst_pe_1_4_2_n18), .S(npu_inst_pe_1_4_2_n7), .Z(
        npu_inst_int_data_x_4__2__1_) );
  MUX2_X1 npu_inst_pe_1_4_2_U142 ( .A(npu_inst_pe_1_4_2_n20), .B(
        npu_inst_pe_1_4_2_n19), .S(npu_inst_pe_1_4_2_n5), .Z(
        npu_inst_pe_1_4_2_n21) );
  MUX2_X1 npu_inst_pe_1_4_2_U141 ( .A(npu_inst_pe_1_4_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_2_n3), .Z(
        npu_inst_pe_1_4_2_n20) );
  MUX2_X1 npu_inst_pe_1_4_2_U140 ( .A(npu_inst_pe_1_4_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_2_n3), .Z(
        npu_inst_pe_1_4_2_n19) );
  MUX2_X1 npu_inst_pe_1_4_2_U139 ( .A(npu_inst_pe_1_4_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_2_n3), .Z(
        npu_inst_pe_1_4_2_n18) );
  MUX2_X1 npu_inst_pe_1_4_2_U138 ( .A(npu_inst_pe_1_4_2_n17), .B(
        npu_inst_pe_1_4_2_n14), .S(npu_inst_pe_1_4_2_n7), .Z(
        npu_inst_int_data_x_4__2__0_) );
  MUX2_X1 npu_inst_pe_1_4_2_U137 ( .A(npu_inst_pe_1_4_2_n16), .B(
        npu_inst_pe_1_4_2_n15), .S(npu_inst_pe_1_4_2_n5), .Z(
        npu_inst_pe_1_4_2_n17) );
  MUX2_X1 npu_inst_pe_1_4_2_U136 ( .A(npu_inst_pe_1_4_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_2_n3), .Z(
        npu_inst_pe_1_4_2_n16) );
  MUX2_X1 npu_inst_pe_1_4_2_U135 ( .A(npu_inst_pe_1_4_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_2_n3), .Z(
        npu_inst_pe_1_4_2_n15) );
  MUX2_X1 npu_inst_pe_1_4_2_U134 ( .A(npu_inst_pe_1_4_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_2_n3), .Z(
        npu_inst_pe_1_4_2_n14) );
  XOR2_X1 npu_inst_pe_1_4_2_U133 ( .A(npu_inst_pe_1_4_2_int_data_0_), .B(
        npu_inst_int_data_res_4__2__0_), .Z(npu_inst_pe_1_4_2_N73) );
  AND2_X1 npu_inst_pe_1_4_2_U132 ( .A1(npu_inst_int_data_res_4__2__0_), .A2(
        npu_inst_pe_1_4_2_int_data_0_), .ZN(npu_inst_pe_1_4_2_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_2_U131 ( .A(npu_inst_int_data_res_4__2__0_), .B(
        npu_inst_pe_1_4_2_n12), .ZN(npu_inst_pe_1_4_2_N65) );
  OR2_X1 npu_inst_pe_1_4_2_U130 ( .A1(npu_inst_pe_1_4_2_n12), .A2(
        npu_inst_int_data_res_4__2__0_), .ZN(npu_inst_pe_1_4_2_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_2_U129 ( .A(npu_inst_int_data_res_4__2__2_), .B(
        npu_inst_pe_1_4_2_add_79_carry_2_), .Z(npu_inst_pe_1_4_2_N75) );
  AND2_X1 npu_inst_pe_1_4_2_U128 ( .A1(npu_inst_pe_1_4_2_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_4__2__2_), .ZN(
        npu_inst_pe_1_4_2_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_2_U127 ( .A(npu_inst_int_data_res_4__2__3_), .B(
        npu_inst_pe_1_4_2_add_79_carry_3_), .Z(npu_inst_pe_1_4_2_N76) );
  AND2_X1 npu_inst_pe_1_4_2_U126 ( .A1(npu_inst_pe_1_4_2_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_4__2__3_), .ZN(
        npu_inst_pe_1_4_2_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_2_U125 ( .A(npu_inst_int_data_res_4__2__4_), .B(
        npu_inst_pe_1_4_2_add_79_carry_4_), .Z(npu_inst_pe_1_4_2_N77) );
  AND2_X1 npu_inst_pe_1_4_2_U124 ( .A1(npu_inst_pe_1_4_2_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_4__2__4_), .ZN(
        npu_inst_pe_1_4_2_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_2_U123 ( .A(npu_inst_int_data_res_4__2__5_), .B(
        npu_inst_pe_1_4_2_add_79_carry_5_), .Z(npu_inst_pe_1_4_2_N78) );
  AND2_X1 npu_inst_pe_1_4_2_U122 ( .A1(npu_inst_pe_1_4_2_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_4__2__5_), .ZN(
        npu_inst_pe_1_4_2_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_2_U121 ( .A(npu_inst_int_data_res_4__2__6_), .B(
        npu_inst_pe_1_4_2_add_79_carry_6_), .Z(npu_inst_pe_1_4_2_N79) );
  AND2_X1 npu_inst_pe_1_4_2_U120 ( .A1(npu_inst_pe_1_4_2_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_4__2__6_), .ZN(
        npu_inst_pe_1_4_2_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_2_U119 ( .A(npu_inst_int_data_res_4__2__7_), .B(
        npu_inst_pe_1_4_2_add_79_carry_7_), .Z(npu_inst_pe_1_4_2_N80) );
  XNOR2_X1 npu_inst_pe_1_4_2_U118 ( .A(npu_inst_pe_1_4_2_sub_77_carry_2_), .B(
        npu_inst_int_data_res_4__2__2_), .ZN(npu_inst_pe_1_4_2_N67) );
  OR2_X1 npu_inst_pe_1_4_2_U117 ( .A1(npu_inst_int_data_res_4__2__2_), .A2(
        npu_inst_pe_1_4_2_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_4_2_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_2_U116 ( .A(npu_inst_pe_1_4_2_sub_77_carry_3_), .B(
        npu_inst_int_data_res_4__2__3_), .ZN(npu_inst_pe_1_4_2_N68) );
  OR2_X1 npu_inst_pe_1_4_2_U115 ( .A1(npu_inst_int_data_res_4__2__3_), .A2(
        npu_inst_pe_1_4_2_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_4_2_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_2_U114 ( .A(npu_inst_pe_1_4_2_sub_77_carry_4_), .B(
        npu_inst_int_data_res_4__2__4_), .ZN(npu_inst_pe_1_4_2_N69) );
  OR2_X1 npu_inst_pe_1_4_2_U113 ( .A1(npu_inst_int_data_res_4__2__4_), .A2(
        npu_inst_pe_1_4_2_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_4_2_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_2_U112 ( .A(npu_inst_pe_1_4_2_sub_77_carry_5_), .B(
        npu_inst_int_data_res_4__2__5_), .ZN(npu_inst_pe_1_4_2_N70) );
  OR2_X1 npu_inst_pe_1_4_2_U111 ( .A1(npu_inst_int_data_res_4__2__5_), .A2(
        npu_inst_pe_1_4_2_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_4_2_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_2_U110 ( .A(npu_inst_pe_1_4_2_sub_77_carry_6_), .B(
        npu_inst_int_data_res_4__2__6_), .ZN(npu_inst_pe_1_4_2_N71) );
  OR2_X1 npu_inst_pe_1_4_2_U109 ( .A1(npu_inst_int_data_res_4__2__6_), .A2(
        npu_inst_pe_1_4_2_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_4_2_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_2_U108 ( .A(npu_inst_int_data_res_4__2__7_), .B(
        npu_inst_pe_1_4_2_sub_77_carry_7_), .ZN(npu_inst_pe_1_4_2_N72) );
  INV_X1 npu_inst_pe_1_4_2_U107 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_4_2_n6)
         );
  INV_X1 npu_inst_pe_1_4_2_U106 ( .A(npu_inst_pe_1_4_2_n6), .ZN(
        npu_inst_pe_1_4_2_n5) );
  INV_X1 npu_inst_pe_1_4_2_U105 ( .A(npu_inst_n38), .ZN(npu_inst_pe_1_4_2_n2)
         );
  AOI22_X1 npu_inst_pe_1_4_2_U104 ( .A1(npu_inst_int_data_y_5__2__0_), .A2(
        npu_inst_pe_1_4_2_n58), .B1(npu_inst_pe_1_4_2_n118), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_2_n57) );
  INV_X1 npu_inst_pe_1_4_2_U103 ( .A(npu_inst_pe_1_4_2_n57), .ZN(
        npu_inst_pe_1_4_2_n107) );
  AOI22_X1 npu_inst_pe_1_4_2_U102 ( .A1(npu_inst_int_data_y_5__2__0_), .A2(
        npu_inst_pe_1_4_2_n54), .B1(npu_inst_pe_1_4_2_n117), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_2_n53) );
  INV_X1 npu_inst_pe_1_4_2_U99 ( .A(npu_inst_pe_1_4_2_n53), .ZN(
        npu_inst_pe_1_4_2_n108) );
  AOI22_X1 npu_inst_pe_1_4_2_U98 ( .A1(npu_inst_int_data_y_5__2__0_), .A2(
        npu_inst_pe_1_4_2_n50), .B1(npu_inst_pe_1_4_2_n116), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_2_n49) );
  INV_X1 npu_inst_pe_1_4_2_U97 ( .A(npu_inst_pe_1_4_2_n49), .ZN(
        npu_inst_pe_1_4_2_n109) );
  AOI22_X1 npu_inst_pe_1_4_2_U96 ( .A1(npu_inst_int_data_y_5__2__0_), .A2(
        npu_inst_pe_1_4_2_n46), .B1(npu_inst_pe_1_4_2_n115), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_2_n45) );
  INV_X1 npu_inst_pe_1_4_2_U95 ( .A(npu_inst_pe_1_4_2_n45), .ZN(
        npu_inst_pe_1_4_2_n110) );
  AOI22_X1 npu_inst_pe_1_4_2_U94 ( .A1(npu_inst_int_data_y_5__2__0_), .A2(
        npu_inst_pe_1_4_2_n42), .B1(npu_inst_pe_1_4_2_n114), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_2_n41) );
  INV_X1 npu_inst_pe_1_4_2_U93 ( .A(npu_inst_pe_1_4_2_n41), .ZN(
        npu_inst_pe_1_4_2_n111) );
  AOI22_X1 npu_inst_pe_1_4_2_U92 ( .A1(npu_inst_int_data_y_5__2__1_), .A2(
        npu_inst_pe_1_4_2_n58), .B1(npu_inst_pe_1_4_2_n118), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_2_n59) );
  INV_X1 npu_inst_pe_1_4_2_U91 ( .A(npu_inst_pe_1_4_2_n59), .ZN(
        npu_inst_pe_1_4_2_n101) );
  AOI22_X1 npu_inst_pe_1_4_2_U90 ( .A1(npu_inst_int_data_y_5__2__1_), .A2(
        npu_inst_pe_1_4_2_n54), .B1(npu_inst_pe_1_4_2_n117), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_2_n55) );
  INV_X1 npu_inst_pe_1_4_2_U89 ( .A(npu_inst_pe_1_4_2_n55), .ZN(
        npu_inst_pe_1_4_2_n102) );
  AOI22_X1 npu_inst_pe_1_4_2_U88 ( .A1(npu_inst_int_data_y_5__2__1_), .A2(
        npu_inst_pe_1_4_2_n50), .B1(npu_inst_pe_1_4_2_n116), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_2_n51) );
  INV_X1 npu_inst_pe_1_4_2_U87 ( .A(npu_inst_pe_1_4_2_n51), .ZN(
        npu_inst_pe_1_4_2_n103) );
  AOI22_X1 npu_inst_pe_1_4_2_U86 ( .A1(npu_inst_int_data_y_5__2__1_), .A2(
        npu_inst_pe_1_4_2_n46), .B1(npu_inst_pe_1_4_2_n115), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_2_n47) );
  INV_X1 npu_inst_pe_1_4_2_U85 ( .A(npu_inst_pe_1_4_2_n47), .ZN(
        npu_inst_pe_1_4_2_n104) );
  AOI22_X1 npu_inst_pe_1_4_2_U84 ( .A1(npu_inst_int_data_y_5__2__1_), .A2(
        npu_inst_pe_1_4_2_n42), .B1(npu_inst_pe_1_4_2_n114), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_2_n43) );
  INV_X1 npu_inst_pe_1_4_2_U83 ( .A(npu_inst_pe_1_4_2_n43), .ZN(
        npu_inst_pe_1_4_2_n105) );
  AOI22_X1 npu_inst_pe_1_4_2_U82 ( .A1(npu_inst_pe_1_4_2_n38), .A2(
        npu_inst_int_data_y_5__2__1_), .B1(npu_inst_pe_1_4_2_n113), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_2_n39) );
  INV_X1 npu_inst_pe_1_4_2_U81 ( .A(npu_inst_pe_1_4_2_n39), .ZN(
        npu_inst_pe_1_4_2_n106) );
  AND2_X1 npu_inst_pe_1_4_2_U80 ( .A1(npu_inst_pe_1_4_2_N93), .A2(npu_inst_n38), .ZN(npu_inst_int_data_y_4__2__0_) );
  NAND2_X1 npu_inst_pe_1_4_2_U79 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_2_n60), .ZN(npu_inst_pe_1_4_2_n74) );
  OAI21_X1 npu_inst_pe_1_4_2_U78 ( .B1(npu_inst_pe_1_4_2_n63), .B2(
        npu_inst_pe_1_4_2_n60), .A(npu_inst_pe_1_4_2_n74), .ZN(
        npu_inst_pe_1_4_2_n97) );
  NAND2_X1 npu_inst_pe_1_4_2_U77 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_2_n60), .ZN(npu_inst_pe_1_4_2_n73) );
  OAI21_X1 npu_inst_pe_1_4_2_U76 ( .B1(npu_inst_pe_1_4_2_n61), .B2(
        npu_inst_pe_1_4_2_n60), .A(npu_inst_pe_1_4_2_n73), .ZN(
        npu_inst_pe_1_4_2_n96) );
  NAND2_X1 npu_inst_pe_1_4_2_U75 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_2_n56), .ZN(npu_inst_pe_1_4_2_n72) );
  OAI21_X1 npu_inst_pe_1_4_2_U74 ( .B1(npu_inst_pe_1_4_2_n63), .B2(
        npu_inst_pe_1_4_2_n56), .A(npu_inst_pe_1_4_2_n72), .ZN(
        npu_inst_pe_1_4_2_n95) );
  NAND2_X1 npu_inst_pe_1_4_2_U73 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_2_n56), .ZN(npu_inst_pe_1_4_2_n71) );
  OAI21_X1 npu_inst_pe_1_4_2_U72 ( .B1(npu_inst_pe_1_4_2_n61), .B2(
        npu_inst_pe_1_4_2_n56), .A(npu_inst_pe_1_4_2_n71), .ZN(
        npu_inst_pe_1_4_2_n94) );
  NAND2_X1 npu_inst_pe_1_4_2_U71 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_2_n52), .ZN(npu_inst_pe_1_4_2_n70) );
  OAI21_X1 npu_inst_pe_1_4_2_U70 ( .B1(npu_inst_pe_1_4_2_n63), .B2(
        npu_inst_pe_1_4_2_n52), .A(npu_inst_pe_1_4_2_n70), .ZN(
        npu_inst_pe_1_4_2_n93) );
  NAND2_X1 npu_inst_pe_1_4_2_U69 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_2_n52), .ZN(npu_inst_pe_1_4_2_n69) );
  OAI21_X1 npu_inst_pe_1_4_2_U68 ( .B1(npu_inst_pe_1_4_2_n61), .B2(
        npu_inst_pe_1_4_2_n52), .A(npu_inst_pe_1_4_2_n69), .ZN(
        npu_inst_pe_1_4_2_n92) );
  NAND2_X1 npu_inst_pe_1_4_2_U67 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_2_n48), .ZN(npu_inst_pe_1_4_2_n68) );
  OAI21_X1 npu_inst_pe_1_4_2_U66 ( .B1(npu_inst_pe_1_4_2_n63), .B2(
        npu_inst_pe_1_4_2_n48), .A(npu_inst_pe_1_4_2_n68), .ZN(
        npu_inst_pe_1_4_2_n91) );
  NAND2_X1 npu_inst_pe_1_4_2_U65 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_2_n48), .ZN(npu_inst_pe_1_4_2_n67) );
  OAI21_X1 npu_inst_pe_1_4_2_U64 ( .B1(npu_inst_pe_1_4_2_n61), .B2(
        npu_inst_pe_1_4_2_n48), .A(npu_inst_pe_1_4_2_n67), .ZN(
        npu_inst_pe_1_4_2_n90) );
  NAND2_X1 npu_inst_pe_1_4_2_U63 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_2_n44), .ZN(npu_inst_pe_1_4_2_n66) );
  OAI21_X1 npu_inst_pe_1_4_2_U62 ( .B1(npu_inst_pe_1_4_2_n63), .B2(
        npu_inst_pe_1_4_2_n44), .A(npu_inst_pe_1_4_2_n66), .ZN(
        npu_inst_pe_1_4_2_n89) );
  NAND2_X1 npu_inst_pe_1_4_2_U61 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_2_n44), .ZN(npu_inst_pe_1_4_2_n65) );
  OAI21_X1 npu_inst_pe_1_4_2_U60 ( .B1(npu_inst_pe_1_4_2_n61), .B2(
        npu_inst_pe_1_4_2_n44), .A(npu_inst_pe_1_4_2_n65), .ZN(
        npu_inst_pe_1_4_2_n88) );
  NAND2_X1 npu_inst_pe_1_4_2_U59 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_2_n40), .ZN(npu_inst_pe_1_4_2_n64) );
  OAI21_X1 npu_inst_pe_1_4_2_U58 ( .B1(npu_inst_pe_1_4_2_n63), .B2(
        npu_inst_pe_1_4_2_n40), .A(npu_inst_pe_1_4_2_n64), .ZN(
        npu_inst_pe_1_4_2_n87) );
  NAND2_X1 npu_inst_pe_1_4_2_U57 ( .A1(npu_inst_pe_1_4_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_2_n40), .ZN(npu_inst_pe_1_4_2_n62) );
  OAI21_X1 npu_inst_pe_1_4_2_U56 ( .B1(npu_inst_pe_1_4_2_n61), .B2(
        npu_inst_pe_1_4_2_n40), .A(npu_inst_pe_1_4_2_n62), .ZN(
        npu_inst_pe_1_4_2_n86) );
  AOI22_X1 npu_inst_pe_1_4_2_U55 ( .A1(npu_inst_pe_1_4_2_n38), .A2(
        npu_inst_int_data_y_5__2__0_), .B1(npu_inst_pe_1_4_2_n113), .B2(
        npu_inst_pe_1_4_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_2_n37) );
  INV_X1 npu_inst_pe_1_4_2_U54 ( .A(npu_inst_pe_1_4_2_n37), .ZN(
        npu_inst_pe_1_4_2_n112) );
  AND2_X1 npu_inst_pe_1_4_2_U53 ( .A1(npu_inst_n38), .A2(npu_inst_pe_1_4_2_N94), .ZN(npu_inst_int_data_y_4__2__1_) );
  AOI222_X1 npu_inst_pe_1_4_2_U52 ( .A1(npu_inst_int_data_res_5__2__0_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N73), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N65), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n84) );
  INV_X1 npu_inst_pe_1_4_2_U51 ( .A(npu_inst_pe_1_4_2_n84), .ZN(
        npu_inst_pe_1_4_2_n100) );
  AOI222_X1 npu_inst_pe_1_4_2_U50 ( .A1(npu_inst_pe_1_4_2_n1), .A2(
        npu_inst_int_data_res_5__2__7_), .B1(npu_inst_pe_1_4_2_N80), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N72), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n75) );
  INV_X1 npu_inst_pe_1_4_2_U49 ( .A(npu_inst_pe_1_4_2_n75), .ZN(
        npu_inst_pe_1_4_2_n32) );
  AOI222_X1 npu_inst_pe_1_4_2_U48 ( .A1(npu_inst_int_data_res_5__2__1_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N74), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N66), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n83) );
  INV_X1 npu_inst_pe_1_4_2_U47 ( .A(npu_inst_pe_1_4_2_n83), .ZN(
        npu_inst_pe_1_4_2_n99) );
  AOI222_X1 npu_inst_pe_1_4_2_U46 ( .A1(npu_inst_int_data_res_5__2__3_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N76), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N68), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n81) );
  INV_X1 npu_inst_pe_1_4_2_U45 ( .A(npu_inst_pe_1_4_2_n81), .ZN(
        npu_inst_pe_1_4_2_n36) );
  AOI222_X1 npu_inst_pe_1_4_2_U44 ( .A1(npu_inst_int_data_res_5__2__4_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N77), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N69), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n80) );
  INV_X1 npu_inst_pe_1_4_2_U43 ( .A(npu_inst_pe_1_4_2_n80), .ZN(
        npu_inst_pe_1_4_2_n35) );
  AOI222_X1 npu_inst_pe_1_4_2_U42 ( .A1(npu_inst_int_data_res_5__2__5_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N78), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N70), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n79) );
  INV_X1 npu_inst_pe_1_4_2_U41 ( .A(npu_inst_pe_1_4_2_n79), .ZN(
        npu_inst_pe_1_4_2_n34) );
  AOI222_X1 npu_inst_pe_1_4_2_U40 ( .A1(npu_inst_int_data_res_5__2__6_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N79), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N71), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n78) );
  INV_X1 npu_inst_pe_1_4_2_U39 ( .A(npu_inst_pe_1_4_2_n78), .ZN(
        npu_inst_pe_1_4_2_n33) );
  AND2_X1 npu_inst_pe_1_4_2_U38 ( .A1(npu_inst_int_data_x_4__2__1_), .A2(
        npu_inst_pe_1_4_2_int_q_weight_1_), .ZN(npu_inst_pe_1_4_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_2_U37 ( .A1(npu_inst_int_data_x_4__2__0_), .A2(
        npu_inst_pe_1_4_2_int_q_weight_1_), .ZN(npu_inst_pe_1_4_2_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_4_2_U36 ( .A(npu_inst_pe_1_4_2_int_data_1_), .ZN(
        npu_inst_pe_1_4_2_n13) );
  NOR3_X1 npu_inst_pe_1_4_2_U35 ( .A1(npu_inst_pe_1_4_2_n26), .A2(npu_inst_n38), .A3(npu_inst_int_ckg[29]), .ZN(npu_inst_pe_1_4_2_n85) );
  OR2_X1 npu_inst_pe_1_4_2_U34 ( .A1(npu_inst_pe_1_4_2_n85), .A2(
        npu_inst_pe_1_4_2_n1), .ZN(npu_inst_pe_1_4_2_N84) );
  AOI222_X1 npu_inst_pe_1_4_2_U33 ( .A1(npu_inst_int_data_res_5__2__2_), .A2(
        npu_inst_pe_1_4_2_n1), .B1(npu_inst_pe_1_4_2_N75), .B2(
        npu_inst_pe_1_4_2_n76), .C1(npu_inst_pe_1_4_2_N67), .C2(
        npu_inst_pe_1_4_2_n77), .ZN(npu_inst_pe_1_4_2_n82) );
  INV_X1 npu_inst_pe_1_4_2_U32 ( .A(npu_inst_pe_1_4_2_n82), .ZN(
        npu_inst_pe_1_4_2_n98) );
  AOI22_X1 npu_inst_pe_1_4_2_U31 ( .A1(npu_inst_n38), .A2(
        npu_inst_int_data_y_5__2__1_), .B1(npu_inst_pe_1_4_2_n2), .B2(
        npu_inst_int_data_x_4__3__1_), .ZN(npu_inst_pe_1_4_2_n63) );
  AOI22_X1 npu_inst_pe_1_4_2_U30 ( .A1(npu_inst_n38), .A2(
        npu_inst_int_data_y_5__2__0_), .B1(npu_inst_pe_1_4_2_n2), .B2(
        npu_inst_int_data_x_4__3__0_), .ZN(npu_inst_pe_1_4_2_n61) );
  INV_X1 npu_inst_pe_1_4_2_U29 ( .A(npu_inst_pe_1_4_2_int_data_0_), .ZN(
        npu_inst_pe_1_4_2_n12) );
  INV_X1 npu_inst_pe_1_4_2_U28 ( .A(npu_inst_n51), .ZN(npu_inst_pe_1_4_2_n4)
         );
  OR3_X1 npu_inst_pe_1_4_2_U27 ( .A1(npu_inst_pe_1_4_2_n5), .A2(
        npu_inst_pe_1_4_2_n7), .A3(npu_inst_pe_1_4_2_n4), .ZN(
        npu_inst_pe_1_4_2_n56) );
  OR3_X1 npu_inst_pe_1_4_2_U26 ( .A1(npu_inst_pe_1_4_2_n4), .A2(
        npu_inst_pe_1_4_2_n7), .A3(npu_inst_pe_1_4_2_n6), .ZN(
        npu_inst_pe_1_4_2_n48) );
  INV_X1 npu_inst_pe_1_4_2_U25 ( .A(npu_inst_pe_1_4_2_n4), .ZN(
        npu_inst_pe_1_4_2_n3) );
  OR3_X1 npu_inst_pe_1_4_2_U24 ( .A1(npu_inst_pe_1_4_2_n3), .A2(
        npu_inst_pe_1_4_2_n7), .A3(npu_inst_pe_1_4_2_n6), .ZN(
        npu_inst_pe_1_4_2_n52) );
  OR3_X1 npu_inst_pe_1_4_2_U23 ( .A1(npu_inst_pe_1_4_2_n5), .A2(
        npu_inst_pe_1_4_2_n7), .A3(npu_inst_pe_1_4_2_n3), .ZN(
        npu_inst_pe_1_4_2_n60) );
  BUF_X1 npu_inst_pe_1_4_2_U22 ( .A(npu_inst_n20), .Z(npu_inst_pe_1_4_2_n1) );
  NOR2_X1 npu_inst_pe_1_4_2_U21 ( .A1(npu_inst_pe_1_4_2_n60), .A2(
        npu_inst_pe_1_4_2_n2), .ZN(npu_inst_pe_1_4_2_n58) );
  NOR2_X1 npu_inst_pe_1_4_2_U20 ( .A1(npu_inst_pe_1_4_2_n56), .A2(
        npu_inst_pe_1_4_2_n2), .ZN(npu_inst_pe_1_4_2_n54) );
  NOR2_X1 npu_inst_pe_1_4_2_U19 ( .A1(npu_inst_pe_1_4_2_n52), .A2(
        npu_inst_pe_1_4_2_n2), .ZN(npu_inst_pe_1_4_2_n50) );
  NOR2_X1 npu_inst_pe_1_4_2_U18 ( .A1(npu_inst_pe_1_4_2_n48), .A2(
        npu_inst_pe_1_4_2_n2), .ZN(npu_inst_pe_1_4_2_n46) );
  NOR2_X1 npu_inst_pe_1_4_2_U17 ( .A1(npu_inst_pe_1_4_2_n40), .A2(
        npu_inst_pe_1_4_2_n2), .ZN(npu_inst_pe_1_4_2_n38) );
  NOR2_X1 npu_inst_pe_1_4_2_U16 ( .A1(npu_inst_pe_1_4_2_n44), .A2(
        npu_inst_pe_1_4_2_n2), .ZN(npu_inst_pe_1_4_2_n42) );
  BUF_X1 npu_inst_pe_1_4_2_U15 ( .A(npu_inst_n81), .Z(npu_inst_pe_1_4_2_n7) );
  INV_X1 npu_inst_pe_1_4_2_U14 ( .A(npu_inst_n106), .ZN(npu_inst_pe_1_4_2_n11)
         );
  INV_X1 npu_inst_pe_1_4_2_U13 ( .A(npu_inst_pe_1_4_2_n38), .ZN(
        npu_inst_pe_1_4_2_n113) );
  INV_X1 npu_inst_pe_1_4_2_U12 ( .A(npu_inst_pe_1_4_2_n58), .ZN(
        npu_inst_pe_1_4_2_n118) );
  INV_X1 npu_inst_pe_1_4_2_U11 ( .A(npu_inst_pe_1_4_2_n54), .ZN(
        npu_inst_pe_1_4_2_n117) );
  INV_X1 npu_inst_pe_1_4_2_U10 ( .A(npu_inst_pe_1_4_2_n50), .ZN(
        npu_inst_pe_1_4_2_n116) );
  INV_X1 npu_inst_pe_1_4_2_U9 ( .A(npu_inst_pe_1_4_2_n46), .ZN(
        npu_inst_pe_1_4_2_n115) );
  INV_X1 npu_inst_pe_1_4_2_U8 ( .A(npu_inst_pe_1_4_2_n42), .ZN(
        npu_inst_pe_1_4_2_n114) );
  BUF_X1 npu_inst_pe_1_4_2_U7 ( .A(npu_inst_pe_1_4_2_n11), .Z(
        npu_inst_pe_1_4_2_n10) );
  BUF_X1 npu_inst_pe_1_4_2_U6 ( .A(npu_inst_pe_1_4_2_n11), .Z(
        npu_inst_pe_1_4_2_n9) );
  BUF_X1 npu_inst_pe_1_4_2_U5 ( .A(npu_inst_pe_1_4_2_n11), .Z(
        npu_inst_pe_1_4_2_n8) );
  NOR2_X1 npu_inst_pe_1_4_2_U4 ( .A1(npu_inst_pe_1_4_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_2_n1), .ZN(npu_inst_pe_1_4_2_n76) );
  NOR2_X1 npu_inst_pe_1_4_2_U3 ( .A1(npu_inst_pe_1_4_2_n27), .A2(
        npu_inst_pe_1_4_2_n1), .ZN(npu_inst_pe_1_4_2_n77) );
  FA_X1 npu_inst_pe_1_4_2_sub_77_U2_1 ( .A(npu_inst_int_data_res_4__2__1_), 
        .B(npu_inst_pe_1_4_2_n13), .CI(npu_inst_pe_1_4_2_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_4_2_sub_77_carry_2_), .S(npu_inst_pe_1_4_2_N66) );
  FA_X1 npu_inst_pe_1_4_2_add_79_U1_1 ( .A(npu_inst_int_data_res_4__2__1_), 
        .B(npu_inst_pe_1_4_2_int_data_1_), .CI(
        npu_inst_pe_1_4_2_add_79_carry_1_), .CO(
        npu_inst_pe_1_4_2_add_79_carry_2_), .S(npu_inst_pe_1_4_2_N74) );
  NAND3_X1 npu_inst_pe_1_4_2_U101 ( .A1(npu_inst_pe_1_4_2_n4), .A2(
        npu_inst_pe_1_4_2_n6), .A3(npu_inst_pe_1_4_2_n7), .ZN(
        npu_inst_pe_1_4_2_n44) );
  NAND3_X1 npu_inst_pe_1_4_2_U100 ( .A1(npu_inst_pe_1_4_2_n3), .A2(
        npu_inst_pe_1_4_2_n6), .A3(npu_inst_pe_1_4_2_n7), .ZN(
        npu_inst_pe_1_4_2_n40) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_2_n33), .CK(
        npu_inst_pe_1_4_2_net3696), .RN(npu_inst_pe_1_4_2_n8), .Q(
        npu_inst_int_data_res_4__2__6_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_2_n34), .CK(
        npu_inst_pe_1_4_2_net3696), .RN(npu_inst_pe_1_4_2_n8), .Q(
        npu_inst_int_data_res_4__2__5_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_2_n35), .CK(
        npu_inst_pe_1_4_2_net3696), .RN(npu_inst_pe_1_4_2_n8), .Q(
        npu_inst_int_data_res_4__2__4_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_2_n36), .CK(
        npu_inst_pe_1_4_2_net3696), .RN(npu_inst_pe_1_4_2_n8), .Q(
        npu_inst_int_data_res_4__2__3_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_2_n98), .CK(
        npu_inst_pe_1_4_2_net3696), .RN(npu_inst_pe_1_4_2_n8), .Q(
        npu_inst_int_data_res_4__2__2_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_2_n99), .CK(
        npu_inst_pe_1_4_2_net3696), .RN(npu_inst_pe_1_4_2_n8), .Q(
        npu_inst_int_data_res_4__2__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_2_n32), .CK(
        npu_inst_pe_1_4_2_net3696), .RN(npu_inst_pe_1_4_2_n8), .Q(
        npu_inst_int_data_res_4__2__7_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_2_n100), 
        .CK(npu_inst_pe_1_4_2_net3696), .RN(npu_inst_pe_1_4_2_n8), .Q(
        npu_inst_int_data_res_4__2__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_weight_reg_0_ ( .D(npu_inst_n92), .CK(
        npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n8), .Q(
        npu_inst_pe_1_4_2_int_q_weight_0_), .QN(npu_inst_pe_1_4_2_n27) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_weight_reg_1_ ( .D(npu_inst_n98), .CK(
        npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n8), .Q(
        npu_inst_pe_1_4_2_int_q_weight_1_), .QN(npu_inst_pe_1_4_2_n26) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_2_n112), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n8), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_2_n106), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n8), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_2_n111), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_2_n105), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_2_n110), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_2_n104), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_2_n109), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_2_n103), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_2_n108), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_2_n102), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_2_n107), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_2_n101), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_2_n86), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_2_n87), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n9), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_2_n88), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_2_n89), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_2_n90), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_2_n91), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_2_n92), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_2_n93), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_2_n94), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_2_n95), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_2_n96), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_2_n97), 
        .CK(npu_inst_pe_1_4_2_net3702), .RN(npu_inst_pe_1_4_2_n10), .Q(
        npu_inst_pe_1_4_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_2_net3696) );
  CLKGATETST_X1 npu_inst_pe_1_4_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n45), .SE(1'b0), .GCK(npu_inst_pe_1_4_2_net3702) );
  MUX2_X1 npu_inst_pe_1_4_3_U153 ( .A(npu_inst_pe_1_4_3_n31), .B(
        npu_inst_pe_1_4_3_n28), .S(npu_inst_pe_1_4_3_n7), .Z(
        npu_inst_pe_1_4_3_N93) );
  MUX2_X1 npu_inst_pe_1_4_3_U152 ( .A(npu_inst_pe_1_4_3_n30), .B(
        npu_inst_pe_1_4_3_n29), .S(npu_inst_pe_1_4_3_n5), .Z(
        npu_inst_pe_1_4_3_n31) );
  MUX2_X1 npu_inst_pe_1_4_3_U151 ( .A(npu_inst_pe_1_4_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_3_n3), .Z(
        npu_inst_pe_1_4_3_n30) );
  MUX2_X1 npu_inst_pe_1_4_3_U150 ( .A(npu_inst_pe_1_4_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_3_n3), .Z(
        npu_inst_pe_1_4_3_n29) );
  MUX2_X1 npu_inst_pe_1_4_3_U149 ( .A(npu_inst_pe_1_4_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_3_n3), .Z(
        npu_inst_pe_1_4_3_n28) );
  MUX2_X1 npu_inst_pe_1_4_3_U148 ( .A(npu_inst_pe_1_4_3_n25), .B(
        npu_inst_pe_1_4_3_n22), .S(npu_inst_pe_1_4_3_n7), .Z(
        npu_inst_pe_1_4_3_N94) );
  MUX2_X1 npu_inst_pe_1_4_3_U147 ( .A(npu_inst_pe_1_4_3_n24), .B(
        npu_inst_pe_1_4_3_n23), .S(npu_inst_pe_1_4_3_n5), .Z(
        npu_inst_pe_1_4_3_n25) );
  MUX2_X1 npu_inst_pe_1_4_3_U146 ( .A(npu_inst_pe_1_4_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_3_n3), .Z(
        npu_inst_pe_1_4_3_n24) );
  MUX2_X1 npu_inst_pe_1_4_3_U145 ( .A(npu_inst_pe_1_4_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_3_n3), .Z(
        npu_inst_pe_1_4_3_n23) );
  MUX2_X1 npu_inst_pe_1_4_3_U144 ( .A(npu_inst_pe_1_4_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_3_n3), .Z(
        npu_inst_pe_1_4_3_n22) );
  MUX2_X1 npu_inst_pe_1_4_3_U143 ( .A(npu_inst_pe_1_4_3_n21), .B(
        npu_inst_pe_1_4_3_n18), .S(npu_inst_pe_1_4_3_n7), .Z(
        npu_inst_int_data_x_4__3__1_) );
  MUX2_X1 npu_inst_pe_1_4_3_U142 ( .A(npu_inst_pe_1_4_3_n20), .B(
        npu_inst_pe_1_4_3_n19), .S(npu_inst_pe_1_4_3_n5), .Z(
        npu_inst_pe_1_4_3_n21) );
  MUX2_X1 npu_inst_pe_1_4_3_U141 ( .A(npu_inst_pe_1_4_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_3_n3), .Z(
        npu_inst_pe_1_4_3_n20) );
  MUX2_X1 npu_inst_pe_1_4_3_U140 ( .A(npu_inst_pe_1_4_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_3_n3), .Z(
        npu_inst_pe_1_4_3_n19) );
  MUX2_X1 npu_inst_pe_1_4_3_U139 ( .A(npu_inst_pe_1_4_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_3_n3), .Z(
        npu_inst_pe_1_4_3_n18) );
  MUX2_X1 npu_inst_pe_1_4_3_U138 ( .A(npu_inst_pe_1_4_3_n17), .B(
        npu_inst_pe_1_4_3_n14), .S(npu_inst_pe_1_4_3_n7), .Z(
        npu_inst_int_data_x_4__3__0_) );
  MUX2_X1 npu_inst_pe_1_4_3_U137 ( .A(npu_inst_pe_1_4_3_n16), .B(
        npu_inst_pe_1_4_3_n15), .S(npu_inst_pe_1_4_3_n5), .Z(
        npu_inst_pe_1_4_3_n17) );
  MUX2_X1 npu_inst_pe_1_4_3_U136 ( .A(npu_inst_pe_1_4_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_3_n3), .Z(
        npu_inst_pe_1_4_3_n16) );
  MUX2_X1 npu_inst_pe_1_4_3_U135 ( .A(npu_inst_pe_1_4_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_3_n3), .Z(
        npu_inst_pe_1_4_3_n15) );
  MUX2_X1 npu_inst_pe_1_4_3_U134 ( .A(npu_inst_pe_1_4_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_3_n3), .Z(
        npu_inst_pe_1_4_3_n14) );
  XOR2_X1 npu_inst_pe_1_4_3_U133 ( .A(npu_inst_pe_1_4_3_int_data_0_), .B(
        npu_inst_int_data_res_4__3__0_), .Z(npu_inst_pe_1_4_3_N73) );
  AND2_X1 npu_inst_pe_1_4_3_U132 ( .A1(npu_inst_int_data_res_4__3__0_), .A2(
        npu_inst_pe_1_4_3_int_data_0_), .ZN(npu_inst_pe_1_4_3_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_3_U131 ( .A(npu_inst_int_data_res_4__3__0_), .B(
        npu_inst_pe_1_4_3_n12), .ZN(npu_inst_pe_1_4_3_N65) );
  OR2_X1 npu_inst_pe_1_4_3_U130 ( .A1(npu_inst_pe_1_4_3_n12), .A2(
        npu_inst_int_data_res_4__3__0_), .ZN(npu_inst_pe_1_4_3_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_3_U129 ( .A(npu_inst_int_data_res_4__3__2_), .B(
        npu_inst_pe_1_4_3_add_79_carry_2_), .Z(npu_inst_pe_1_4_3_N75) );
  AND2_X1 npu_inst_pe_1_4_3_U128 ( .A1(npu_inst_pe_1_4_3_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_4__3__2_), .ZN(
        npu_inst_pe_1_4_3_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_3_U127 ( .A(npu_inst_int_data_res_4__3__3_), .B(
        npu_inst_pe_1_4_3_add_79_carry_3_), .Z(npu_inst_pe_1_4_3_N76) );
  AND2_X1 npu_inst_pe_1_4_3_U126 ( .A1(npu_inst_pe_1_4_3_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_4__3__3_), .ZN(
        npu_inst_pe_1_4_3_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_3_U125 ( .A(npu_inst_int_data_res_4__3__4_), .B(
        npu_inst_pe_1_4_3_add_79_carry_4_), .Z(npu_inst_pe_1_4_3_N77) );
  AND2_X1 npu_inst_pe_1_4_3_U124 ( .A1(npu_inst_pe_1_4_3_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_4__3__4_), .ZN(
        npu_inst_pe_1_4_3_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_3_U123 ( .A(npu_inst_int_data_res_4__3__5_), .B(
        npu_inst_pe_1_4_3_add_79_carry_5_), .Z(npu_inst_pe_1_4_3_N78) );
  AND2_X1 npu_inst_pe_1_4_3_U122 ( .A1(npu_inst_pe_1_4_3_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_4__3__5_), .ZN(
        npu_inst_pe_1_4_3_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_3_U121 ( .A(npu_inst_int_data_res_4__3__6_), .B(
        npu_inst_pe_1_4_3_add_79_carry_6_), .Z(npu_inst_pe_1_4_3_N79) );
  AND2_X1 npu_inst_pe_1_4_3_U120 ( .A1(npu_inst_pe_1_4_3_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_4__3__6_), .ZN(
        npu_inst_pe_1_4_3_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_3_U119 ( .A(npu_inst_int_data_res_4__3__7_), .B(
        npu_inst_pe_1_4_3_add_79_carry_7_), .Z(npu_inst_pe_1_4_3_N80) );
  XNOR2_X1 npu_inst_pe_1_4_3_U118 ( .A(npu_inst_pe_1_4_3_sub_77_carry_2_), .B(
        npu_inst_int_data_res_4__3__2_), .ZN(npu_inst_pe_1_4_3_N67) );
  OR2_X1 npu_inst_pe_1_4_3_U117 ( .A1(npu_inst_int_data_res_4__3__2_), .A2(
        npu_inst_pe_1_4_3_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_4_3_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_3_U116 ( .A(npu_inst_pe_1_4_3_sub_77_carry_3_), .B(
        npu_inst_int_data_res_4__3__3_), .ZN(npu_inst_pe_1_4_3_N68) );
  OR2_X1 npu_inst_pe_1_4_3_U115 ( .A1(npu_inst_int_data_res_4__3__3_), .A2(
        npu_inst_pe_1_4_3_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_4_3_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_3_U114 ( .A(npu_inst_pe_1_4_3_sub_77_carry_4_), .B(
        npu_inst_int_data_res_4__3__4_), .ZN(npu_inst_pe_1_4_3_N69) );
  OR2_X1 npu_inst_pe_1_4_3_U113 ( .A1(npu_inst_int_data_res_4__3__4_), .A2(
        npu_inst_pe_1_4_3_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_4_3_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_3_U112 ( .A(npu_inst_pe_1_4_3_sub_77_carry_5_), .B(
        npu_inst_int_data_res_4__3__5_), .ZN(npu_inst_pe_1_4_3_N70) );
  OR2_X1 npu_inst_pe_1_4_3_U111 ( .A1(npu_inst_int_data_res_4__3__5_), .A2(
        npu_inst_pe_1_4_3_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_4_3_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_3_U110 ( .A(npu_inst_pe_1_4_3_sub_77_carry_6_), .B(
        npu_inst_int_data_res_4__3__6_), .ZN(npu_inst_pe_1_4_3_N71) );
  OR2_X1 npu_inst_pe_1_4_3_U109 ( .A1(npu_inst_int_data_res_4__3__6_), .A2(
        npu_inst_pe_1_4_3_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_4_3_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_3_U108 ( .A(npu_inst_int_data_res_4__3__7_), .B(
        npu_inst_pe_1_4_3_sub_77_carry_7_), .ZN(npu_inst_pe_1_4_3_N72) );
  INV_X1 npu_inst_pe_1_4_3_U107 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_4_3_n6)
         );
  INV_X1 npu_inst_pe_1_4_3_U106 ( .A(npu_inst_pe_1_4_3_n6), .ZN(
        npu_inst_pe_1_4_3_n5) );
  INV_X1 npu_inst_pe_1_4_3_U105 ( .A(npu_inst_n38), .ZN(npu_inst_pe_1_4_3_n2)
         );
  AOI22_X1 npu_inst_pe_1_4_3_U104 ( .A1(npu_inst_int_data_y_5__3__0_), .A2(
        npu_inst_pe_1_4_3_n58), .B1(npu_inst_pe_1_4_3_n118), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_3_n57) );
  INV_X1 npu_inst_pe_1_4_3_U103 ( .A(npu_inst_pe_1_4_3_n57), .ZN(
        npu_inst_pe_1_4_3_n107) );
  AOI22_X1 npu_inst_pe_1_4_3_U102 ( .A1(npu_inst_int_data_y_5__3__0_), .A2(
        npu_inst_pe_1_4_3_n54), .B1(npu_inst_pe_1_4_3_n117), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_3_n53) );
  INV_X1 npu_inst_pe_1_4_3_U99 ( .A(npu_inst_pe_1_4_3_n53), .ZN(
        npu_inst_pe_1_4_3_n108) );
  AOI22_X1 npu_inst_pe_1_4_3_U98 ( .A1(npu_inst_int_data_y_5__3__0_), .A2(
        npu_inst_pe_1_4_3_n50), .B1(npu_inst_pe_1_4_3_n116), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_3_n49) );
  INV_X1 npu_inst_pe_1_4_3_U97 ( .A(npu_inst_pe_1_4_3_n49), .ZN(
        npu_inst_pe_1_4_3_n109) );
  AOI22_X1 npu_inst_pe_1_4_3_U96 ( .A1(npu_inst_int_data_y_5__3__0_), .A2(
        npu_inst_pe_1_4_3_n46), .B1(npu_inst_pe_1_4_3_n115), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_3_n45) );
  INV_X1 npu_inst_pe_1_4_3_U95 ( .A(npu_inst_pe_1_4_3_n45), .ZN(
        npu_inst_pe_1_4_3_n110) );
  AOI22_X1 npu_inst_pe_1_4_3_U94 ( .A1(npu_inst_int_data_y_5__3__0_), .A2(
        npu_inst_pe_1_4_3_n42), .B1(npu_inst_pe_1_4_3_n114), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_3_n41) );
  INV_X1 npu_inst_pe_1_4_3_U93 ( .A(npu_inst_pe_1_4_3_n41), .ZN(
        npu_inst_pe_1_4_3_n111) );
  AOI22_X1 npu_inst_pe_1_4_3_U92 ( .A1(npu_inst_int_data_y_5__3__1_), .A2(
        npu_inst_pe_1_4_3_n58), .B1(npu_inst_pe_1_4_3_n118), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_3_n59) );
  INV_X1 npu_inst_pe_1_4_3_U91 ( .A(npu_inst_pe_1_4_3_n59), .ZN(
        npu_inst_pe_1_4_3_n101) );
  AOI22_X1 npu_inst_pe_1_4_3_U90 ( .A1(npu_inst_int_data_y_5__3__1_), .A2(
        npu_inst_pe_1_4_3_n54), .B1(npu_inst_pe_1_4_3_n117), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_3_n55) );
  INV_X1 npu_inst_pe_1_4_3_U89 ( .A(npu_inst_pe_1_4_3_n55), .ZN(
        npu_inst_pe_1_4_3_n102) );
  AOI22_X1 npu_inst_pe_1_4_3_U88 ( .A1(npu_inst_int_data_y_5__3__1_), .A2(
        npu_inst_pe_1_4_3_n50), .B1(npu_inst_pe_1_4_3_n116), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_3_n51) );
  INV_X1 npu_inst_pe_1_4_3_U87 ( .A(npu_inst_pe_1_4_3_n51), .ZN(
        npu_inst_pe_1_4_3_n103) );
  AOI22_X1 npu_inst_pe_1_4_3_U86 ( .A1(npu_inst_int_data_y_5__3__1_), .A2(
        npu_inst_pe_1_4_3_n46), .B1(npu_inst_pe_1_4_3_n115), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_3_n47) );
  INV_X1 npu_inst_pe_1_4_3_U85 ( .A(npu_inst_pe_1_4_3_n47), .ZN(
        npu_inst_pe_1_4_3_n104) );
  AOI22_X1 npu_inst_pe_1_4_3_U84 ( .A1(npu_inst_int_data_y_5__3__1_), .A2(
        npu_inst_pe_1_4_3_n42), .B1(npu_inst_pe_1_4_3_n114), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_3_n43) );
  INV_X1 npu_inst_pe_1_4_3_U83 ( .A(npu_inst_pe_1_4_3_n43), .ZN(
        npu_inst_pe_1_4_3_n105) );
  AOI22_X1 npu_inst_pe_1_4_3_U82 ( .A1(npu_inst_pe_1_4_3_n38), .A2(
        npu_inst_int_data_y_5__3__1_), .B1(npu_inst_pe_1_4_3_n113), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_3_n39) );
  INV_X1 npu_inst_pe_1_4_3_U81 ( .A(npu_inst_pe_1_4_3_n39), .ZN(
        npu_inst_pe_1_4_3_n106) );
  AND2_X1 npu_inst_pe_1_4_3_U80 ( .A1(npu_inst_pe_1_4_3_N93), .A2(npu_inst_n38), .ZN(npu_inst_int_data_y_4__3__0_) );
  NAND2_X1 npu_inst_pe_1_4_3_U79 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_3_n60), .ZN(npu_inst_pe_1_4_3_n74) );
  OAI21_X1 npu_inst_pe_1_4_3_U78 ( .B1(npu_inst_pe_1_4_3_n63), .B2(
        npu_inst_pe_1_4_3_n60), .A(npu_inst_pe_1_4_3_n74), .ZN(
        npu_inst_pe_1_4_3_n97) );
  NAND2_X1 npu_inst_pe_1_4_3_U77 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_3_n60), .ZN(npu_inst_pe_1_4_3_n73) );
  OAI21_X1 npu_inst_pe_1_4_3_U76 ( .B1(npu_inst_pe_1_4_3_n61), .B2(
        npu_inst_pe_1_4_3_n60), .A(npu_inst_pe_1_4_3_n73), .ZN(
        npu_inst_pe_1_4_3_n96) );
  NAND2_X1 npu_inst_pe_1_4_3_U75 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_3_n56), .ZN(npu_inst_pe_1_4_3_n72) );
  OAI21_X1 npu_inst_pe_1_4_3_U74 ( .B1(npu_inst_pe_1_4_3_n63), .B2(
        npu_inst_pe_1_4_3_n56), .A(npu_inst_pe_1_4_3_n72), .ZN(
        npu_inst_pe_1_4_3_n95) );
  NAND2_X1 npu_inst_pe_1_4_3_U73 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_3_n56), .ZN(npu_inst_pe_1_4_3_n71) );
  OAI21_X1 npu_inst_pe_1_4_3_U72 ( .B1(npu_inst_pe_1_4_3_n61), .B2(
        npu_inst_pe_1_4_3_n56), .A(npu_inst_pe_1_4_3_n71), .ZN(
        npu_inst_pe_1_4_3_n94) );
  NAND2_X1 npu_inst_pe_1_4_3_U71 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_3_n52), .ZN(npu_inst_pe_1_4_3_n70) );
  OAI21_X1 npu_inst_pe_1_4_3_U70 ( .B1(npu_inst_pe_1_4_3_n63), .B2(
        npu_inst_pe_1_4_3_n52), .A(npu_inst_pe_1_4_3_n70), .ZN(
        npu_inst_pe_1_4_3_n93) );
  NAND2_X1 npu_inst_pe_1_4_3_U69 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_3_n52), .ZN(npu_inst_pe_1_4_3_n69) );
  OAI21_X1 npu_inst_pe_1_4_3_U68 ( .B1(npu_inst_pe_1_4_3_n61), .B2(
        npu_inst_pe_1_4_3_n52), .A(npu_inst_pe_1_4_3_n69), .ZN(
        npu_inst_pe_1_4_3_n92) );
  NAND2_X1 npu_inst_pe_1_4_3_U67 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_3_n48), .ZN(npu_inst_pe_1_4_3_n68) );
  OAI21_X1 npu_inst_pe_1_4_3_U66 ( .B1(npu_inst_pe_1_4_3_n63), .B2(
        npu_inst_pe_1_4_3_n48), .A(npu_inst_pe_1_4_3_n68), .ZN(
        npu_inst_pe_1_4_3_n91) );
  NAND2_X1 npu_inst_pe_1_4_3_U65 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_3_n48), .ZN(npu_inst_pe_1_4_3_n67) );
  OAI21_X1 npu_inst_pe_1_4_3_U64 ( .B1(npu_inst_pe_1_4_3_n61), .B2(
        npu_inst_pe_1_4_3_n48), .A(npu_inst_pe_1_4_3_n67), .ZN(
        npu_inst_pe_1_4_3_n90) );
  NAND2_X1 npu_inst_pe_1_4_3_U63 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_3_n44), .ZN(npu_inst_pe_1_4_3_n66) );
  OAI21_X1 npu_inst_pe_1_4_3_U62 ( .B1(npu_inst_pe_1_4_3_n63), .B2(
        npu_inst_pe_1_4_3_n44), .A(npu_inst_pe_1_4_3_n66), .ZN(
        npu_inst_pe_1_4_3_n89) );
  NAND2_X1 npu_inst_pe_1_4_3_U61 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_3_n44), .ZN(npu_inst_pe_1_4_3_n65) );
  OAI21_X1 npu_inst_pe_1_4_3_U60 ( .B1(npu_inst_pe_1_4_3_n61), .B2(
        npu_inst_pe_1_4_3_n44), .A(npu_inst_pe_1_4_3_n65), .ZN(
        npu_inst_pe_1_4_3_n88) );
  NAND2_X1 npu_inst_pe_1_4_3_U59 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_3_n40), .ZN(npu_inst_pe_1_4_3_n64) );
  OAI21_X1 npu_inst_pe_1_4_3_U58 ( .B1(npu_inst_pe_1_4_3_n63), .B2(
        npu_inst_pe_1_4_3_n40), .A(npu_inst_pe_1_4_3_n64), .ZN(
        npu_inst_pe_1_4_3_n87) );
  NAND2_X1 npu_inst_pe_1_4_3_U57 ( .A1(npu_inst_pe_1_4_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_3_n40), .ZN(npu_inst_pe_1_4_3_n62) );
  OAI21_X1 npu_inst_pe_1_4_3_U56 ( .B1(npu_inst_pe_1_4_3_n61), .B2(
        npu_inst_pe_1_4_3_n40), .A(npu_inst_pe_1_4_3_n62), .ZN(
        npu_inst_pe_1_4_3_n86) );
  AOI22_X1 npu_inst_pe_1_4_3_U55 ( .A1(npu_inst_pe_1_4_3_n38), .A2(
        npu_inst_int_data_y_5__3__0_), .B1(npu_inst_pe_1_4_3_n113), .B2(
        npu_inst_pe_1_4_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_3_n37) );
  INV_X1 npu_inst_pe_1_4_3_U54 ( .A(npu_inst_pe_1_4_3_n37), .ZN(
        npu_inst_pe_1_4_3_n112) );
  AND2_X1 npu_inst_pe_1_4_3_U53 ( .A1(npu_inst_n38), .A2(npu_inst_pe_1_4_3_N94), .ZN(npu_inst_int_data_y_4__3__1_) );
  AOI222_X1 npu_inst_pe_1_4_3_U52 ( .A1(npu_inst_int_data_res_5__3__0_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N73), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N65), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n84) );
  INV_X1 npu_inst_pe_1_4_3_U51 ( .A(npu_inst_pe_1_4_3_n84), .ZN(
        npu_inst_pe_1_4_3_n100) );
  AOI222_X1 npu_inst_pe_1_4_3_U50 ( .A1(npu_inst_pe_1_4_3_n1), .A2(
        npu_inst_int_data_res_5__3__7_), .B1(npu_inst_pe_1_4_3_N80), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N72), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n75) );
  INV_X1 npu_inst_pe_1_4_3_U49 ( .A(npu_inst_pe_1_4_3_n75), .ZN(
        npu_inst_pe_1_4_3_n32) );
  AOI222_X1 npu_inst_pe_1_4_3_U48 ( .A1(npu_inst_int_data_res_5__3__1_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N74), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N66), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n83) );
  INV_X1 npu_inst_pe_1_4_3_U47 ( .A(npu_inst_pe_1_4_3_n83), .ZN(
        npu_inst_pe_1_4_3_n99) );
  AOI222_X1 npu_inst_pe_1_4_3_U46 ( .A1(npu_inst_int_data_res_5__3__3_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N76), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N68), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n81) );
  INV_X1 npu_inst_pe_1_4_3_U45 ( .A(npu_inst_pe_1_4_3_n81), .ZN(
        npu_inst_pe_1_4_3_n36) );
  AOI222_X1 npu_inst_pe_1_4_3_U44 ( .A1(npu_inst_int_data_res_5__3__4_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N77), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N69), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n80) );
  INV_X1 npu_inst_pe_1_4_3_U43 ( .A(npu_inst_pe_1_4_3_n80), .ZN(
        npu_inst_pe_1_4_3_n35) );
  AOI222_X1 npu_inst_pe_1_4_3_U42 ( .A1(npu_inst_int_data_res_5__3__5_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N78), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N70), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n79) );
  INV_X1 npu_inst_pe_1_4_3_U41 ( .A(npu_inst_pe_1_4_3_n79), .ZN(
        npu_inst_pe_1_4_3_n34) );
  AOI222_X1 npu_inst_pe_1_4_3_U40 ( .A1(npu_inst_int_data_res_5__3__6_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N79), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N71), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n78) );
  INV_X1 npu_inst_pe_1_4_3_U39 ( .A(npu_inst_pe_1_4_3_n78), .ZN(
        npu_inst_pe_1_4_3_n33) );
  AND2_X1 npu_inst_pe_1_4_3_U38 ( .A1(npu_inst_int_data_x_4__3__1_), .A2(
        npu_inst_pe_1_4_3_int_q_weight_1_), .ZN(npu_inst_pe_1_4_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_3_U37 ( .A1(npu_inst_int_data_x_4__3__0_), .A2(
        npu_inst_pe_1_4_3_int_q_weight_1_), .ZN(npu_inst_pe_1_4_3_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_4_3_U36 ( .A(npu_inst_pe_1_4_3_int_data_1_), .ZN(
        npu_inst_pe_1_4_3_n13) );
  NOR3_X1 npu_inst_pe_1_4_3_U35 ( .A1(npu_inst_pe_1_4_3_n26), .A2(npu_inst_n38), .A3(npu_inst_int_ckg[28]), .ZN(npu_inst_pe_1_4_3_n85) );
  OR2_X1 npu_inst_pe_1_4_3_U34 ( .A1(npu_inst_pe_1_4_3_n85), .A2(
        npu_inst_pe_1_4_3_n1), .ZN(npu_inst_pe_1_4_3_N84) );
  AOI222_X1 npu_inst_pe_1_4_3_U33 ( .A1(npu_inst_int_data_res_5__3__2_), .A2(
        npu_inst_pe_1_4_3_n1), .B1(npu_inst_pe_1_4_3_N75), .B2(
        npu_inst_pe_1_4_3_n76), .C1(npu_inst_pe_1_4_3_N67), .C2(
        npu_inst_pe_1_4_3_n77), .ZN(npu_inst_pe_1_4_3_n82) );
  INV_X1 npu_inst_pe_1_4_3_U32 ( .A(npu_inst_pe_1_4_3_n82), .ZN(
        npu_inst_pe_1_4_3_n98) );
  AOI22_X1 npu_inst_pe_1_4_3_U31 ( .A1(npu_inst_n38), .A2(
        npu_inst_int_data_y_5__3__1_), .B1(npu_inst_pe_1_4_3_n2), .B2(
        npu_inst_int_data_x_4__4__1_), .ZN(npu_inst_pe_1_4_3_n63) );
  AOI22_X1 npu_inst_pe_1_4_3_U30 ( .A1(npu_inst_n38), .A2(
        npu_inst_int_data_y_5__3__0_), .B1(npu_inst_pe_1_4_3_n2), .B2(
        npu_inst_int_data_x_4__4__0_), .ZN(npu_inst_pe_1_4_3_n61) );
  INV_X1 npu_inst_pe_1_4_3_U29 ( .A(npu_inst_pe_1_4_3_int_data_0_), .ZN(
        npu_inst_pe_1_4_3_n12) );
  INV_X1 npu_inst_pe_1_4_3_U28 ( .A(npu_inst_n51), .ZN(npu_inst_pe_1_4_3_n4)
         );
  OR3_X1 npu_inst_pe_1_4_3_U27 ( .A1(npu_inst_pe_1_4_3_n5), .A2(
        npu_inst_pe_1_4_3_n7), .A3(npu_inst_pe_1_4_3_n4), .ZN(
        npu_inst_pe_1_4_3_n56) );
  OR3_X1 npu_inst_pe_1_4_3_U26 ( .A1(npu_inst_pe_1_4_3_n4), .A2(
        npu_inst_pe_1_4_3_n7), .A3(npu_inst_pe_1_4_3_n6), .ZN(
        npu_inst_pe_1_4_3_n48) );
  INV_X1 npu_inst_pe_1_4_3_U25 ( .A(npu_inst_pe_1_4_3_n4), .ZN(
        npu_inst_pe_1_4_3_n3) );
  OR3_X1 npu_inst_pe_1_4_3_U24 ( .A1(npu_inst_pe_1_4_3_n3), .A2(
        npu_inst_pe_1_4_3_n7), .A3(npu_inst_pe_1_4_3_n6), .ZN(
        npu_inst_pe_1_4_3_n52) );
  OR3_X1 npu_inst_pe_1_4_3_U23 ( .A1(npu_inst_pe_1_4_3_n5), .A2(
        npu_inst_pe_1_4_3_n7), .A3(npu_inst_pe_1_4_3_n3), .ZN(
        npu_inst_pe_1_4_3_n60) );
  BUF_X1 npu_inst_pe_1_4_3_U22 ( .A(npu_inst_n20), .Z(npu_inst_pe_1_4_3_n1) );
  NOR2_X1 npu_inst_pe_1_4_3_U21 ( .A1(npu_inst_pe_1_4_3_n60), .A2(
        npu_inst_pe_1_4_3_n2), .ZN(npu_inst_pe_1_4_3_n58) );
  NOR2_X1 npu_inst_pe_1_4_3_U20 ( .A1(npu_inst_pe_1_4_3_n56), .A2(
        npu_inst_pe_1_4_3_n2), .ZN(npu_inst_pe_1_4_3_n54) );
  NOR2_X1 npu_inst_pe_1_4_3_U19 ( .A1(npu_inst_pe_1_4_3_n52), .A2(
        npu_inst_pe_1_4_3_n2), .ZN(npu_inst_pe_1_4_3_n50) );
  NOR2_X1 npu_inst_pe_1_4_3_U18 ( .A1(npu_inst_pe_1_4_3_n48), .A2(
        npu_inst_pe_1_4_3_n2), .ZN(npu_inst_pe_1_4_3_n46) );
  NOR2_X1 npu_inst_pe_1_4_3_U17 ( .A1(npu_inst_pe_1_4_3_n40), .A2(
        npu_inst_pe_1_4_3_n2), .ZN(npu_inst_pe_1_4_3_n38) );
  NOR2_X1 npu_inst_pe_1_4_3_U16 ( .A1(npu_inst_pe_1_4_3_n44), .A2(
        npu_inst_pe_1_4_3_n2), .ZN(npu_inst_pe_1_4_3_n42) );
  BUF_X1 npu_inst_pe_1_4_3_U15 ( .A(npu_inst_n81), .Z(npu_inst_pe_1_4_3_n7) );
  INV_X1 npu_inst_pe_1_4_3_U14 ( .A(npu_inst_n106), .ZN(npu_inst_pe_1_4_3_n11)
         );
  INV_X1 npu_inst_pe_1_4_3_U13 ( .A(npu_inst_pe_1_4_3_n38), .ZN(
        npu_inst_pe_1_4_3_n113) );
  INV_X1 npu_inst_pe_1_4_3_U12 ( .A(npu_inst_pe_1_4_3_n58), .ZN(
        npu_inst_pe_1_4_3_n118) );
  INV_X1 npu_inst_pe_1_4_3_U11 ( .A(npu_inst_pe_1_4_3_n54), .ZN(
        npu_inst_pe_1_4_3_n117) );
  INV_X1 npu_inst_pe_1_4_3_U10 ( .A(npu_inst_pe_1_4_3_n50), .ZN(
        npu_inst_pe_1_4_3_n116) );
  INV_X1 npu_inst_pe_1_4_3_U9 ( .A(npu_inst_pe_1_4_3_n46), .ZN(
        npu_inst_pe_1_4_3_n115) );
  INV_X1 npu_inst_pe_1_4_3_U8 ( .A(npu_inst_pe_1_4_3_n42), .ZN(
        npu_inst_pe_1_4_3_n114) );
  BUF_X1 npu_inst_pe_1_4_3_U7 ( .A(npu_inst_pe_1_4_3_n11), .Z(
        npu_inst_pe_1_4_3_n10) );
  BUF_X1 npu_inst_pe_1_4_3_U6 ( .A(npu_inst_pe_1_4_3_n11), .Z(
        npu_inst_pe_1_4_3_n9) );
  BUF_X1 npu_inst_pe_1_4_3_U5 ( .A(npu_inst_pe_1_4_3_n11), .Z(
        npu_inst_pe_1_4_3_n8) );
  NOR2_X1 npu_inst_pe_1_4_3_U4 ( .A1(npu_inst_pe_1_4_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_3_n1), .ZN(npu_inst_pe_1_4_3_n76) );
  NOR2_X1 npu_inst_pe_1_4_3_U3 ( .A1(npu_inst_pe_1_4_3_n27), .A2(
        npu_inst_pe_1_4_3_n1), .ZN(npu_inst_pe_1_4_3_n77) );
  FA_X1 npu_inst_pe_1_4_3_sub_77_U2_1 ( .A(npu_inst_int_data_res_4__3__1_), 
        .B(npu_inst_pe_1_4_3_n13), .CI(npu_inst_pe_1_4_3_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_4_3_sub_77_carry_2_), .S(npu_inst_pe_1_4_3_N66) );
  FA_X1 npu_inst_pe_1_4_3_add_79_U1_1 ( .A(npu_inst_int_data_res_4__3__1_), 
        .B(npu_inst_pe_1_4_3_int_data_1_), .CI(
        npu_inst_pe_1_4_3_add_79_carry_1_), .CO(
        npu_inst_pe_1_4_3_add_79_carry_2_), .S(npu_inst_pe_1_4_3_N74) );
  NAND3_X1 npu_inst_pe_1_4_3_U101 ( .A1(npu_inst_pe_1_4_3_n4), .A2(
        npu_inst_pe_1_4_3_n6), .A3(npu_inst_pe_1_4_3_n7), .ZN(
        npu_inst_pe_1_4_3_n44) );
  NAND3_X1 npu_inst_pe_1_4_3_U100 ( .A1(npu_inst_pe_1_4_3_n3), .A2(
        npu_inst_pe_1_4_3_n6), .A3(npu_inst_pe_1_4_3_n7), .ZN(
        npu_inst_pe_1_4_3_n40) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_3_n33), .CK(
        npu_inst_pe_1_4_3_net3673), .RN(npu_inst_pe_1_4_3_n8), .Q(
        npu_inst_int_data_res_4__3__6_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_3_n34), .CK(
        npu_inst_pe_1_4_3_net3673), .RN(npu_inst_pe_1_4_3_n8), .Q(
        npu_inst_int_data_res_4__3__5_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_3_n35), .CK(
        npu_inst_pe_1_4_3_net3673), .RN(npu_inst_pe_1_4_3_n8), .Q(
        npu_inst_int_data_res_4__3__4_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_3_n36), .CK(
        npu_inst_pe_1_4_3_net3673), .RN(npu_inst_pe_1_4_3_n8), .Q(
        npu_inst_int_data_res_4__3__3_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_3_n98), .CK(
        npu_inst_pe_1_4_3_net3673), .RN(npu_inst_pe_1_4_3_n8), .Q(
        npu_inst_int_data_res_4__3__2_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_3_n99), .CK(
        npu_inst_pe_1_4_3_net3673), .RN(npu_inst_pe_1_4_3_n8), .Q(
        npu_inst_int_data_res_4__3__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_3_n32), .CK(
        npu_inst_pe_1_4_3_net3673), .RN(npu_inst_pe_1_4_3_n8), .Q(
        npu_inst_int_data_res_4__3__7_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_3_n100), 
        .CK(npu_inst_pe_1_4_3_net3673), .RN(npu_inst_pe_1_4_3_n8), .Q(
        npu_inst_int_data_res_4__3__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_weight_reg_0_ ( .D(npu_inst_n92), .CK(
        npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n8), .Q(
        npu_inst_pe_1_4_3_int_q_weight_0_), .QN(npu_inst_pe_1_4_3_n27) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_weight_reg_1_ ( .D(npu_inst_n98), .CK(
        npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n8), .Q(
        npu_inst_pe_1_4_3_int_q_weight_1_), .QN(npu_inst_pe_1_4_3_n26) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_3_n112), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n8), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_3_n106), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n8), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_3_n111), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_3_n105), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_3_n110), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_3_n104), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_3_n109), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_3_n103), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_3_n108), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_3_n102), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_3_n107), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_3_n101), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_3_n86), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_3_n87), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n9), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_3_n88), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_3_n89), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_3_n90), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_3_n91), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_3_n92), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_3_n93), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_3_n94), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_3_n95), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_3_n96), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_3_n97), 
        .CK(npu_inst_pe_1_4_3_net3679), .RN(npu_inst_pe_1_4_3_n10), .Q(
        npu_inst_pe_1_4_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_3_net3673) );
  CLKGATETST_X1 npu_inst_pe_1_4_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n45), .SE(1'b0), .GCK(npu_inst_pe_1_4_3_net3679) );
  MUX2_X1 npu_inst_pe_1_4_4_U153 ( .A(npu_inst_pe_1_4_4_n31), .B(
        npu_inst_pe_1_4_4_n28), .S(npu_inst_pe_1_4_4_n7), .Z(
        npu_inst_pe_1_4_4_N93) );
  MUX2_X1 npu_inst_pe_1_4_4_U152 ( .A(npu_inst_pe_1_4_4_n30), .B(
        npu_inst_pe_1_4_4_n29), .S(npu_inst_pe_1_4_4_n5), .Z(
        npu_inst_pe_1_4_4_n31) );
  MUX2_X1 npu_inst_pe_1_4_4_U151 ( .A(npu_inst_pe_1_4_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_4_n3), .Z(
        npu_inst_pe_1_4_4_n30) );
  MUX2_X1 npu_inst_pe_1_4_4_U150 ( .A(npu_inst_pe_1_4_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_4_n3), .Z(
        npu_inst_pe_1_4_4_n29) );
  MUX2_X1 npu_inst_pe_1_4_4_U149 ( .A(npu_inst_pe_1_4_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_4_n3), .Z(
        npu_inst_pe_1_4_4_n28) );
  MUX2_X1 npu_inst_pe_1_4_4_U148 ( .A(npu_inst_pe_1_4_4_n25), .B(
        npu_inst_pe_1_4_4_n22), .S(npu_inst_pe_1_4_4_n7), .Z(
        npu_inst_pe_1_4_4_N94) );
  MUX2_X1 npu_inst_pe_1_4_4_U147 ( .A(npu_inst_pe_1_4_4_n24), .B(
        npu_inst_pe_1_4_4_n23), .S(npu_inst_pe_1_4_4_n5), .Z(
        npu_inst_pe_1_4_4_n25) );
  MUX2_X1 npu_inst_pe_1_4_4_U146 ( .A(npu_inst_pe_1_4_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_4_n3), .Z(
        npu_inst_pe_1_4_4_n24) );
  MUX2_X1 npu_inst_pe_1_4_4_U145 ( .A(npu_inst_pe_1_4_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_4_n3), .Z(
        npu_inst_pe_1_4_4_n23) );
  MUX2_X1 npu_inst_pe_1_4_4_U144 ( .A(npu_inst_pe_1_4_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_4_n3), .Z(
        npu_inst_pe_1_4_4_n22) );
  MUX2_X1 npu_inst_pe_1_4_4_U143 ( .A(npu_inst_pe_1_4_4_n21), .B(
        npu_inst_pe_1_4_4_n18), .S(npu_inst_pe_1_4_4_n7), .Z(
        npu_inst_int_data_x_4__4__1_) );
  MUX2_X1 npu_inst_pe_1_4_4_U142 ( .A(npu_inst_pe_1_4_4_n20), .B(
        npu_inst_pe_1_4_4_n19), .S(npu_inst_pe_1_4_4_n5), .Z(
        npu_inst_pe_1_4_4_n21) );
  MUX2_X1 npu_inst_pe_1_4_4_U141 ( .A(npu_inst_pe_1_4_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_4_n3), .Z(
        npu_inst_pe_1_4_4_n20) );
  MUX2_X1 npu_inst_pe_1_4_4_U140 ( .A(npu_inst_pe_1_4_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_4_n3), .Z(
        npu_inst_pe_1_4_4_n19) );
  MUX2_X1 npu_inst_pe_1_4_4_U139 ( .A(npu_inst_pe_1_4_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_4_n3), .Z(
        npu_inst_pe_1_4_4_n18) );
  MUX2_X1 npu_inst_pe_1_4_4_U138 ( .A(npu_inst_pe_1_4_4_n17), .B(
        npu_inst_pe_1_4_4_n14), .S(npu_inst_pe_1_4_4_n7), .Z(
        npu_inst_int_data_x_4__4__0_) );
  MUX2_X1 npu_inst_pe_1_4_4_U137 ( .A(npu_inst_pe_1_4_4_n16), .B(
        npu_inst_pe_1_4_4_n15), .S(npu_inst_pe_1_4_4_n5), .Z(
        npu_inst_pe_1_4_4_n17) );
  MUX2_X1 npu_inst_pe_1_4_4_U136 ( .A(npu_inst_pe_1_4_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_4_n3), .Z(
        npu_inst_pe_1_4_4_n16) );
  MUX2_X1 npu_inst_pe_1_4_4_U135 ( .A(npu_inst_pe_1_4_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_4_n3), .Z(
        npu_inst_pe_1_4_4_n15) );
  MUX2_X1 npu_inst_pe_1_4_4_U134 ( .A(npu_inst_pe_1_4_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_4_n3), .Z(
        npu_inst_pe_1_4_4_n14) );
  XOR2_X1 npu_inst_pe_1_4_4_U133 ( .A(npu_inst_pe_1_4_4_int_data_0_), .B(
        npu_inst_int_data_res_4__4__0_), .Z(npu_inst_pe_1_4_4_N73) );
  AND2_X1 npu_inst_pe_1_4_4_U132 ( .A1(npu_inst_int_data_res_4__4__0_), .A2(
        npu_inst_pe_1_4_4_int_data_0_), .ZN(npu_inst_pe_1_4_4_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_4_U131 ( .A(npu_inst_int_data_res_4__4__0_), .B(
        npu_inst_pe_1_4_4_n12), .ZN(npu_inst_pe_1_4_4_N65) );
  OR2_X1 npu_inst_pe_1_4_4_U130 ( .A1(npu_inst_pe_1_4_4_n12), .A2(
        npu_inst_int_data_res_4__4__0_), .ZN(npu_inst_pe_1_4_4_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_4_U129 ( .A(npu_inst_int_data_res_4__4__2_), .B(
        npu_inst_pe_1_4_4_add_79_carry_2_), .Z(npu_inst_pe_1_4_4_N75) );
  AND2_X1 npu_inst_pe_1_4_4_U128 ( .A1(npu_inst_pe_1_4_4_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_4__4__2_), .ZN(
        npu_inst_pe_1_4_4_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_4_U127 ( .A(npu_inst_int_data_res_4__4__3_), .B(
        npu_inst_pe_1_4_4_add_79_carry_3_), .Z(npu_inst_pe_1_4_4_N76) );
  AND2_X1 npu_inst_pe_1_4_4_U126 ( .A1(npu_inst_pe_1_4_4_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_4__4__3_), .ZN(
        npu_inst_pe_1_4_4_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_4_U125 ( .A(npu_inst_int_data_res_4__4__4_), .B(
        npu_inst_pe_1_4_4_add_79_carry_4_), .Z(npu_inst_pe_1_4_4_N77) );
  AND2_X1 npu_inst_pe_1_4_4_U124 ( .A1(npu_inst_pe_1_4_4_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_4__4__4_), .ZN(
        npu_inst_pe_1_4_4_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_4_U123 ( .A(npu_inst_int_data_res_4__4__5_), .B(
        npu_inst_pe_1_4_4_add_79_carry_5_), .Z(npu_inst_pe_1_4_4_N78) );
  AND2_X1 npu_inst_pe_1_4_4_U122 ( .A1(npu_inst_pe_1_4_4_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_4__4__5_), .ZN(
        npu_inst_pe_1_4_4_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_4_U121 ( .A(npu_inst_int_data_res_4__4__6_), .B(
        npu_inst_pe_1_4_4_add_79_carry_6_), .Z(npu_inst_pe_1_4_4_N79) );
  AND2_X1 npu_inst_pe_1_4_4_U120 ( .A1(npu_inst_pe_1_4_4_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_4__4__6_), .ZN(
        npu_inst_pe_1_4_4_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_4_U119 ( .A(npu_inst_int_data_res_4__4__7_), .B(
        npu_inst_pe_1_4_4_add_79_carry_7_), .Z(npu_inst_pe_1_4_4_N80) );
  XNOR2_X1 npu_inst_pe_1_4_4_U118 ( .A(npu_inst_pe_1_4_4_sub_77_carry_2_), .B(
        npu_inst_int_data_res_4__4__2_), .ZN(npu_inst_pe_1_4_4_N67) );
  OR2_X1 npu_inst_pe_1_4_4_U117 ( .A1(npu_inst_int_data_res_4__4__2_), .A2(
        npu_inst_pe_1_4_4_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_4_4_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_4_U116 ( .A(npu_inst_pe_1_4_4_sub_77_carry_3_), .B(
        npu_inst_int_data_res_4__4__3_), .ZN(npu_inst_pe_1_4_4_N68) );
  OR2_X1 npu_inst_pe_1_4_4_U115 ( .A1(npu_inst_int_data_res_4__4__3_), .A2(
        npu_inst_pe_1_4_4_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_4_4_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_4_U114 ( .A(npu_inst_pe_1_4_4_sub_77_carry_4_), .B(
        npu_inst_int_data_res_4__4__4_), .ZN(npu_inst_pe_1_4_4_N69) );
  OR2_X1 npu_inst_pe_1_4_4_U113 ( .A1(npu_inst_int_data_res_4__4__4_), .A2(
        npu_inst_pe_1_4_4_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_4_4_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_4_U112 ( .A(npu_inst_pe_1_4_4_sub_77_carry_5_), .B(
        npu_inst_int_data_res_4__4__5_), .ZN(npu_inst_pe_1_4_4_N70) );
  OR2_X1 npu_inst_pe_1_4_4_U111 ( .A1(npu_inst_int_data_res_4__4__5_), .A2(
        npu_inst_pe_1_4_4_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_4_4_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_4_U110 ( .A(npu_inst_pe_1_4_4_sub_77_carry_6_), .B(
        npu_inst_int_data_res_4__4__6_), .ZN(npu_inst_pe_1_4_4_N71) );
  OR2_X1 npu_inst_pe_1_4_4_U109 ( .A1(npu_inst_int_data_res_4__4__6_), .A2(
        npu_inst_pe_1_4_4_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_4_4_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_4_U108 ( .A(npu_inst_int_data_res_4__4__7_), .B(
        npu_inst_pe_1_4_4_sub_77_carry_7_), .ZN(npu_inst_pe_1_4_4_N72) );
  INV_X1 npu_inst_pe_1_4_4_U107 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_4_4_n6)
         );
  INV_X1 npu_inst_pe_1_4_4_U106 ( .A(npu_inst_pe_1_4_4_n6), .ZN(
        npu_inst_pe_1_4_4_n5) );
  INV_X1 npu_inst_pe_1_4_4_U105 ( .A(npu_inst_n37), .ZN(npu_inst_pe_1_4_4_n2)
         );
  AOI22_X1 npu_inst_pe_1_4_4_U104 ( .A1(npu_inst_int_data_y_5__4__0_), .A2(
        npu_inst_pe_1_4_4_n58), .B1(npu_inst_pe_1_4_4_n118), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_4_n57) );
  INV_X1 npu_inst_pe_1_4_4_U103 ( .A(npu_inst_pe_1_4_4_n57), .ZN(
        npu_inst_pe_1_4_4_n107) );
  AOI22_X1 npu_inst_pe_1_4_4_U102 ( .A1(npu_inst_int_data_y_5__4__0_), .A2(
        npu_inst_pe_1_4_4_n54), .B1(npu_inst_pe_1_4_4_n117), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_4_n53) );
  INV_X1 npu_inst_pe_1_4_4_U99 ( .A(npu_inst_pe_1_4_4_n53), .ZN(
        npu_inst_pe_1_4_4_n108) );
  AOI22_X1 npu_inst_pe_1_4_4_U98 ( .A1(npu_inst_int_data_y_5__4__0_), .A2(
        npu_inst_pe_1_4_4_n50), .B1(npu_inst_pe_1_4_4_n116), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_4_n49) );
  INV_X1 npu_inst_pe_1_4_4_U97 ( .A(npu_inst_pe_1_4_4_n49), .ZN(
        npu_inst_pe_1_4_4_n109) );
  AOI22_X1 npu_inst_pe_1_4_4_U96 ( .A1(npu_inst_int_data_y_5__4__0_), .A2(
        npu_inst_pe_1_4_4_n46), .B1(npu_inst_pe_1_4_4_n115), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_4_n45) );
  INV_X1 npu_inst_pe_1_4_4_U95 ( .A(npu_inst_pe_1_4_4_n45), .ZN(
        npu_inst_pe_1_4_4_n110) );
  AOI22_X1 npu_inst_pe_1_4_4_U94 ( .A1(npu_inst_int_data_y_5__4__0_), .A2(
        npu_inst_pe_1_4_4_n42), .B1(npu_inst_pe_1_4_4_n114), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_4_n41) );
  INV_X1 npu_inst_pe_1_4_4_U93 ( .A(npu_inst_pe_1_4_4_n41), .ZN(
        npu_inst_pe_1_4_4_n111) );
  AOI22_X1 npu_inst_pe_1_4_4_U92 ( .A1(npu_inst_int_data_y_5__4__1_), .A2(
        npu_inst_pe_1_4_4_n58), .B1(npu_inst_pe_1_4_4_n118), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_4_n59) );
  INV_X1 npu_inst_pe_1_4_4_U91 ( .A(npu_inst_pe_1_4_4_n59), .ZN(
        npu_inst_pe_1_4_4_n101) );
  AOI22_X1 npu_inst_pe_1_4_4_U90 ( .A1(npu_inst_int_data_y_5__4__1_), .A2(
        npu_inst_pe_1_4_4_n54), .B1(npu_inst_pe_1_4_4_n117), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_4_n55) );
  INV_X1 npu_inst_pe_1_4_4_U89 ( .A(npu_inst_pe_1_4_4_n55), .ZN(
        npu_inst_pe_1_4_4_n102) );
  AOI22_X1 npu_inst_pe_1_4_4_U88 ( .A1(npu_inst_int_data_y_5__4__1_), .A2(
        npu_inst_pe_1_4_4_n50), .B1(npu_inst_pe_1_4_4_n116), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_4_n51) );
  INV_X1 npu_inst_pe_1_4_4_U87 ( .A(npu_inst_pe_1_4_4_n51), .ZN(
        npu_inst_pe_1_4_4_n103) );
  AOI22_X1 npu_inst_pe_1_4_4_U86 ( .A1(npu_inst_int_data_y_5__4__1_), .A2(
        npu_inst_pe_1_4_4_n46), .B1(npu_inst_pe_1_4_4_n115), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_4_n47) );
  INV_X1 npu_inst_pe_1_4_4_U85 ( .A(npu_inst_pe_1_4_4_n47), .ZN(
        npu_inst_pe_1_4_4_n104) );
  AOI22_X1 npu_inst_pe_1_4_4_U84 ( .A1(npu_inst_int_data_y_5__4__1_), .A2(
        npu_inst_pe_1_4_4_n42), .B1(npu_inst_pe_1_4_4_n114), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_4_n43) );
  INV_X1 npu_inst_pe_1_4_4_U83 ( .A(npu_inst_pe_1_4_4_n43), .ZN(
        npu_inst_pe_1_4_4_n105) );
  AOI22_X1 npu_inst_pe_1_4_4_U82 ( .A1(npu_inst_pe_1_4_4_n38), .A2(
        npu_inst_int_data_y_5__4__1_), .B1(npu_inst_pe_1_4_4_n113), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_4_n39) );
  INV_X1 npu_inst_pe_1_4_4_U81 ( .A(npu_inst_pe_1_4_4_n39), .ZN(
        npu_inst_pe_1_4_4_n106) );
  NOR3_X1 npu_inst_pe_1_4_4_U80 ( .A1(npu_inst_pe_1_4_4_n26), .A2(npu_inst_n37), .A3(npu_inst_int_ckg[27]), .ZN(npu_inst_pe_1_4_4_n85) );
  OR2_X1 npu_inst_pe_1_4_4_U79 ( .A1(npu_inst_pe_1_4_4_n85), .A2(
        npu_inst_pe_1_4_4_n1), .ZN(npu_inst_pe_1_4_4_N84) );
  AND2_X1 npu_inst_pe_1_4_4_U78 ( .A1(npu_inst_pe_1_4_4_N93), .A2(npu_inst_n37), .ZN(npu_inst_int_data_y_4__4__0_) );
  NAND2_X1 npu_inst_pe_1_4_4_U77 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_4_n60), .ZN(npu_inst_pe_1_4_4_n74) );
  OAI21_X1 npu_inst_pe_1_4_4_U76 ( .B1(npu_inst_pe_1_4_4_n63), .B2(
        npu_inst_pe_1_4_4_n60), .A(npu_inst_pe_1_4_4_n74), .ZN(
        npu_inst_pe_1_4_4_n97) );
  NAND2_X1 npu_inst_pe_1_4_4_U75 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_4_n60), .ZN(npu_inst_pe_1_4_4_n73) );
  OAI21_X1 npu_inst_pe_1_4_4_U74 ( .B1(npu_inst_pe_1_4_4_n61), .B2(
        npu_inst_pe_1_4_4_n60), .A(npu_inst_pe_1_4_4_n73), .ZN(
        npu_inst_pe_1_4_4_n96) );
  NAND2_X1 npu_inst_pe_1_4_4_U73 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_4_n56), .ZN(npu_inst_pe_1_4_4_n72) );
  OAI21_X1 npu_inst_pe_1_4_4_U72 ( .B1(npu_inst_pe_1_4_4_n63), .B2(
        npu_inst_pe_1_4_4_n56), .A(npu_inst_pe_1_4_4_n72), .ZN(
        npu_inst_pe_1_4_4_n95) );
  NAND2_X1 npu_inst_pe_1_4_4_U71 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_4_n56), .ZN(npu_inst_pe_1_4_4_n71) );
  OAI21_X1 npu_inst_pe_1_4_4_U70 ( .B1(npu_inst_pe_1_4_4_n61), .B2(
        npu_inst_pe_1_4_4_n56), .A(npu_inst_pe_1_4_4_n71), .ZN(
        npu_inst_pe_1_4_4_n94) );
  NAND2_X1 npu_inst_pe_1_4_4_U69 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_4_n52), .ZN(npu_inst_pe_1_4_4_n70) );
  OAI21_X1 npu_inst_pe_1_4_4_U68 ( .B1(npu_inst_pe_1_4_4_n63), .B2(
        npu_inst_pe_1_4_4_n52), .A(npu_inst_pe_1_4_4_n70), .ZN(
        npu_inst_pe_1_4_4_n93) );
  NAND2_X1 npu_inst_pe_1_4_4_U67 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_4_n52), .ZN(npu_inst_pe_1_4_4_n69) );
  OAI21_X1 npu_inst_pe_1_4_4_U66 ( .B1(npu_inst_pe_1_4_4_n61), .B2(
        npu_inst_pe_1_4_4_n52), .A(npu_inst_pe_1_4_4_n69), .ZN(
        npu_inst_pe_1_4_4_n92) );
  NAND2_X1 npu_inst_pe_1_4_4_U65 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_4_n48), .ZN(npu_inst_pe_1_4_4_n68) );
  OAI21_X1 npu_inst_pe_1_4_4_U64 ( .B1(npu_inst_pe_1_4_4_n63), .B2(
        npu_inst_pe_1_4_4_n48), .A(npu_inst_pe_1_4_4_n68), .ZN(
        npu_inst_pe_1_4_4_n91) );
  NAND2_X1 npu_inst_pe_1_4_4_U63 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_4_n48), .ZN(npu_inst_pe_1_4_4_n67) );
  OAI21_X1 npu_inst_pe_1_4_4_U62 ( .B1(npu_inst_pe_1_4_4_n61), .B2(
        npu_inst_pe_1_4_4_n48), .A(npu_inst_pe_1_4_4_n67), .ZN(
        npu_inst_pe_1_4_4_n90) );
  NAND2_X1 npu_inst_pe_1_4_4_U61 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_4_n44), .ZN(npu_inst_pe_1_4_4_n66) );
  OAI21_X1 npu_inst_pe_1_4_4_U60 ( .B1(npu_inst_pe_1_4_4_n63), .B2(
        npu_inst_pe_1_4_4_n44), .A(npu_inst_pe_1_4_4_n66), .ZN(
        npu_inst_pe_1_4_4_n89) );
  NAND2_X1 npu_inst_pe_1_4_4_U59 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_4_n44), .ZN(npu_inst_pe_1_4_4_n65) );
  OAI21_X1 npu_inst_pe_1_4_4_U58 ( .B1(npu_inst_pe_1_4_4_n61), .B2(
        npu_inst_pe_1_4_4_n44), .A(npu_inst_pe_1_4_4_n65), .ZN(
        npu_inst_pe_1_4_4_n88) );
  NAND2_X1 npu_inst_pe_1_4_4_U57 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_4_n40), .ZN(npu_inst_pe_1_4_4_n64) );
  OAI21_X1 npu_inst_pe_1_4_4_U56 ( .B1(npu_inst_pe_1_4_4_n63), .B2(
        npu_inst_pe_1_4_4_n40), .A(npu_inst_pe_1_4_4_n64), .ZN(
        npu_inst_pe_1_4_4_n87) );
  NAND2_X1 npu_inst_pe_1_4_4_U55 ( .A1(npu_inst_pe_1_4_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_4_n40), .ZN(npu_inst_pe_1_4_4_n62) );
  OAI21_X1 npu_inst_pe_1_4_4_U54 ( .B1(npu_inst_pe_1_4_4_n61), .B2(
        npu_inst_pe_1_4_4_n40), .A(npu_inst_pe_1_4_4_n62), .ZN(
        npu_inst_pe_1_4_4_n86) );
  AOI22_X1 npu_inst_pe_1_4_4_U53 ( .A1(npu_inst_pe_1_4_4_n38), .A2(
        npu_inst_int_data_y_5__4__0_), .B1(npu_inst_pe_1_4_4_n113), .B2(
        npu_inst_pe_1_4_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_4_n37) );
  INV_X1 npu_inst_pe_1_4_4_U52 ( .A(npu_inst_pe_1_4_4_n37), .ZN(
        npu_inst_pe_1_4_4_n112) );
  AND2_X1 npu_inst_pe_1_4_4_U51 ( .A1(npu_inst_n37), .A2(npu_inst_pe_1_4_4_N94), .ZN(npu_inst_int_data_y_4__4__1_) );
  AOI222_X1 npu_inst_pe_1_4_4_U50 ( .A1(npu_inst_int_data_res_5__4__0_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N73), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N65), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n84) );
  INV_X1 npu_inst_pe_1_4_4_U49 ( .A(npu_inst_pe_1_4_4_n84), .ZN(
        npu_inst_pe_1_4_4_n100) );
  AOI222_X1 npu_inst_pe_1_4_4_U48 ( .A1(npu_inst_pe_1_4_4_n1), .A2(
        npu_inst_int_data_res_5__4__7_), .B1(npu_inst_pe_1_4_4_N80), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N72), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n75) );
  INV_X1 npu_inst_pe_1_4_4_U47 ( .A(npu_inst_pe_1_4_4_n75), .ZN(
        npu_inst_pe_1_4_4_n32) );
  AOI222_X1 npu_inst_pe_1_4_4_U46 ( .A1(npu_inst_int_data_res_5__4__1_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N74), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N66), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n83) );
  INV_X1 npu_inst_pe_1_4_4_U45 ( .A(npu_inst_pe_1_4_4_n83), .ZN(
        npu_inst_pe_1_4_4_n99) );
  AOI222_X1 npu_inst_pe_1_4_4_U44 ( .A1(npu_inst_int_data_res_5__4__3_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N76), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N68), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n81) );
  INV_X1 npu_inst_pe_1_4_4_U43 ( .A(npu_inst_pe_1_4_4_n81), .ZN(
        npu_inst_pe_1_4_4_n36) );
  AOI222_X1 npu_inst_pe_1_4_4_U42 ( .A1(npu_inst_int_data_res_5__4__4_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N77), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N69), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n80) );
  INV_X1 npu_inst_pe_1_4_4_U41 ( .A(npu_inst_pe_1_4_4_n80), .ZN(
        npu_inst_pe_1_4_4_n35) );
  AOI222_X1 npu_inst_pe_1_4_4_U40 ( .A1(npu_inst_int_data_res_5__4__5_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N78), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N70), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n79) );
  INV_X1 npu_inst_pe_1_4_4_U39 ( .A(npu_inst_pe_1_4_4_n79), .ZN(
        npu_inst_pe_1_4_4_n34) );
  AOI222_X1 npu_inst_pe_1_4_4_U38 ( .A1(npu_inst_int_data_res_5__4__6_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N79), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N71), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n78) );
  INV_X1 npu_inst_pe_1_4_4_U37 ( .A(npu_inst_pe_1_4_4_n78), .ZN(
        npu_inst_pe_1_4_4_n33) );
  AND2_X1 npu_inst_pe_1_4_4_U36 ( .A1(npu_inst_int_data_x_4__4__1_), .A2(
        npu_inst_pe_1_4_4_int_q_weight_1_), .ZN(npu_inst_pe_1_4_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_4_U35 ( .A1(npu_inst_int_data_x_4__4__0_), .A2(
        npu_inst_pe_1_4_4_int_q_weight_1_), .ZN(npu_inst_pe_1_4_4_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_4_4_U34 ( .A(npu_inst_pe_1_4_4_int_data_1_), .ZN(
        npu_inst_pe_1_4_4_n13) );
  AOI222_X1 npu_inst_pe_1_4_4_U33 ( .A1(npu_inst_int_data_res_5__4__2_), .A2(
        npu_inst_pe_1_4_4_n1), .B1(npu_inst_pe_1_4_4_N75), .B2(
        npu_inst_pe_1_4_4_n76), .C1(npu_inst_pe_1_4_4_N67), .C2(
        npu_inst_pe_1_4_4_n77), .ZN(npu_inst_pe_1_4_4_n82) );
  INV_X1 npu_inst_pe_1_4_4_U32 ( .A(npu_inst_pe_1_4_4_n82), .ZN(
        npu_inst_pe_1_4_4_n98) );
  AOI22_X1 npu_inst_pe_1_4_4_U31 ( .A1(npu_inst_n37), .A2(
        npu_inst_int_data_y_5__4__1_), .B1(npu_inst_pe_1_4_4_n2), .B2(
        npu_inst_int_data_x_4__5__1_), .ZN(npu_inst_pe_1_4_4_n63) );
  AOI22_X1 npu_inst_pe_1_4_4_U30 ( .A1(npu_inst_n37), .A2(
        npu_inst_int_data_y_5__4__0_), .B1(npu_inst_pe_1_4_4_n2), .B2(
        npu_inst_int_data_x_4__5__0_), .ZN(npu_inst_pe_1_4_4_n61) );
  INV_X1 npu_inst_pe_1_4_4_U29 ( .A(npu_inst_pe_1_4_4_int_data_0_), .ZN(
        npu_inst_pe_1_4_4_n12) );
  INV_X1 npu_inst_pe_1_4_4_U28 ( .A(npu_inst_n51), .ZN(npu_inst_pe_1_4_4_n4)
         );
  OR3_X1 npu_inst_pe_1_4_4_U27 ( .A1(npu_inst_pe_1_4_4_n5), .A2(
        npu_inst_pe_1_4_4_n7), .A3(npu_inst_pe_1_4_4_n4), .ZN(
        npu_inst_pe_1_4_4_n56) );
  OR3_X1 npu_inst_pe_1_4_4_U26 ( .A1(npu_inst_pe_1_4_4_n4), .A2(
        npu_inst_pe_1_4_4_n7), .A3(npu_inst_pe_1_4_4_n6), .ZN(
        npu_inst_pe_1_4_4_n48) );
  INV_X1 npu_inst_pe_1_4_4_U25 ( .A(npu_inst_pe_1_4_4_n4), .ZN(
        npu_inst_pe_1_4_4_n3) );
  OR3_X1 npu_inst_pe_1_4_4_U24 ( .A1(npu_inst_pe_1_4_4_n3), .A2(
        npu_inst_pe_1_4_4_n7), .A3(npu_inst_pe_1_4_4_n6), .ZN(
        npu_inst_pe_1_4_4_n52) );
  OR3_X1 npu_inst_pe_1_4_4_U23 ( .A1(npu_inst_pe_1_4_4_n5), .A2(
        npu_inst_pe_1_4_4_n7), .A3(npu_inst_pe_1_4_4_n3), .ZN(
        npu_inst_pe_1_4_4_n60) );
  BUF_X1 npu_inst_pe_1_4_4_U22 ( .A(npu_inst_n20), .Z(npu_inst_pe_1_4_4_n1) );
  NOR2_X1 npu_inst_pe_1_4_4_U21 ( .A1(npu_inst_pe_1_4_4_n60), .A2(
        npu_inst_pe_1_4_4_n2), .ZN(npu_inst_pe_1_4_4_n58) );
  NOR2_X1 npu_inst_pe_1_4_4_U20 ( .A1(npu_inst_pe_1_4_4_n56), .A2(
        npu_inst_pe_1_4_4_n2), .ZN(npu_inst_pe_1_4_4_n54) );
  NOR2_X1 npu_inst_pe_1_4_4_U19 ( .A1(npu_inst_pe_1_4_4_n52), .A2(
        npu_inst_pe_1_4_4_n2), .ZN(npu_inst_pe_1_4_4_n50) );
  NOR2_X1 npu_inst_pe_1_4_4_U18 ( .A1(npu_inst_pe_1_4_4_n48), .A2(
        npu_inst_pe_1_4_4_n2), .ZN(npu_inst_pe_1_4_4_n46) );
  NOR2_X1 npu_inst_pe_1_4_4_U17 ( .A1(npu_inst_pe_1_4_4_n40), .A2(
        npu_inst_pe_1_4_4_n2), .ZN(npu_inst_pe_1_4_4_n38) );
  NOR2_X1 npu_inst_pe_1_4_4_U16 ( .A1(npu_inst_pe_1_4_4_n44), .A2(
        npu_inst_pe_1_4_4_n2), .ZN(npu_inst_pe_1_4_4_n42) );
  BUF_X1 npu_inst_pe_1_4_4_U15 ( .A(npu_inst_n80), .Z(npu_inst_pe_1_4_4_n7) );
  INV_X1 npu_inst_pe_1_4_4_U14 ( .A(npu_inst_n106), .ZN(npu_inst_pe_1_4_4_n11)
         );
  INV_X1 npu_inst_pe_1_4_4_U13 ( .A(npu_inst_pe_1_4_4_n38), .ZN(
        npu_inst_pe_1_4_4_n113) );
  INV_X1 npu_inst_pe_1_4_4_U12 ( .A(npu_inst_pe_1_4_4_n58), .ZN(
        npu_inst_pe_1_4_4_n118) );
  INV_X1 npu_inst_pe_1_4_4_U11 ( .A(npu_inst_pe_1_4_4_n54), .ZN(
        npu_inst_pe_1_4_4_n117) );
  INV_X1 npu_inst_pe_1_4_4_U10 ( .A(npu_inst_pe_1_4_4_n50), .ZN(
        npu_inst_pe_1_4_4_n116) );
  INV_X1 npu_inst_pe_1_4_4_U9 ( .A(npu_inst_pe_1_4_4_n46), .ZN(
        npu_inst_pe_1_4_4_n115) );
  INV_X1 npu_inst_pe_1_4_4_U8 ( .A(npu_inst_pe_1_4_4_n42), .ZN(
        npu_inst_pe_1_4_4_n114) );
  BUF_X1 npu_inst_pe_1_4_4_U7 ( .A(npu_inst_pe_1_4_4_n11), .Z(
        npu_inst_pe_1_4_4_n10) );
  BUF_X1 npu_inst_pe_1_4_4_U6 ( .A(npu_inst_pe_1_4_4_n11), .Z(
        npu_inst_pe_1_4_4_n9) );
  BUF_X1 npu_inst_pe_1_4_4_U5 ( .A(npu_inst_pe_1_4_4_n11), .Z(
        npu_inst_pe_1_4_4_n8) );
  NOR2_X1 npu_inst_pe_1_4_4_U4 ( .A1(npu_inst_pe_1_4_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_4_n1), .ZN(npu_inst_pe_1_4_4_n76) );
  NOR2_X1 npu_inst_pe_1_4_4_U3 ( .A1(npu_inst_pe_1_4_4_n27), .A2(
        npu_inst_pe_1_4_4_n1), .ZN(npu_inst_pe_1_4_4_n77) );
  FA_X1 npu_inst_pe_1_4_4_sub_77_U2_1 ( .A(npu_inst_int_data_res_4__4__1_), 
        .B(npu_inst_pe_1_4_4_n13), .CI(npu_inst_pe_1_4_4_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_4_4_sub_77_carry_2_), .S(npu_inst_pe_1_4_4_N66) );
  FA_X1 npu_inst_pe_1_4_4_add_79_U1_1 ( .A(npu_inst_int_data_res_4__4__1_), 
        .B(npu_inst_pe_1_4_4_int_data_1_), .CI(
        npu_inst_pe_1_4_4_add_79_carry_1_), .CO(
        npu_inst_pe_1_4_4_add_79_carry_2_), .S(npu_inst_pe_1_4_4_N74) );
  NAND3_X1 npu_inst_pe_1_4_4_U101 ( .A1(npu_inst_pe_1_4_4_n4), .A2(
        npu_inst_pe_1_4_4_n6), .A3(npu_inst_pe_1_4_4_n7), .ZN(
        npu_inst_pe_1_4_4_n44) );
  NAND3_X1 npu_inst_pe_1_4_4_U100 ( .A1(npu_inst_pe_1_4_4_n3), .A2(
        npu_inst_pe_1_4_4_n6), .A3(npu_inst_pe_1_4_4_n7), .ZN(
        npu_inst_pe_1_4_4_n40) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_4_n33), .CK(
        npu_inst_pe_1_4_4_net3650), .RN(npu_inst_pe_1_4_4_n8), .Q(
        npu_inst_int_data_res_4__4__6_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_4_n34), .CK(
        npu_inst_pe_1_4_4_net3650), .RN(npu_inst_pe_1_4_4_n8), .Q(
        npu_inst_int_data_res_4__4__5_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_4_n35), .CK(
        npu_inst_pe_1_4_4_net3650), .RN(npu_inst_pe_1_4_4_n8), .Q(
        npu_inst_int_data_res_4__4__4_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_4_n36), .CK(
        npu_inst_pe_1_4_4_net3650), .RN(npu_inst_pe_1_4_4_n8), .Q(
        npu_inst_int_data_res_4__4__3_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_4_n98), .CK(
        npu_inst_pe_1_4_4_net3650), .RN(npu_inst_pe_1_4_4_n8), .Q(
        npu_inst_int_data_res_4__4__2_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_4_n99), .CK(
        npu_inst_pe_1_4_4_net3650), .RN(npu_inst_pe_1_4_4_n8), .Q(
        npu_inst_int_data_res_4__4__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_4_n32), .CK(
        npu_inst_pe_1_4_4_net3650), .RN(npu_inst_pe_1_4_4_n8), .Q(
        npu_inst_int_data_res_4__4__7_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_4_n100), 
        .CK(npu_inst_pe_1_4_4_net3650), .RN(npu_inst_pe_1_4_4_n8), .Q(
        npu_inst_int_data_res_4__4__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_weight_reg_0_ ( .D(npu_inst_n92), .CK(
        npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n8), .Q(
        npu_inst_pe_1_4_4_int_q_weight_0_), .QN(npu_inst_pe_1_4_4_n27) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_weight_reg_1_ ( .D(npu_inst_n98), .CK(
        npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n8), .Q(
        npu_inst_pe_1_4_4_int_q_weight_1_), .QN(npu_inst_pe_1_4_4_n26) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_4_n112), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n8), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_4_n106), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n8), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_4_n111), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_4_n105), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_4_n110), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_4_n104), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_4_n109), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_4_n103), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_4_n108), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_4_n102), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_4_n107), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_4_n101), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_4_n86), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_4_n87), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n9), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_4_n88), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_4_n89), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_4_n90), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_4_n91), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_4_n92), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_4_n93), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_4_n94), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_4_n95), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_4_n96), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_4_n97), 
        .CK(npu_inst_pe_1_4_4_net3656), .RN(npu_inst_pe_1_4_4_n10), .Q(
        npu_inst_pe_1_4_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_4_net3650) );
  CLKGATETST_X1 npu_inst_pe_1_4_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n45), .SE(1'b0), .GCK(npu_inst_pe_1_4_4_net3656) );
  MUX2_X1 npu_inst_pe_1_4_5_U153 ( .A(npu_inst_pe_1_4_5_n31), .B(
        npu_inst_pe_1_4_5_n28), .S(npu_inst_pe_1_4_5_n7), .Z(
        npu_inst_pe_1_4_5_N93) );
  MUX2_X1 npu_inst_pe_1_4_5_U152 ( .A(npu_inst_pe_1_4_5_n30), .B(
        npu_inst_pe_1_4_5_n29), .S(npu_inst_pe_1_4_5_n5), .Z(
        npu_inst_pe_1_4_5_n31) );
  MUX2_X1 npu_inst_pe_1_4_5_U151 ( .A(npu_inst_pe_1_4_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_5_n3), .Z(
        npu_inst_pe_1_4_5_n30) );
  MUX2_X1 npu_inst_pe_1_4_5_U150 ( .A(npu_inst_pe_1_4_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_5_n3), .Z(
        npu_inst_pe_1_4_5_n29) );
  MUX2_X1 npu_inst_pe_1_4_5_U149 ( .A(npu_inst_pe_1_4_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_5_n3), .Z(
        npu_inst_pe_1_4_5_n28) );
  MUX2_X1 npu_inst_pe_1_4_5_U148 ( .A(npu_inst_pe_1_4_5_n25), .B(
        npu_inst_pe_1_4_5_n22), .S(npu_inst_pe_1_4_5_n7), .Z(
        npu_inst_pe_1_4_5_N94) );
  MUX2_X1 npu_inst_pe_1_4_5_U147 ( .A(npu_inst_pe_1_4_5_n24), .B(
        npu_inst_pe_1_4_5_n23), .S(npu_inst_pe_1_4_5_n5), .Z(
        npu_inst_pe_1_4_5_n25) );
  MUX2_X1 npu_inst_pe_1_4_5_U146 ( .A(npu_inst_pe_1_4_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_5_n3), .Z(
        npu_inst_pe_1_4_5_n24) );
  MUX2_X1 npu_inst_pe_1_4_5_U145 ( .A(npu_inst_pe_1_4_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_5_n3), .Z(
        npu_inst_pe_1_4_5_n23) );
  MUX2_X1 npu_inst_pe_1_4_5_U144 ( .A(npu_inst_pe_1_4_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_5_n3), .Z(
        npu_inst_pe_1_4_5_n22) );
  MUX2_X1 npu_inst_pe_1_4_5_U143 ( .A(npu_inst_pe_1_4_5_n21), .B(
        npu_inst_pe_1_4_5_n18), .S(npu_inst_pe_1_4_5_n7), .Z(
        npu_inst_int_data_x_4__5__1_) );
  MUX2_X1 npu_inst_pe_1_4_5_U142 ( .A(npu_inst_pe_1_4_5_n20), .B(
        npu_inst_pe_1_4_5_n19), .S(npu_inst_pe_1_4_5_n5), .Z(
        npu_inst_pe_1_4_5_n21) );
  MUX2_X1 npu_inst_pe_1_4_5_U141 ( .A(npu_inst_pe_1_4_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_5_n3), .Z(
        npu_inst_pe_1_4_5_n20) );
  MUX2_X1 npu_inst_pe_1_4_5_U140 ( .A(npu_inst_pe_1_4_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_5_n3), .Z(
        npu_inst_pe_1_4_5_n19) );
  MUX2_X1 npu_inst_pe_1_4_5_U139 ( .A(npu_inst_pe_1_4_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_5_n3), .Z(
        npu_inst_pe_1_4_5_n18) );
  MUX2_X1 npu_inst_pe_1_4_5_U138 ( .A(npu_inst_pe_1_4_5_n17), .B(
        npu_inst_pe_1_4_5_n14), .S(npu_inst_pe_1_4_5_n7), .Z(
        npu_inst_int_data_x_4__5__0_) );
  MUX2_X1 npu_inst_pe_1_4_5_U137 ( .A(npu_inst_pe_1_4_5_n16), .B(
        npu_inst_pe_1_4_5_n15), .S(npu_inst_pe_1_4_5_n5), .Z(
        npu_inst_pe_1_4_5_n17) );
  MUX2_X1 npu_inst_pe_1_4_5_U136 ( .A(npu_inst_pe_1_4_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_5_n3), .Z(
        npu_inst_pe_1_4_5_n16) );
  MUX2_X1 npu_inst_pe_1_4_5_U135 ( .A(npu_inst_pe_1_4_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_5_n3), .Z(
        npu_inst_pe_1_4_5_n15) );
  MUX2_X1 npu_inst_pe_1_4_5_U134 ( .A(npu_inst_pe_1_4_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_5_n3), .Z(
        npu_inst_pe_1_4_5_n14) );
  XOR2_X1 npu_inst_pe_1_4_5_U133 ( .A(npu_inst_pe_1_4_5_int_data_0_), .B(
        npu_inst_int_data_res_4__5__0_), .Z(npu_inst_pe_1_4_5_N73) );
  AND2_X1 npu_inst_pe_1_4_5_U132 ( .A1(npu_inst_int_data_res_4__5__0_), .A2(
        npu_inst_pe_1_4_5_int_data_0_), .ZN(npu_inst_pe_1_4_5_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_5_U131 ( .A(npu_inst_int_data_res_4__5__0_), .B(
        npu_inst_pe_1_4_5_n12), .ZN(npu_inst_pe_1_4_5_N65) );
  OR2_X1 npu_inst_pe_1_4_5_U130 ( .A1(npu_inst_pe_1_4_5_n12), .A2(
        npu_inst_int_data_res_4__5__0_), .ZN(npu_inst_pe_1_4_5_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_5_U129 ( .A(npu_inst_int_data_res_4__5__2_), .B(
        npu_inst_pe_1_4_5_add_79_carry_2_), .Z(npu_inst_pe_1_4_5_N75) );
  AND2_X1 npu_inst_pe_1_4_5_U128 ( .A1(npu_inst_pe_1_4_5_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_4__5__2_), .ZN(
        npu_inst_pe_1_4_5_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_5_U127 ( .A(npu_inst_int_data_res_4__5__3_), .B(
        npu_inst_pe_1_4_5_add_79_carry_3_), .Z(npu_inst_pe_1_4_5_N76) );
  AND2_X1 npu_inst_pe_1_4_5_U126 ( .A1(npu_inst_pe_1_4_5_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_4__5__3_), .ZN(
        npu_inst_pe_1_4_5_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_5_U125 ( .A(npu_inst_int_data_res_4__5__4_), .B(
        npu_inst_pe_1_4_5_add_79_carry_4_), .Z(npu_inst_pe_1_4_5_N77) );
  AND2_X1 npu_inst_pe_1_4_5_U124 ( .A1(npu_inst_pe_1_4_5_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_4__5__4_), .ZN(
        npu_inst_pe_1_4_5_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_5_U123 ( .A(npu_inst_int_data_res_4__5__5_), .B(
        npu_inst_pe_1_4_5_add_79_carry_5_), .Z(npu_inst_pe_1_4_5_N78) );
  AND2_X1 npu_inst_pe_1_4_5_U122 ( .A1(npu_inst_pe_1_4_5_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_4__5__5_), .ZN(
        npu_inst_pe_1_4_5_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_5_U121 ( .A(npu_inst_int_data_res_4__5__6_), .B(
        npu_inst_pe_1_4_5_add_79_carry_6_), .Z(npu_inst_pe_1_4_5_N79) );
  AND2_X1 npu_inst_pe_1_4_5_U120 ( .A1(npu_inst_pe_1_4_5_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_4__5__6_), .ZN(
        npu_inst_pe_1_4_5_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_5_U119 ( .A(npu_inst_int_data_res_4__5__7_), .B(
        npu_inst_pe_1_4_5_add_79_carry_7_), .Z(npu_inst_pe_1_4_5_N80) );
  XNOR2_X1 npu_inst_pe_1_4_5_U118 ( .A(npu_inst_pe_1_4_5_sub_77_carry_2_), .B(
        npu_inst_int_data_res_4__5__2_), .ZN(npu_inst_pe_1_4_5_N67) );
  OR2_X1 npu_inst_pe_1_4_5_U117 ( .A1(npu_inst_int_data_res_4__5__2_), .A2(
        npu_inst_pe_1_4_5_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_4_5_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_5_U116 ( .A(npu_inst_pe_1_4_5_sub_77_carry_3_), .B(
        npu_inst_int_data_res_4__5__3_), .ZN(npu_inst_pe_1_4_5_N68) );
  OR2_X1 npu_inst_pe_1_4_5_U115 ( .A1(npu_inst_int_data_res_4__5__3_), .A2(
        npu_inst_pe_1_4_5_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_4_5_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_5_U114 ( .A(npu_inst_pe_1_4_5_sub_77_carry_4_), .B(
        npu_inst_int_data_res_4__5__4_), .ZN(npu_inst_pe_1_4_5_N69) );
  OR2_X1 npu_inst_pe_1_4_5_U113 ( .A1(npu_inst_int_data_res_4__5__4_), .A2(
        npu_inst_pe_1_4_5_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_4_5_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_5_U112 ( .A(npu_inst_pe_1_4_5_sub_77_carry_5_), .B(
        npu_inst_int_data_res_4__5__5_), .ZN(npu_inst_pe_1_4_5_N70) );
  OR2_X1 npu_inst_pe_1_4_5_U111 ( .A1(npu_inst_int_data_res_4__5__5_), .A2(
        npu_inst_pe_1_4_5_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_4_5_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_5_U110 ( .A(npu_inst_pe_1_4_5_sub_77_carry_6_), .B(
        npu_inst_int_data_res_4__5__6_), .ZN(npu_inst_pe_1_4_5_N71) );
  OR2_X1 npu_inst_pe_1_4_5_U109 ( .A1(npu_inst_int_data_res_4__5__6_), .A2(
        npu_inst_pe_1_4_5_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_4_5_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_5_U108 ( .A(npu_inst_int_data_res_4__5__7_), .B(
        npu_inst_pe_1_4_5_sub_77_carry_7_), .ZN(npu_inst_pe_1_4_5_N72) );
  INV_X1 npu_inst_pe_1_4_5_U107 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_4_5_n6)
         );
  INV_X1 npu_inst_pe_1_4_5_U106 ( .A(npu_inst_pe_1_4_5_n6), .ZN(
        npu_inst_pe_1_4_5_n5) );
  INV_X1 npu_inst_pe_1_4_5_U105 ( .A(npu_inst_n37), .ZN(npu_inst_pe_1_4_5_n2)
         );
  AOI22_X1 npu_inst_pe_1_4_5_U104 ( .A1(npu_inst_int_data_y_5__5__0_), .A2(
        npu_inst_pe_1_4_5_n58), .B1(npu_inst_pe_1_4_5_n118), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_5_n57) );
  INV_X1 npu_inst_pe_1_4_5_U103 ( .A(npu_inst_pe_1_4_5_n57), .ZN(
        npu_inst_pe_1_4_5_n107) );
  AOI22_X1 npu_inst_pe_1_4_5_U102 ( .A1(npu_inst_int_data_y_5__5__0_), .A2(
        npu_inst_pe_1_4_5_n54), .B1(npu_inst_pe_1_4_5_n117), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_5_n53) );
  INV_X1 npu_inst_pe_1_4_5_U99 ( .A(npu_inst_pe_1_4_5_n53), .ZN(
        npu_inst_pe_1_4_5_n108) );
  AOI22_X1 npu_inst_pe_1_4_5_U98 ( .A1(npu_inst_int_data_y_5__5__0_), .A2(
        npu_inst_pe_1_4_5_n50), .B1(npu_inst_pe_1_4_5_n116), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_5_n49) );
  INV_X1 npu_inst_pe_1_4_5_U97 ( .A(npu_inst_pe_1_4_5_n49), .ZN(
        npu_inst_pe_1_4_5_n109) );
  AOI22_X1 npu_inst_pe_1_4_5_U96 ( .A1(npu_inst_int_data_y_5__5__0_), .A2(
        npu_inst_pe_1_4_5_n46), .B1(npu_inst_pe_1_4_5_n115), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_5_n45) );
  INV_X1 npu_inst_pe_1_4_5_U95 ( .A(npu_inst_pe_1_4_5_n45), .ZN(
        npu_inst_pe_1_4_5_n110) );
  AOI22_X1 npu_inst_pe_1_4_5_U94 ( .A1(npu_inst_int_data_y_5__5__0_), .A2(
        npu_inst_pe_1_4_5_n42), .B1(npu_inst_pe_1_4_5_n114), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_5_n41) );
  INV_X1 npu_inst_pe_1_4_5_U93 ( .A(npu_inst_pe_1_4_5_n41), .ZN(
        npu_inst_pe_1_4_5_n111) );
  AOI22_X1 npu_inst_pe_1_4_5_U92 ( .A1(npu_inst_int_data_y_5__5__1_), .A2(
        npu_inst_pe_1_4_5_n58), .B1(npu_inst_pe_1_4_5_n118), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_5_n59) );
  INV_X1 npu_inst_pe_1_4_5_U91 ( .A(npu_inst_pe_1_4_5_n59), .ZN(
        npu_inst_pe_1_4_5_n101) );
  AOI22_X1 npu_inst_pe_1_4_5_U90 ( .A1(npu_inst_int_data_y_5__5__1_), .A2(
        npu_inst_pe_1_4_5_n54), .B1(npu_inst_pe_1_4_5_n117), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_5_n55) );
  INV_X1 npu_inst_pe_1_4_5_U89 ( .A(npu_inst_pe_1_4_5_n55), .ZN(
        npu_inst_pe_1_4_5_n102) );
  AOI22_X1 npu_inst_pe_1_4_5_U88 ( .A1(npu_inst_int_data_y_5__5__1_), .A2(
        npu_inst_pe_1_4_5_n50), .B1(npu_inst_pe_1_4_5_n116), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_5_n51) );
  INV_X1 npu_inst_pe_1_4_5_U87 ( .A(npu_inst_pe_1_4_5_n51), .ZN(
        npu_inst_pe_1_4_5_n103) );
  AOI22_X1 npu_inst_pe_1_4_5_U86 ( .A1(npu_inst_int_data_y_5__5__1_), .A2(
        npu_inst_pe_1_4_5_n46), .B1(npu_inst_pe_1_4_5_n115), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_5_n47) );
  INV_X1 npu_inst_pe_1_4_5_U85 ( .A(npu_inst_pe_1_4_5_n47), .ZN(
        npu_inst_pe_1_4_5_n104) );
  AOI22_X1 npu_inst_pe_1_4_5_U84 ( .A1(npu_inst_int_data_y_5__5__1_), .A2(
        npu_inst_pe_1_4_5_n42), .B1(npu_inst_pe_1_4_5_n114), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_5_n43) );
  INV_X1 npu_inst_pe_1_4_5_U83 ( .A(npu_inst_pe_1_4_5_n43), .ZN(
        npu_inst_pe_1_4_5_n105) );
  AOI22_X1 npu_inst_pe_1_4_5_U82 ( .A1(npu_inst_pe_1_4_5_n38), .A2(
        npu_inst_int_data_y_5__5__1_), .B1(npu_inst_pe_1_4_5_n113), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_5_n39) );
  INV_X1 npu_inst_pe_1_4_5_U81 ( .A(npu_inst_pe_1_4_5_n39), .ZN(
        npu_inst_pe_1_4_5_n106) );
  AND2_X1 npu_inst_pe_1_4_5_U80 ( .A1(npu_inst_pe_1_4_5_N93), .A2(npu_inst_n37), .ZN(npu_inst_int_data_y_4__5__0_) );
  NAND2_X1 npu_inst_pe_1_4_5_U79 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_5_n60), .ZN(npu_inst_pe_1_4_5_n74) );
  OAI21_X1 npu_inst_pe_1_4_5_U78 ( .B1(npu_inst_pe_1_4_5_n63), .B2(
        npu_inst_pe_1_4_5_n60), .A(npu_inst_pe_1_4_5_n74), .ZN(
        npu_inst_pe_1_4_5_n97) );
  NAND2_X1 npu_inst_pe_1_4_5_U77 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_5_n60), .ZN(npu_inst_pe_1_4_5_n73) );
  OAI21_X1 npu_inst_pe_1_4_5_U76 ( .B1(npu_inst_pe_1_4_5_n61), .B2(
        npu_inst_pe_1_4_5_n60), .A(npu_inst_pe_1_4_5_n73), .ZN(
        npu_inst_pe_1_4_5_n96) );
  NAND2_X1 npu_inst_pe_1_4_5_U75 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_5_n56), .ZN(npu_inst_pe_1_4_5_n72) );
  OAI21_X1 npu_inst_pe_1_4_5_U74 ( .B1(npu_inst_pe_1_4_5_n63), .B2(
        npu_inst_pe_1_4_5_n56), .A(npu_inst_pe_1_4_5_n72), .ZN(
        npu_inst_pe_1_4_5_n95) );
  NAND2_X1 npu_inst_pe_1_4_5_U73 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_5_n56), .ZN(npu_inst_pe_1_4_5_n71) );
  OAI21_X1 npu_inst_pe_1_4_5_U72 ( .B1(npu_inst_pe_1_4_5_n61), .B2(
        npu_inst_pe_1_4_5_n56), .A(npu_inst_pe_1_4_5_n71), .ZN(
        npu_inst_pe_1_4_5_n94) );
  NAND2_X1 npu_inst_pe_1_4_5_U71 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_5_n52), .ZN(npu_inst_pe_1_4_5_n70) );
  OAI21_X1 npu_inst_pe_1_4_5_U70 ( .B1(npu_inst_pe_1_4_5_n63), .B2(
        npu_inst_pe_1_4_5_n52), .A(npu_inst_pe_1_4_5_n70), .ZN(
        npu_inst_pe_1_4_5_n93) );
  NAND2_X1 npu_inst_pe_1_4_5_U69 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_5_n52), .ZN(npu_inst_pe_1_4_5_n69) );
  OAI21_X1 npu_inst_pe_1_4_5_U68 ( .B1(npu_inst_pe_1_4_5_n61), .B2(
        npu_inst_pe_1_4_5_n52), .A(npu_inst_pe_1_4_5_n69), .ZN(
        npu_inst_pe_1_4_5_n92) );
  NAND2_X1 npu_inst_pe_1_4_5_U67 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_5_n48), .ZN(npu_inst_pe_1_4_5_n68) );
  OAI21_X1 npu_inst_pe_1_4_5_U66 ( .B1(npu_inst_pe_1_4_5_n63), .B2(
        npu_inst_pe_1_4_5_n48), .A(npu_inst_pe_1_4_5_n68), .ZN(
        npu_inst_pe_1_4_5_n91) );
  NAND2_X1 npu_inst_pe_1_4_5_U65 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_5_n48), .ZN(npu_inst_pe_1_4_5_n67) );
  OAI21_X1 npu_inst_pe_1_4_5_U64 ( .B1(npu_inst_pe_1_4_5_n61), .B2(
        npu_inst_pe_1_4_5_n48), .A(npu_inst_pe_1_4_5_n67), .ZN(
        npu_inst_pe_1_4_5_n90) );
  NAND2_X1 npu_inst_pe_1_4_5_U63 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_5_n44), .ZN(npu_inst_pe_1_4_5_n66) );
  OAI21_X1 npu_inst_pe_1_4_5_U62 ( .B1(npu_inst_pe_1_4_5_n63), .B2(
        npu_inst_pe_1_4_5_n44), .A(npu_inst_pe_1_4_5_n66), .ZN(
        npu_inst_pe_1_4_5_n89) );
  NAND2_X1 npu_inst_pe_1_4_5_U61 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_5_n44), .ZN(npu_inst_pe_1_4_5_n65) );
  OAI21_X1 npu_inst_pe_1_4_5_U60 ( .B1(npu_inst_pe_1_4_5_n61), .B2(
        npu_inst_pe_1_4_5_n44), .A(npu_inst_pe_1_4_5_n65), .ZN(
        npu_inst_pe_1_4_5_n88) );
  NAND2_X1 npu_inst_pe_1_4_5_U59 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_5_n40), .ZN(npu_inst_pe_1_4_5_n64) );
  OAI21_X1 npu_inst_pe_1_4_5_U58 ( .B1(npu_inst_pe_1_4_5_n63), .B2(
        npu_inst_pe_1_4_5_n40), .A(npu_inst_pe_1_4_5_n64), .ZN(
        npu_inst_pe_1_4_5_n87) );
  NAND2_X1 npu_inst_pe_1_4_5_U57 ( .A1(npu_inst_pe_1_4_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_5_n40), .ZN(npu_inst_pe_1_4_5_n62) );
  OAI21_X1 npu_inst_pe_1_4_5_U56 ( .B1(npu_inst_pe_1_4_5_n61), .B2(
        npu_inst_pe_1_4_5_n40), .A(npu_inst_pe_1_4_5_n62), .ZN(
        npu_inst_pe_1_4_5_n86) );
  AOI22_X1 npu_inst_pe_1_4_5_U55 ( .A1(npu_inst_pe_1_4_5_n38), .A2(
        npu_inst_int_data_y_5__5__0_), .B1(npu_inst_pe_1_4_5_n113), .B2(
        npu_inst_pe_1_4_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_5_n37) );
  INV_X1 npu_inst_pe_1_4_5_U54 ( .A(npu_inst_pe_1_4_5_n37), .ZN(
        npu_inst_pe_1_4_5_n112) );
  AND2_X1 npu_inst_pe_1_4_5_U53 ( .A1(npu_inst_n37), .A2(npu_inst_pe_1_4_5_N94), .ZN(npu_inst_int_data_y_4__5__1_) );
  AOI222_X1 npu_inst_pe_1_4_5_U52 ( .A1(npu_inst_int_data_res_5__5__0_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N73), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N65), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n84) );
  INV_X1 npu_inst_pe_1_4_5_U51 ( .A(npu_inst_pe_1_4_5_n84), .ZN(
        npu_inst_pe_1_4_5_n100) );
  AOI222_X1 npu_inst_pe_1_4_5_U50 ( .A1(npu_inst_pe_1_4_5_n1), .A2(
        npu_inst_int_data_res_5__5__7_), .B1(npu_inst_pe_1_4_5_N80), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N72), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n75) );
  INV_X1 npu_inst_pe_1_4_5_U49 ( .A(npu_inst_pe_1_4_5_n75), .ZN(
        npu_inst_pe_1_4_5_n32) );
  AOI222_X1 npu_inst_pe_1_4_5_U48 ( .A1(npu_inst_int_data_res_5__5__1_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N74), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N66), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n83) );
  INV_X1 npu_inst_pe_1_4_5_U47 ( .A(npu_inst_pe_1_4_5_n83), .ZN(
        npu_inst_pe_1_4_5_n99) );
  AOI222_X1 npu_inst_pe_1_4_5_U46 ( .A1(npu_inst_int_data_res_5__5__3_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N76), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N68), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n81) );
  INV_X1 npu_inst_pe_1_4_5_U45 ( .A(npu_inst_pe_1_4_5_n81), .ZN(
        npu_inst_pe_1_4_5_n36) );
  AOI222_X1 npu_inst_pe_1_4_5_U44 ( .A1(npu_inst_int_data_res_5__5__4_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N77), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N69), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n80) );
  INV_X1 npu_inst_pe_1_4_5_U43 ( .A(npu_inst_pe_1_4_5_n80), .ZN(
        npu_inst_pe_1_4_5_n35) );
  AOI222_X1 npu_inst_pe_1_4_5_U42 ( .A1(npu_inst_int_data_res_5__5__5_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N78), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N70), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n79) );
  INV_X1 npu_inst_pe_1_4_5_U41 ( .A(npu_inst_pe_1_4_5_n79), .ZN(
        npu_inst_pe_1_4_5_n34) );
  AOI222_X1 npu_inst_pe_1_4_5_U40 ( .A1(npu_inst_int_data_res_5__5__6_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N79), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N71), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n78) );
  INV_X1 npu_inst_pe_1_4_5_U39 ( .A(npu_inst_pe_1_4_5_n78), .ZN(
        npu_inst_pe_1_4_5_n33) );
  AND2_X1 npu_inst_pe_1_4_5_U38 ( .A1(npu_inst_int_data_x_4__5__1_), .A2(
        npu_inst_pe_1_4_5_int_q_weight_1_), .ZN(npu_inst_pe_1_4_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_5_U37 ( .A1(npu_inst_int_data_x_4__5__0_), .A2(
        npu_inst_pe_1_4_5_int_q_weight_1_), .ZN(npu_inst_pe_1_4_5_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_4_5_U36 ( .A(npu_inst_pe_1_4_5_int_data_1_), .ZN(
        npu_inst_pe_1_4_5_n13) );
  NOR3_X1 npu_inst_pe_1_4_5_U35 ( .A1(npu_inst_pe_1_4_5_n26), .A2(npu_inst_n37), .A3(npu_inst_int_ckg[26]), .ZN(npu_inst_pe_1_4_5_n85) );
  OR2_X1 npu_inst_pe_1_4_5_U34 ( .A1(npu_inst_pe_1_4_5_n85), .A2(
        npu_inst_pe_1_4_5_n1), .ZN(npu_inst_pe_1_4_5_N84) );
  AOI222_X1 npu_inst_pe_1_4_5_U33 ( .A1(npu_inst_int_data_res_5__5__2_), .A2(
        npu_inst_pe_1_4_5_n1), .B1(npu_inst_pe_1_4_5_N75), .B2(
        npu_inst_pe_1_4_5_n76), .C1(npu_inst_pe_1_4_5_N67), .C2(
        npu_inst_pe_1_4_5_n77), .ZN(npu_inst_pe_1_4_5_n82) );
  INV_X1 npu_inst_pe_1_4_5_U32 ( .A(npu_inst_pe_1_4_5_n82), .ZN(
        npu_inst_pe_1_4_5_n98) );
  AOI22_X1 npu_inst_pe_1_4_5_U31 ( .A1(npu_inst_n37), .A2(
        npu_inst_int_data_y_5__5__1_), .B1(npu_inst_pe_1_4_5_n2), .B2(
        npu_inst_int_data_x_4__6__1_), .ZN(npu_inst_pe_1_4_5_n63) );
  AOI22_X1 npu_inst_pe_1_4_5_U30 ( .A1(npu_inst_n37), .A2(
        npu_inst_int_data_y_5__5__0_), .B1(npu_inst_pe_1_4_5_n2), .B2(
        npu_inst_int_data_x_4__6__0_), .ZN(npu_inst_pe_1_4_5_n61) );
  INV_X1 npu_inst_pe_1_4_5_U29 ( .A(npu_inst_pe_1_4_5_int_data_0_), .ZN(
        npu_inst_pe_1_4_5_n12) );
  INV_X1 npu_inst_pe_1_4_5_U28 ( .A(npu_inst_n51), .ZN(npu_inst_pe_1_4_5_n4)
         );
  OR3_X1 npu_inst_pe_1_4_5_U27 ( .A1(npu_inst_pe_1_4_5_n5), .A2(
        npu_inst_pe_1_4_5_n7), .A3(npu_inst_pe_1_4_5_n4), .ZN(
        npu_inst_pe_1_4_5_n56) );
  OR3_X1 npu_inst_pe_1_4_5_U26 ( .A1(npu_inst_pe_1_4_5_n4), .A2(
        npu_inst_pe_1_4_5_n7), .A3(npu_inst_pe_1_4_5_n6), .ZN(
        npu_inst_pe_1_4_5_n48) );
  INV_X1 npu_inst_pe_1_4_5_U25 ( .A(npu_inst_pe_1_4_5_n4), .ZN(
        npu_inst_pe_1_4_5_n3) );
  OR3_X1 npu_inst_pe_1_4_5_U24 ( .A1(npu_inst_pe_1_4_5_n3), .A2(
        npu_inst_pe_1_4_5_n7), .A3(npu_inst_pe_1_4_5_n6), .ZN(
        npu_inst_pe_1_4_5_n52) );
  OR3_X1 npu_inst_pe_1_4_5_U23 ( .A1(npu_inst_pe_1_4_5_n5), .A2(
        npu_inst_pe_1_4_5_n7), .A3(npu_inst_pe_1_4_5_n3), .ZN(
        npu_inst_pe_1_4_5_n60) );
  BUF_X1 npu_inst_pe_1_4_5_U22 ( .A(npu_inst_n19), .Z(npu_inst_pe_1_4_5_n1) );
  NOR2_X1 npu_inst_pe_1_4_5_U21 ( .A1(npu_inst_pe_1_4_5_n60), .A2(
        npu_inst_pe_1_4_5_n2), .ZN(npu_inst_pe_1_4_5_n58) );
  NOR2_X1 npu_inst_pe_1_4_5_U20 ( .A1(npu_inst_pe_1_4_5_n56), .A2(
        npu_inst_pe_1_4_5_n2), .ZN(npu_inst_pe_1_4_5_n54) );
  NOR2_X1 npu_inst_pe_1_4_5_U19 ( .A1(npu_inst_pe_1_4_5_n52), .A2(
        npu_inst_pe_1_4_5_n2), .ZN(npu_inst_pe_1_4_5_n50) );
  NOR2_X1 npu_inst_pe_1_4_5_U18 ( .A1(npu_inst_pe_1_4_5_n48), .A2(
        npu_inst_pe_1_4_5_n2), .ZN(npu_inst_pe_1_4_5_n46) );
  NOR2_X1 npu_inst_pe_1_4_5_U17 ( .A1(npu_inst_pe_1_4_5_n40), .A2(
        npu_inst_pe_1_4_5_n2), .ZN(npu_inst_pe_1_4_5_n38) );
  NOR2_X1 npu_inst_pe_1_4_5_U16 ( .A1(npu_inst_pe_1_4_5_n44), .A2(
        npu_inst_pe_1_4_5_n2), .ZN(npu_inst_pe_1_4_5_n42) );
  BUF_X1 npu_inst_pe_1_4_5_U15 ( .A(npu_inst_n80), .Z(npu_inst_pe_1_4_5_n7) );
  INV_X1 npu_inst_pe_1_4_5_U14 ( .A(npu_inst_n106), .ZN(npu_inst_pe_1_4_5_n11)
         );
  INV_X1 npu_inst_pe_1_4_5_U13 ( .A(npu_inst_pe_1_4_5_n38), .ZN(
        npu_inst_pe_1_4_5_n113) );
  INV_X1 npu_inst_pe_1_4_5_U12 ( .A(npu_inst_pe_1_4_5_n58), .ZN(
        npu_inst_pe_1_4_5_n118) );
  INV_X1 npu_inst_pe_1_4_5_U11 ( .A(npu_inst_pe_1_4_5_n54), .ZN(
        npu_inst_pe_1_4_5_n117) );
  INV_X1 npu_inst_pe_1_4_5_U10 ( .A(npu_inst_pe_1_4_5_n50), .ZN(
        npu_inst_pe_1_4_5_n116) );
  INV_X1 npu_inst_pe_1_4_5_U9 ( .A(npu_inst_pe_1_4_5_n46), .ZN(
        npu_inst_pe_1_4_5_n115) );
  INV_X1 npu_inst_pe_1_4_5_U8 ( .A(npu_inst_pe_1_4_5_n42), .ZN(
        npu_inst_pe_1_4_5_n114) );
  BUF_X1 npu_inst_pe_1_4_5_U7 ( .A(npu_inst_pe_1_4_5_n11), .Z(
        npu_inst_pe_1_4_5_n10) );
  BUF_X1 npu_inst_pe_1_4_5_U6 ( .A(npu_inst_pe_1_4_5_n11), .Z(
        npu_inst_pe_1_4_5_n9) );
  BUF_X1 npu_inst_pe_1_4_5_U5 ( .A(npu_inst_pe_1_4_5_n11), .Z(
        npu_inst_pe_1_4_5_n8) );
  NOR2_X1 npu_inst_pe_1_4_5_U4 ( .A1(npu_inst_pe_1_4_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_5_n1), .ZN(npu_inst_pe_1_4_5_n76) );
  NOR2_X1 npu_inst_pe_1_4_5_U3 ( .A1(npu_inst_pe_1_4_5_n27), .A2(
        npu_inst_pe_1_4_5_n1), .ZN(npu_inst_pe_1_4_5_n77) );
  FA_X1 npu_inst_pe_1_4_5_sub_77_U2_1 ( .A(npu_inst_int_data_res_4__5__1_), 
        .B(npu_inst_pe_1_4_5_n13), .CI(npu_inst_pe_1_4_5_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_4_5_sub_77_carry_2_), .S(npu_inst_pe_1_4_5_N66) );
  FA_X1 npu_inst_pe_1_4_5_add_79_U1_1 ( .A(npu_inst_int_data_res_4__5__1_), 
        .B(npu_inst_pe_1_4_5_int_data_1_), .CI(
        npu_inst_pe_1_4_5_add_79_carry_1_), .CO(
        npu_inst_pe_1_4_5_add_79_carry_2_), .S(npu_inst_pe_1_4_5_N74) );
  NAND3_X1 npu_inst_pe_1_4_5_U101 ( .A1(npu_inst_pe_1_4_5_n4), .A2(
        npu_inst_pe_1_4_5_n6), .A3(npu_inst_pe_1_4_5_n7), .ZN(
        npu_inst_pe_1_4_5_n44) );
  NAND3_X1 npu_inst_pe_1_4_5_U100 ( .A1(npu_inst_pe_1_4_5_n3), .A2(
        npu_inst_pe_1_4_5_n6), .A3(npu_inst_pe_1_4_5_n7), .ZN(
        npu_inst_pe_1_4_5_n40) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_5_n33), .CK(
        npu_inst_pe_1_4_5_net3627), .RN(npu_inst_pe_1_4_5_n8), .Q(
        npu_inst_int_data_res_4__5__6_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_5_n34), .CK(
        npu_inst_pe_1_4_5_net3627), .RN(npu_inst_pe_1_4_5_n8), .Q(
        npu_inst_int_data_res_4__5__5_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_5_n35), .CK(
        npu_inst_pe_1_4_5_net3627), .RN(npu_inst_pe_1_4_5_n8), .Q(
        npu_inst_int_data_res_4__5__4_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_5_n36), .CK(
        npu_inst_pe_1_4_5_net3627), .RN(npu_inst_pe_1_4_5_n8), .Q(
        npu_inst_int_data_res_4__5__3_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_5_n98), .CK(
        npu_inst_pe_1_4_5_net3627), .RN(npu_inst_pe_1_4_5_n8), .Q(
        npu_inst_int_data_res_4__5__2_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_5_n99), .CK(
        npu_inst_pe_1_4_5_net3627), .RN(npu_inst_pe_1_4_5_n8), .Q(
        npu_inst_int_data_res_4__5__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_5_n32), .CK(
        npu_inst_pe_1_4_5_net3627), .RN(npu_inst_pe_1_4_5_n8), .Q(
        npu_inst_int_data_res_4__5__7_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_5_n100), 
        .CK(npu_inst_pe_1_4_5_net3627), .RN(npu_inst_pe_1_4_5_n8), .Q(
        npu_inst_int_data_res_4__5__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_weight_reg_0_ ( .D(npu_inst_n92), .CK(
        npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n8), .Q(
        npu_inst_pe_1_4_5_int_q_weight_0_), .QN(npu_inst_pe_1_4_5_n27) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_weight_reg_1_ ( .D(npu_inst_n98), .CK(
        npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n8), .Q(
        npu_inst_pe_1_4_5_int_q_weight_1_), .QN(npu_inst_pe_1_4_5_n26) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_5_n112), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n8), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_5_n106), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n8), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_5_n111), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_5_n105), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_5_n110), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_5_n104), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_5_n109), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_5_n103), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_5_n108), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_5_n102), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_5_n107), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_5_n101), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_5_n86), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_5_n87), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n9), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_5_n88), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_5_n89), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_5_n90), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_5_n91), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_5_n92), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_5_n93), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_5_n94), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_5_n95), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_5_n96), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_5_n97), 
        .CK(npu_inst_pe_1_4_5_net3633), .RN(npu_inst_pe_1_4_5_n10), .Q(
        npu_inst_pe_1_4_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_5_net3627) );
  CLKGATETST_X1 npu_inst_pe_1_4_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n45), .SE(1'b0), .GCK(npu_inst_pe_1_4_5_net3633) );
  MUX2_X1 npu_inst_pe_1_4_6_U153 ( .A(npu_inst_pe_1_4_6_n31), .B(
        npu_inst_pe_1_4_6_n28), .S(npu_inst_pe_1_4_6_n7), .Z(
        npu_inst_pe_1_4_6_N93) );
  MUX2_X1 npu_inst_pe_1_4_6_U152 ( .A(npu_inst_pe_1_4_6_n30), .B(
        npu_inst_pe_1_4_6_n29), .S(npu_inst_pe_1_4_6_n5), .Z(
        npu_inst_pe_1_4_6_n31) );
  MUX2_X1 npu_inst_pe_1_4_6_U151 ( .A(npu_inst_pe_1_4_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_6_n3), .Z(
        npu_inst_pe_1_4_6_n30) );
  MUX2_X1 npu_inst_pe_1_4_6_U150 ( .A(npu_inst_pe_1_4_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_6_n3), .Z(
        npu_inst_pe_1_4_6_n29) );
  MUX2_X1 npu_inst_pe_1_4_6_U149 ( .A(npu_inst_pe_1_4_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_6_n3), .Z(
        npu_inst_pe_1_4_6_n28) );
  MUX2_X1 npu_inst_pe_1_4_6_U148 ( .A(npu_inst_pe_1_4_6_n25), .B(
        npu_inst_pe_1_4_6_n22), .S(npu_inst_pe_1_4_6_n7), .Z(
        npu_inst_pe_1_4_6_N94) );
  MUX2_X1 npu_inst_pe_1_4_6_U147 ( .A(npu_inst_pe_1_4_6_n24), .B(
        npu_inst_pe_1_4_6_n23), .S(npu_inst_pe_1_4_6_n5), .Z(
        npu_inst_pe_1_4_6_n25) );
  MUX2_X1 npu_inst_pe_1_4_6_U146 ( .A(npu_inst_pe_1_4_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_6_n3), .Z(
        npu_inst_pe_1_4_6_n24) );
  MUX2_X1 npu_inst_pe_1_4_6_U145 ( .A(npu_inst_pe_1_4_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_6_n3), .Z(
        npu_inst_pe_1_4_6_n23) );
  MUX2_X1 npu_inst_pe_1_4_6_U144 ( .A(npu_inst_pe_1_4_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_6_n3), .Z(
        npu_inst_pe_1_4_6_n22) );
  MUX2_X1 npu_inst_pe_1_4_6_U143 ( .A(npu_inst_pe_1_4_6_n21), .B(
        npu_inst_pe_1_4_6_n18), .S(npu_inst_pe_1_4_6_n7), .Z(
        npu_inst_int_data_x_4__6__1_) );
  MUX2_X1 npu_inst_pe_1_4_6_U142 ( .A(npu_inst_pe_1_4_6_n20), .B(
        npu_inst_pe_1_4_6_n19), .S(npu_inst_pe_1_4_6_n5), .Z(
        npu_inst_pe_1_4_6_n21) );
  MUX2_X1 npu_inst_pe_1_4_6_U141 ( .A(npu_inst_pe_1_4_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_6_n3), .Z(
        npu_inst_pe_1_4_6_n20) );
  MUX2_X1 npu_inst_pe_1_4_6_U140 ( .A(npu_inst_pe_1_4_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_6_n3), .Z(
        npu_inst_pe_1_4_6_n19) );
  MUX2_X1 npu_inst_pe_1_4_6_U139 ( .A(npu_inst_pe_1_4_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_6_n3), .Z(
        npu_inst_pe_1_4_6_n18) );
  MUX2_X1 npu_inst_pe_1_4_6_U138 ( .A(npu_inst_pe_1_4_6_n17), .B(
        npu_inst_pe_1_4_6_n14), .S(npu_inst_pe_1_4_6_n7), .Z(
        npu_inst_int_data_x_4__6__0_) );
  MUX2_X1 npu_inst_pe_1_4_6_U137 ( .A(npu_inst_pe_1_4_6_n16), .B(
        npu_inst_pe_1_4_6_n15), .S(npu_inst_pe_1_4_6_n5), .Z(
        npu_inst_pe_1_4_6_n17) );
  MUX2_X1 npu_inst_pe_1_4_6_U136 ( .A(npu_inst_pe_1_4_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_6_n3), .Z(
        npu_inst_pe_1_4_6_n16) );
  MUX2_X1 npu_inst_pe_1_4_6_U135 ( .A(npu_inst_pe_1_4_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_6_n3), .Z(
        npu_inst_pe_1_4_6_n15) );
  MUX2_X1 npu_inst_pe_1_4_6_U134 ( .A(npu_inst_pe_1_4_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_6_n3), .Z(
        npu_inst_pe_1_4_6_n14) );
  XOR2_X1 npu_inst_pe_1_4_6_U133 ( .A(npu_inst_pe_1_4_6_int_data_0_), .B(
        npu_inst_int_data_res_4__6__0_), .Z(npu_inst_pe_1_4_6_N73) );
  AND2_X1 npu_inst_pe_1_4_6_U132 ( .A1(npu_inst_int_data_res_4__6__0_), .A2(
        npu_inst_pe_1_4_6_int_data_0_), .ZN(npu_inst_pe_1_4_6_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_6_U131 ( .A(npu_inst_int_data_res_4__6__0_), .B(
        npu_inst_pe_1_4_6_n12), .ZN(npu_inst_pe_1_4_6_N65) );
  OR2_X1 npu_inst_pe_1_4_6_U130 ( .A1(npu_inst_pe_1_4_6_n12), .A2(
        npu_inst_int_data_res_4__6__0_), .ZN(npu_inst_pe_1_4_6_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_6_U129 ( .A(npu_inst_int_data_res_4__6__2_), .B(
        npu_inst_pe_1_4_6_add_79_carry_2_), .Z(npu_inst_pe_1_4_6_N75) );
  AND2_X1 npu_inst_pe_1_4_6_U128 ( .A1(npu_inst_pe_1_4_6_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_4__6__2_), .ZN(
        npu_inst_pe_1_4_6_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_6_U127 ( .A(npu_inst_int_data_res_4__6__3_), .B(
        npu_inst_pe_1_4_6_add_79_carry_3_), .Z(npu_inst_pe_1_4_6_N76) );
  AND2_X1 npu_inst_pe_1_4_6_U126 ( .A1(npu_inst_pe_1_4_6_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_4__6__3_), .ZN(
        npu_inst_pe_1_4_6_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_6_U125 ( .A(npu_inst_int_data_res_4__6__4_), .B(
        npu_inst_pe_1_4_6_add_79_carry_4_), .Z(npu_inst_pe_1_4_6_N77) );
  AND2_X1 npu_inst_pe_1_4_6_U124 ( .A1(npu_inst_pe_1_4_6_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_4__6__4_), .ZN(
        npu_inst_pe_1_4_6_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_6_U123 ( .A(npu_inst_int_data_res_4__6__5_), .B(
        npu_inst_pe_1_4_6_add_79_carry_5_), .Z(npu_inst_pe_1_4_6_N78) );
  AND2_X1 npu_inst_pe_1_4_6_U122 ( .A1(npu_inst_pe_1_4_6_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_4__6__5_), .ZN(
        npu_inst_pe_1_4_6_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_6_U121 ( .A(npu_inst_int_data_res_4__6__6_), .B(
        npu_inst_pe_1_4_6_add_79_carry_6_), .Z(npu_inst_pe_1_4_6_N79) );
  AND2_X1 npu_inst_pe_1_4_6_U120 ( .A1(npu_inst_pe_1_4_6_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_4__6__6_), .ZN(
        npu_inst_pe_1_4_6_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_6_U119 ( .A(npu_inst_int_data_res_4__6__7_), .B(
        npu_inst_pe_1_4_6_add_79_carry_7_), .Z(npu_inst_pe_1_4_6_N80) );
  XNOR2_X1 npu_inst_pe_1_4_6_U118 ( .A(npu_inst_pe_1_4_6_sub_77_carry_2_), .B(
        npu_inst_int_data_res_4__6__2_), .ZN(npu_inst_pe_1_4_6_N67) );
  OR2_X1 npu_inst_pe_1_4_6_U117 ( .A1(npu_inst_int_data_res_4__6__2_), .A2(
        npu_inst_pe_1_4_6_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_4_6_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_6_U116 ( .A(npu_inst_pe_1_4_6_sub_77_carry_3_), .B(
        npu_inst_int_data_res_4__6__3_), .ZN(npu_inst_pe_1_4_6_N68) );
  OR2_X1 npu_inst_pe_1_4_6_U115 ( .A1(npu_inst_int_data_res_4__6__3_), .A2(
        npu_inst_pe_1_4_6_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_4_6_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_6_U114 ( .A(npu_inst_pe_1_4_6_sub_77_carry_4_), .B(
        npu_inst_int_data_res_4__6__4_), .ZN(npu_inst_pe_1_4_6_N69) );
  OR2_X1 npu_inst_pe_1_4_6_U113 ( .A1(npu_inst_int_data_res_4__6__4_), .A2(
        npu_inst_pe_1_4_6_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_4_6_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_6_U112 ( .A(npu_inst_pe_1_4_6_sub_77_carry_5_), .B(
        npu_inst_int_data_res_4__6__5_), .ZN(npu_inst_pe_1_4_6_N70) );
  OR2_X1 npu_inst_pe_1_4_6_U111 ( .A1(npu_inst_int_data_res_4__6__5_), .A2(
        npu_inst_pe_1_4_6_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_4_6_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_6_U110 ( .A(npu_inst_pe_1_4_6_sub_77_carry_6_), .B(
        npu_inst_int_data_res_4__6__6_), .ZN(npu_inst_pe_1_4_6_N71) );
  OR2_X1 npu_inst_pe_1_4_6_U109 ( .A1(npu_inst_int_data_res_4__6__6_), .A2(
        npu_inst_pe_1_4_6_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_4_6_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_6_U108 ( .A(npu_inst_int_data_res_4__6__7_), .B(
        npu_inst_pe_1_4_6_sub_77_carry_7_), .ZN(npu_inst_pe_1_4_6_N72) );
  INV_X1 npu_inst_pe_1_4_6_U107 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_4_6_n6)
         );
  INV_X1 npu_inst_pe_1_4_6_U106 ( .A(npu_inst_pe_1_4_6_n6), .ZN(
        npu_inst_pe_1_4_6_n5) );
  INV_X1 npu_inst_pe_1_4_6_U105 ( .A(npu_inst_n37), .ZN(npu_inst_pe_1_4_6_n2)
         );
  AOI22_X1 npu_inst_pe_1_4_6_U104 ( .A1(npu_inst_int_data_y_5__6__0_), .A2(
        npu_inst_pe_1_4_6_n58), .B1(npu_inst_pe_1_4_6_n118), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_6_n57) );
  INV_X1 npu_inst_pe_1_4_6_U103 ( .A(npu_inst_pe_1_4_6_n57), .ZN(
        npu_inst_pe_1_4_6_n107) );
  AOI22_X1 npu_inst_pe_1_4_6_U102 ( .A1(npu_inst_int_data_y_5__6__0_), .A2(
        npu_inst_pe_1_4_6_n54), .B1(npu_inst_pe_1_4_6_n117), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_6_n53) );
  INV_X1 npu_inst_pe_1_4_6_U99 ( .A(npu_inst_pe_1_4_6_n53), .ZN(
        npu_inst_pe_1_4_6_n108) );
  AOI22_X1 npu_inst_pe_1_4_6_U98 ( .A1(npu_inst_int_data_y_5__6__0_), .A2(
        npu_inst_pe_1_4_6_n50), .B1(npu_inst_pe_1_4_6_n116), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_6_n49) );
  INV_X1 npu_inst_pe_1_4_6_U97 ( .A(npu_inst_pe_1_4_6_n49), .ZN(
        npu_inst_pe_1_4_6_n109) );
  AOI22_X1 npu_inst_pe_1_4_6_U96 ( .A1(npu_inst_int_data_y_5__6__0_), .A2(
        npu_inst_pe_1_4_6_n46), .B1(npu_inst_pe_1_4_6_n115), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_6_n45) );
  INV_X1 npu_inst_pe_1_4_6_U95 ( .A(npu_inst_pe_1_4_6_n45), .ZN(
        npu_inst_pe_1_4_6_n110) );
  AOI22_X1 npu_inst_pe_1_4_6_U94 ( .A1(npu_inst_int_data_y_5__6__0_), .A2(
        npu_inst_pe_1_4_6_n42), .B1(npu_inst_pe_1_4_6_n114), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_6_n41) );
  INV_X1 npu_inst_pe_1_4_6_U93 ( .A(npu_inst_pe_1_4_6_n41), .ZN(
        npu_inst_pe_1_4_6_n111) );
  AOI22_X1 npu_inst_pe_1_4_6_U92 ( .A1(npu_inst_int_data_y_5__6__1_), .A2(
        npu_inst_pe_1_4_6_n58), .B1(npu_inst_pe_1_4_6_n118), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_6_n59) );
  INV_X1 npu_inst_pe_1_4_6_U91 ( .A(npu_inst_pe_1_4_6_n59), .ZN(
        npu_inst_pe_1_4_6_n101) );
  AOI22_X1 npu_inst_pe_1_4_6_U90 ( .A1(npu_inst_int_data_y_5__6__1_), .A2(
        npu_inst_pe_1_4_6_n54), .B1(npu_inst_pe_1_4_6_n117), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_6_n55) );
  INV_X1 npu_inst_pe_1_4_6_U89 ( .A(npu_inst_pe_1_4_6_n55), .ZN(
        npu_inst_pe_1_4_6_n102) );
  AOI22_X1 npu_inst_pe_1_4_6_U88 ( .A1(npu_inst_int_data_y_5__6__1_), .A2(
        npu_inst_pe_1_4_6_n50), .B1(npu_inst_pe_1_4_6_n116), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_6_n51) );
  INV_X1 npu_inst_pe_1_4_6_U87 ( .A(npu_inst_pe_1_4_6_n51), .ZN(
        npu_inst_pe_1_4_6_n103) );
  AOI22_X1 npu_inst_pe_1_4_6_U86 ( .A1(npu_inst_int_data_y_5__6__1_), .A2(
        npu_inst_pe_1_4_6_n46), .B1(npu_inst_pe_1_4_6_n115), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_6_n47) );
  INV_X1 npu_inst_pe_1_4_6_U85 ( .A(npu_inst_pe_1_4_6_n47), .ZN(
        npu_inst_pe_1_4_6_n104) );
  AOI22_X1 npu_inst_pe_1_4_6_U84 ( .A1(npu_inst_int_data_y_5__6__1_), .A2(
        npu_inst_pe_1_4_6_n42), .B1(npu_inst_pe_1_4_6_n114), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_6_n43) );
  INV_X1 npu_inst_pe_1_4_6_U83 ( .A(npu_inst_pe_1_4_6_n43), .ZN(
        npu_inst_pe_1_4_6_n105) );
  AOI22_X1 npu_inst_pe_1_4_6_U82 ( .A1(npu_inst_pe_1_4_6_n38), .A2(
        npu_inst_int_data_y_5__6__1_), .B1(npu_inst_pe_1_4_6_n113), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_6_n39) );
  INV_X1 npu_inst_pe_1_4_6_U81 ( .A(npu_inst_pe_1_4_6_n39), .ZN(
        npu_inst_pe_1_4_6_n106) );
  AND2_X1 npu_inst_pe_1_4_6_U80 ( .A1(npu_inst_pe_1_4_6_N93), .A2(npu_inst_n37), .ZN(npu_inst_int_data_y_4__6__0_) );
  NAND2_X1 npu_inst_pe_1_4_6_U79 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_6_n60), .ZN(npu_inst_pe_1_4_6_n74) );
  OAI21_X1 npu_inst_pe_1_4_6_U78 ( .B1(npu_inst_pe_1_4_6_n63), .B2(
        npu_inst_pe_1_4_6_n60), .A(npu_inst_pe_1_4_6_n74), .ZN(
        npu_inst_pe_1_4_6_n97) );
  NAND2_X1 npu_inst_pe_1_4_6_U77 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_6_n60), .ZN(npu_inst_pe_1_4_6_n73) );
  OAI21_X1 npu_inst_pe_1_4_6_U76 ( .B1(npu_inst_pe_1_4_6_n61), .B2(
        npu_inst_pe_1_4_6_n60), .A(npu_inst_pe_1_4_6_n73), .ZN(
        npu_inst_pe_1_4_6_n96) );
  NAND2_X1 npu_inst_pe_1_4_6_U75 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_6_n56), .ZN(npu_inst_pe_1_4_6_n72) );
  OAI21_X1 npu_inst_pe_1_4_6_U74 ( .B1(npu_inst_pe_1_4_6_n63), .B2(
        npu_inst_pe_1_4_6_n56), .A(npu_inst_pe_1_4_6_n72), .ZN(
        npu_inst_pe_1_4_6_n95) );
  NAND2_X1 npu_inst_pe_1_4_6_U73 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_6_n56), .ZN(npu_inst_pe_1_4_6_n71) );
  OAI21_X1 npu_inst_pe_1_4_6_U72 ( .B1(npu_inst_pe_1_4_6_n61), .B2(
        npu_inst_pe_1_4_6_n56), .A(npu_inst_pe_1_4_6_n71), .ZN(
        npu_inst_pe_1_4_6_n94) );
  NAND2_X1 npu_inst_pe_1_4_6_U71 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_6_n52), .ZN(npu_inst_pe_1_4_6_n70) );
  OAI21_X1 npu_inst_pe_1_4_6_U70 ( .B1(npu_inst_pe_1_4_6_n63), .B2(
        npu_inst_pe_1_4_6_n52), .A(npu_inst_pe_1_4_6_n70), .ZN(
        npu_inst_pe_1_4_6_n93) );
  NAND2_X1 npu_inst_pe_1_4_6_U69 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_6_n52), .ZN(npu_inst_pe_1_4_6_n69) );
  OAI21_X1 npu_inst_pe_1_4_6_U68 ( .B1(npu_inst_pe_1_4_6_n61), .B2(
        npu_inst_pe_1_4_6_n52), .A(npu_inst_pe_1_4_6_n69), .ZN(
        npu_inst_pe_1_4_6_n92) );
  NAND2_X1 npu_inst_pe_1_4_6_U67 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_6_n48), .ZN(npu_inst_pe_1_4_6_n68) );
  OAI21_X1 npu_inst_pe_1_4_6_U66 ( .B1(npu_inst_pe_1_4_6_n63), .B2(
        npu_inst_pe_1_4_6_n48), .A(npu_inst_pe_1_4_6_n68), .ZN(
        npu_inst_pe_1_4_6_n91) );
  NAND2_X1 npu_inst_pe_1_4_6_U65 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_6_n48), .ZN(npu_inst_pe_1_4_6_n67) );
  OAI21_X1 npu_inst_pe_1_4_6_U64 ( .B1(npu_inst_pe_1_4_6_n61), .B2(
        npu_inst_pe_1_4_6_n48), .A(npu_inst_pe_1_4_6_n67), .ZN(
        npu_inst_pe_1_4_6_n90) );
  NAND2_X1 npu_inst_pe_1_4_6_U63 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_6_n44), .ZN(npu_inst_pe_1_4_6_n66) );
  OAI21_X1 npu_inst_pe_1_4_6_U62 ( .B1(npu_inst_pe_1_4_6_n63), .B2(
        npu_inst_pe_1_4_6_n44), .A(npu_inst_pe_1_4_6_n66), .ZN(
        npu_inst_pe_1_4_6_n89) );
  NAND2_X1 npu_inst_pe_1_4_6_U61 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_6_n44), .ZN(npu_inst_pe_1_4_6_n65) );
  OAI21_X1 npu_inst_pe_1_4_6_U60 ( .B1(npu_inst_pe_1_4_6_n61), .B2(
        npu_inst_pe_1_4_6_n44), .A(npu_inst_pe_1_4_6_n65), .ZN(
        npu_inst_pe_1_4_6_n88) );
  NAND2_X1 npu_inst_pe_1_4_6_U59 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_6_n40), .ZN(npu_inst_pe_1_4_6_n64) );
  OAI21_X1 npu_inst_pe_1_4_6_U58 ( .B1(npu_inst_pe_1_4_6_n63), .B2(
        npu_inst_pe_1_4_6_n40), .A(npu_inst_pe_1_4_6_n64), .ZN(
        npu_inst_pe_1_4_6_n87) );
  NAND2_X1 npu_inst_pe_1_4_6_U57 ( .A1(npu_inst_pe_1_4_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_6_n40), .ZN(npu_inst_pe_1_4_6_n62) );
  OAI21_X1 npu_inst_pe_1_4_6_U56 ( .B1(npu_inst_pe_1_4_6_n61), .B2(
        npu_inst_pe_1_4_6_n40), .A(npu_inst_pe_1_4_6_n62), .ZN(
        npu_inst_pe_1_4_6_n86) );
  AOI22_X1 npu_inst_pe_1_4_6_U55 ( .A1(npu_inst_pe_1_4_6_n38), .A2(
        npu_inst_int_data_y_5__6__0_), .B1(npu_inst_pe_1_4_6_n113), .B2(
        npu_inst_pe_1_4_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_6_n37) );
  INV_X1 npu_inst_pe_1_4_6_U54 ( .A(npu_inst_pe_1_4_6_n37), .ZN(
        npu_inst_pe_1_4_6_n112) );
  AND2_X1 npu_inst_pe_1_4_6_U53 ( .A1(npu_inst_n37), .A2(npu_inst_pe_1_4_6_N94), .ZN(npu_inst_int_data_y_4__6__1_) );
  AOI222_X1 npu_inst_pe_1_4_6_U52 ( .A1(npu_inst_int_data_res_5__6__0_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N73), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N65), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n84) );
  INV_X1 npu_inst_pe_1_4_6_U51 ( .A(npu_inst_pe_1_4_6_n84), .ZN(
        npu_inst_pe_1_4_6_n100) );
  AOI222_X1 npu_inst_pe_1_4_6_U50 ( .A1(npu_inst_pe_1_4_6_n1), .A2(
        npu_inst_int_data_res_5__6__7_), .B1(npu_inst_pe_1_4_6_N80), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N72), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n75) );
  INV_X1 npu_inst_pe_1_4_6_U49 ( .A(npu_inst_pe_1_4_6_n75), .ZN(
        npu_inst_pe_1_4_6_n32) );
  AOI222_X1 npu_inst_pe_1_4_6_U48 ( .A1(npu_inst_int_data_res_5__6__1_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N74), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N66), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n83) );
  INV_X1 npu_inst_pe_1_4_6_U47 ( .A(npu_inst_pe_1_4_6_n83), .ZN(
        npu_inst_pe_1_4_6_n99) );
  AOI222_X1 npu_inst_pe_1_4_6_U46 ( .A1(npu_inst_int_data_res_5__6__3_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N76), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N68), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n81) );
  INV_X1 npu_inst_pe_1_4_6_U45 ( .A(npu_inst_pe_1_4_6_n81), .ZN(
        npu_inst_pe_1_4_6_n36) );
  AOI222_X1 npu_inst_pe_1_4_6_U44 ( .A1(npu_inst_int_data_res_5__6__4_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N77), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N69), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n80) );
  INV_X1 npu_inst_pe_1_4_6_U43 ( .A(npu_inst_pe_1_4_6_n80), .ZN(
        npu_inst_pe_1_4_6_n35) );
  AOI222_X1 npu_inst_pe_1_4_6_U42 ( .A1(npu_inst_int_data_res_5__6__5_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N78), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N70), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n79) );
  INV_X1 npu_inst_pe_1_4_6_U41 ( .A(npu_inst_pe_1_4_6_n79), .ZN(
        npu_inst_pe_1_4_6_n34) );
  AOI222_X1 npu_inst_pe_1_4_6_U40 ( .A1(npu_inst_int_data_res_5__6__6_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N79), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N71), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n78) );
  INV_X1 npu_inst_pe_1_4_6_U39 ( .A(npu_inst_pe_1_4_6_n78), .ZN(
        npu_inst_pe_1_4_6_n33) );
  AND2_X1 npu_inst_pe_1_4_6_U38 ( .A1(npu_inst_int_data_x_4__6__1_), .A2(
        npu_inst_pe_1_4_6_int_q_weight_1_), .ZN(npu_inst_pe_1_4_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_6_U37 ( .A1(npu_inst_int_data_x_4__6__0_), .A2(
        npu_inst_pe_1_4_6_int_q_weight_1_), .ZN(npu_inst_pe_1_4_6_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_4_6_U36 ( .A(npu_inst_pe_1_4_6_int_data_1_), .ZN(
        npu_inst_pe_1_4_6_n13) );
  NOR3_X1 npu_inst_pe_1_4_6_U35 ( .A1(npu_inst_pe_1_4_6_n26), .A2(npu_inst_n37), .A3(npu_inst_int_ckg[25]), .ZN(npu_inst_pe_1_4_6_n85) );
  OR2_X1 npu_inst_pe_1_4_6_U34 ( .A1(npu_inst_pe_1_4_6_n85), .A2(
        npu_inst_pe_1_4_6_n1), .ZN(npu_inst_pe_1_4_6_N84) );
  AOI222_X1 npu_inst_pe_1_4_6_U33 ( .A1(npu_inst_int_data_res_5__6__2_), .A2(
        npu_inst_pe_1_4_6_n1), .B1(npu_inst_pe_1_4_6_N75), .B2(
        npu_inst_pe_1_4_6_n76), .C1(npu_inst_pe_1_4_6_N67), .C2(
        npu_inst_pe_1_4_6_n77), .ZN(npu_inst_pe_1_4_6_n82) );
  INV_X1 npu_inst_pe_1_4_6_U32 ( .A(npu_inst_pe_1_4_6_n82), .ZN(
        npu_inst_pe_1_4_6_n98) );
  AOI22_X1 npu_inst_pe_1_4_6_U31 ( .A1(npu_inst_n37), .A2(
        npu_inst_int_data_y_5__6__1_), .B1(npu_inst_pe_1_4_6_n2), .B2(
        npu_inst_int_data_x_4__7__1_), .ZN(npu_inst_pe_1_4_6_n63) );
  AOI22_X1 npu_inst_pe_1_4_6_U30 ( .A1(npu_inst_n37), .A2(
        npu_inst_int_data_y_5__6__0_), .B1(npu_inst_pe_1_4_6_n2), .B2(
        npu_inst_int_data_x_4__7__0_), .ZN(npu_inst_pe_1_4_6_n61) );
  INV_X1 npu_inst_pe_1_4_6_U29 ( .A(npu_inst_pe_1_4_6_int_data_0_), .ZN(
        npu_inst_pe_1_4_6_n12) );
  INV_X1 npu_inst_pe_1_4_6_U28 ( .A(npu_inst_n51), .ZN(npu_inst_pe_1_4_6_n4)
         );
  OR3_X1 npu_inst_pe_1_4_6_U27 ( .A1(npu_inst_pe_1_4_6_n5), .A2(
        npu_inst_pe_1_4_6_n7), .A3(npu_inst_pe_1_4_6_n4), .ZN(
        npu_inst_pe_1_4_6_n56) );
  OR3_X1 npu_inst_pe_1_4_6_U26 ( .A1(npu_inst_pe_1_4_6_n4), .A2(
        npu_inst_pe_1_4_6_n7), .A3(npu_inst_pe_1_4_6_n6), .ZN(
        npu_inst_pe_1_4_6_n48) );
  INV_X1 npu_inst_pe_1_4_6_U25 ( .A(npu_inst_pe_1_4_6_n4), .ZN(
        npu_inst_pe_1_4_6_n3) );
  OR3_X1 npu_inst_pe_1_4_6_U24 ( .A1(npu_inst_pe_1_4_6_n3), .A2(
        npu_inst_pe_1_4_6_n7), .A3(npu_inst_pe_1_4_6_n6), .ZN(
        npu_inst_pe_1_4_6_n52) );
  OR3_X1 npu_inst_pe_1_4_6_U23 ( .A1(npu_inst_pe_1_4_6_n5), .A2(
        npu_inst_pe_1_4_6_n7), .A3(npu_inst_pe_1_4_6_n3), .ZN(
        npu_inst_pe_1_4_6_n60) );
  BUF_X1 npu_inst_pe_1_4_6_U22 ( .A(npu_inst_n19), .Z(npu_inst_pe_1_4_6_n1) );
  NOR2_X1 npu_inst_pe_1_4_6_U21 ( .A1(npu_inst_pe_1_4_6_n60), .A2(
        npu_inst_pe_1_4_6_n2), .ZN(npu_inst_pe_1_4_6_n58) );
  NOR2_X1 npu_inst_pe_1_4_6_U20 ( .A1(npu_inst_pe_1_4_6_n56), .A2(
        npu_inst_pe_1_4_6_n2), .ZN(npu_inst_pe_1_4_6_n54) );
  NOR2_X1 npu_inst_pe_1_4_6_U19 ( .A1(npu_inst_pe_1_4_6_n52), .A2(
        npu_inst_pe_1_4_6_n2), .ZN(npu_inst_pe_1_4_6_n50) );
  NOR2_X1 npu_inst_pe_1_4_6_U18 ( .A1(npu_inst_pe_1_4_6_n48), .A2(
        npu_inst_pe_1_4_6_n2), .ZN(npu_inst_pe_1_4_6_n46) );
  NOR2_X1 npu_inst_pe_1_4_6_U17 ( .A1(npu_inst_pe_1_4_6_n40), .A2(
        npu_inst_pe_1_4_6_n2), .ZN(npu_inst_pe_1_4_6_n38) );
  NOR2_X1 npu_inst_pe_1_4_6_U16 ( .A1(npu_inst_pe_1_4_6_n44), .A2(
        npu_inst_pe_1_4_6_n2), .ZN(npu_inst_pe_1_4_6_n42) );
  BUF_X1 npu_inst_pe_1_4_6_U15 ( .A(npu_inst_n80), .Z(npu_inst_pe_1_4_6_n7) );
  INV_X1 npu_inst_pe_1_4_6_U14 ( .A(npu_inst_n106), .ZN(npu_inst_pe_1_4_6_n11)
         );
  INV_X1 npu_inst_pe_1_4_6_U13 ( .A(npu_inst_pe_1_4_6_n38), .ZN(
        npu_inst_pe_1_4_6_n113) );
  INV_X1 npu_inst_pe_1_4_6_U12 ( .A(npu_inst_pe_1_4_6_n58), .ZN(
        npu_inst_pe_1_4_6_n118) );
  INV_X1 npu_inst_pe_1_4_6_U11 ( .A(npu_inst_pe_1_4_6_n54), .ZN(
        npu_inst_pe_1_4_6_n117) );
  INV_X1 npu_inst_pe_1_4_6_U10 ( .A(npu_inst_pe_1_4_6_n50), .ZN(
        npu_inst_pe_1_4_6_n116) );
  INV_X1 npu_inst_pe_1_4_6_U9 ( .A(npu_inst_pe_1_4_6_n46), .ZN(
        npu_inst_pe_1_4_6_n115) );
  INV_X1 npu_inst_pe_1_4_6_U8 ( .A(npu_inst_pe_1_4_6_n42), .ZN(
        npu_inst_pe_1_4_6_n114) );
  BUF_X1 npu_inst_pe_1_4_6_U7 ( .A(npu_inst_pe_1_4_6_n11), .Z(
        npu_inst_pe_1_4_6_n10) );
  BUF_X1 npu_inst_pe_1_4_6_U6 ( .A(npu_inst_pe_1_4_6_n11), .Z(
        npu_inst_pe_1_4_6_n9) );
  BUF_X1 npu_inst_pe_1_4_6_U5 ( .A(npu_inst_pe_1_4_6_n11), .Z(
        npu_inst_pe_1_4_6_n8) );
  NOR2_X1 npu_inst_pe_1_4_6_U4 ( .A1(npu_inst_pe_1_4_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_6_n1), .ZN(npu_inst_pe_1_4_6_n76) );
  NOR2_X1 npu_inst_pe_1_4_6_U3 ( .A1(npu_inst_pe_1_4_6_n27), .A2(
        npu_inst_pe_1_4_6_n1), .ZN(npu_inst_pe_1_4_6_n77) );
  FA_X1 npu_inst_pe_1_4_6_sub_77_U2_1 ( .A(npu_inst_int_data_res_4__6__1_), 
        .B(npu_inst_pe_1_4_6_n13), .CI(npu_inst_pe_1_4_6_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_4_6_sub_77_carry_2_), .S(npu_inst_pe_1_4_6_N66) );
  FA_X1 npu_inst_pe_1_4_6_add_79_U1_1 ( .A(npu_inst_int_data_res_4__6__1_), 
        .B(npu_inst_pe_1_4_6_int_data_1_), .CI(
        npu_inst_pe_1_4_6_add_79_carry_1_), .CO(
        npu_inst_pe_1_4_6_add_79_carry_2_), .S(npu_inst_pe_1_4_6_N74) );
  NAND3_X1 npu_inst_pe_1_4_6_U101 ( .A1(npu_inst_pe_1_4_6_n4), .A2(
        npu_inst_pe_1_4_6_n6), .A3(npu_inst_pe_1_4_6_n7), .ZN(
        npu_inst_pe_1_4_6_n44) );
  NAND3_X1 npu_inst_pe_1_4_6_U100 ( .A1(npu_inst_pe_1_4_6_n3), .A2(
        npu_inst_pe_1_4_6_n6), .A3(npu_inst_pe_1_4_6_n7), .ZN(
        npu_inst_pe_1_4_6_n40) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_6_n33), .CK(
        npu_inst_pe_1_4_6_net3604), .RN(npu_inst_pe_1_4_6_n8), .Q(
        npu_inst_int_data_res_4__6__6_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_6_n34), .CK(
        npu_inst_pe_1_4_6_net3604), .RN(npu_inst_pe_1_4_6_n8), .Q(
        npu_inst_int_data_res_4__6__5_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_6_n35), .CK(
        npu_inst_pe_1_4_6_net3604), .RN(npu_inst_pe_1_4_6_n8), .Q(
        npu_inst_int_data_res_4__6__4_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_6_n36), .CK(
        npu_inst_pe_1_4_6_net3604), .RN(npu_inst_pe_1_4_6_n8), .Q(
        npu_inst_int_data_res_4__6__3_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_6_n98), .CK(
        npu_inst_pe_1_4_6_net3604), .RN(npu_inst_pe_1_4_6_n8), .Q(
        npu_inst_int_data_res_4__6__2_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_6_n99), .CK(
        npu_inst_pe_1_4_6_net3604), .RN(npu_inst_pe_1_4_6_n8), .Q(
        npu_inst_int_data_res_4__6__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_6_n32), .CK(
        npu_inst_pe_1_4_6_net3604), .RN(npu_inst_pe_1_4_6_n8), .Q(
        npu_inst_int_data_res_4__6__7_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_6_n100), 
        .CK(npu_inst_pe_1_4_6_net3604), .RN(npu_inst_pe_1_4_6_n8), .Q(
        npu_inst_int_data_res_4__6__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_weight_reg_0_ ( .D(npu_inst_n92), .CK(
        npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n8), .Q(
        npu_inst_pe_1_4_6_int_q_weight_0_), .QN(npu_inst_pe_1_4_6_n27) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_weight_reg_1_ ( .D(npu_inst_n98), .CK(
        npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n8), .Q(
        npu_inst_pe_1_4_6_int_q_weight_1_), .QN(npu_inst_pe_1_4_6_n26) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_6_n112), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n8), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_6_n106), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n8), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_6_n111), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_6_n105), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_6_n110), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_6_n104), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_6_n109), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_6_n103), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_6_n108), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_6_n102), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_6_n107), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_6_n101), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_6_n86), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_6_n87), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n9), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_6_n88), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_6_n89), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_6_n90), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_6_n91), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_6_n92), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_6_n93), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_6_n94), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_6_n95), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_6_n96), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_6_n97), 
        .CK(npu_inst_pe_1_4_6_net3610), .RN(npu_inst_pe_1_4_6_n10), .Q(
        npu_inst_pe_1_4_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_6_net3604) );
  CLKGATETST_X1 npu_inst_pe_1_4_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n45), .SE(1'b0), .GCK(npu_inst_pe_1_4_6_net3610) );
  MUX2_X1 npu_inst_pe_1_4_7_U153 ( .A(npu_inst_pe_1_4_7_n31), .B(
        npu_inst_pe_1_4_7_n28), .S(npu_inst_pe_1_4_7_n7), .Z(
        npu_inst_pe_1_4_7_N93) );
  MUX2_X1 npu_inst_pe_1_4_7_U152 ( .A(npu_inst_pe_1_4_7_n30), .B(
        npu_inst_pe_1_4_7_n29), .S(npu_inst_pe_1_4_7_n5), .Z(
        npu_inst_pe_1_4_7_n31) );
  MUX2_X1 npu_inst_pe_1_4_7_U151 ( .A(npu_inst_pe_1_4_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_4_7_n3), .Z(
        npu_inst_pe_1_4_7_n30) );
  MUX2_X1 npu_inst_pe_1_4_7_U150 ( .A(npu_inst_pe_1_4_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_4_7_n3), .Z(
        npu_inst_pe_1_4_7_n29) );
  MUX2_X1 npu_inst_pe_1_4_7_U149 ( .A(npu_inst_pe_1_4_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_4_7_n3), .Z(
        npu_inst_pe_1_4_7_n28) );
  MUX2_X1 npu_inst_pe_1_4_7_U148 ( .A(npu_inst_pe_1_4_7_n25), .B(
        npu_inst_pe_1_4_7_n22), .S(npu_inst_pe_1_4_7_n7), .Z(
        npu_inst_pe_1_4_7_N94) );
  MUX2_X1 npu_inst_pe_1_4_7_U147 ( .A(npu_inst_pe_1_4_7_n24), .B(
        npu_inst_pe_1_4_7_n23), .S(npu_inst_pe_1_4_7_n5), .Z(
        npu_inst_pe_1_4_7_n25) );
  MUX2_X1 npu_inst_pe_1_4_7_U146 ( .A(npu_inst_pe_1_4_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_4_7_n3), .Z(
        npu_inst_pe_1_4_7_n24) );
  MUX2_X1 npu_inst_pe_1_4_7_U145 ( .A(npu_inst_pe_1_4_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_4_7_n3), .Z(
        npu_inst_pe_1_4_7_n23) );
  MUX2_X1 npu_inst_pe_1_4_7_U144 ( .A(npu_inst_pe_1_4_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_4_7_n3), .Z(
        npu_inst_pe_1_4_7_n22) );
  MUX2_X1 npu_inst_pe_1_4_7_U143 ( .A(npu_inst_pe_1_4_7_n21), .B(
        npu_inst_pe_1_4_7_n18), .S(npu_inst_pe_1_4_7_n7), .Z(
        npu_inst_int_data_x_4__7__1_) );
  MUX2_X1 npu_inst_pe_1_4_7_U142 ( .A(npu_inst_pe_1_4_7_n20), .B(
        npu_inst_pe_1_4_7_n19), .S(npu_inst_pe_1_4_7_n5), .Z(
        npu_inst_pe_1_4_7_n21) );
  MUX2_X1 npu_inst_pe_1_4_7_U141 ( .A(npu_inst_pe_1_4_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_4_7_n3), .Z(
        npu_inst_pe_1_4_7_n20) );
  MUX2_X1 npu_inst_pe_1_4_7_U140 ( .A(npu_inst_pe_1_4_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_4_7_n3), .Z(
        npu_inst_pe_1_4_7_n19) );
  MUX2_X1 npu_inst_pe_1_4_7_U139 ( .A(npu_inst_pe_1_4_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_4_7_n3), .Z(
        npu_inst_pe_1_4_7_n18) );
  MUX2_X1 npu_inst_pe_1_4_7_U138 ( .A(npu_inst_pe_1_4_7_n17), .B(
        npu_inst_pe_1_4_7_n14), .S(npu_inst_pe_1_4_7_n7), .Z(
        npu_inst_int_data_x_4__7__0_) );
  MUX2_X1 npu_inst_pe_1_4_7_U137 ( .A(npu_inst_pe_1_4_7_n16), .B(
        npu_inst_pe_1_4_7_n15), .S(npu_inst_pe_1_4_7_n5), .Z(
        npu_inst_pe_1_4_7_n17) );
  MUX2_X1 npu_inst_pe_1_4_7_U136 ( .A(npu_inst_pe_1_4_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_4_7_n3), .Z(
        npu_inst_pe_1_4_7_n16) );
  MUX2_X1 npu_inst_pe_1_4_7_U135 ( .A(npu_inst_pe_1_4_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_4_7_n3), .Z(
        npu_inst_pe_1_4_7_n15) );
  MUX2_X1 npu_inst_pe_1_4_7_U134 ( .A(npu_inst_pe_1_4_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_4_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_4_7_n3), .Z(
        npu_inst_pe_1_4_7_n14) );
  XOR2_X1 npu_inst_pe_1_4_7_U133 ( .A(npu_inst_pe_1_4_7_int_data_0_), .B(
        npu_inst_int_data_res_4__7__0_), .Z(npu_inst_pe_1_4_7_N73) );
  AND2_X1 npu_inst_pe_1_4_7_U132 ( .A1(npu_inst_int_data_res_4__7__0_), .A2(
        npu_inst_pe_1_4_7_int_data_0_), .ZN(npu_inst_pe_1_4_7_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_4_7_U131 ( .A(npu_inst_int_data_res_4__7__0_), .B(
        npu_inst_pe_1_4_7_n12), .ZN(npu_inst_pe_1_4_7_N65) );
  OR2_X1 npu_inst_pe_1_4_7_U130 ( .A1(npu_inst_pe_1_4_7_n12), .A2(
        npu_inst_int_data_res_4__7__0_), .ZN(npu_inst_pe_1_4_7_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_4_7_U129 ( .A(npu_inst_int_data_res_4__7__2_), .B(
        npu_inst_pe_1_4_7_add_79_carry_2_), .Z(npu_inst_pe_1_4_7_N75) );
  AND2_X1 npu_inst_pe_1_4_7_U128 ( .A1(npu_inst_pe_1_4_7_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_4__7__2_), .ZN(
        npu_inst_pe_1_4_7_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_4_7_U127 ( .A(npu_inst_int_data_res_4__7__3_), .B(
        npu_inst_pe_1_4_7_add_79_carry_3_), .Z(npu_inst_pe_1_4_7_N76) );
  AND2_X1 npu_inst_pe_1_4_7_U126 ( .A1(npu_inst_pe_1_4_7_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_4__7__3_), .ZN(
        npu_inst_pe_1_4_7_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_4_7_U125 ( .A(npu_inst_int_data_res_4__7__4_), .B(
        npu_inst_pe_1_4_7_add_79_carry_4_), .Z(npu_inst_pe_1_4_7_N77) );
  AND2_X1 npu_inst_pe_1_4_7_U124 ( .A1(npu_inst_pe_1_4_7_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_4__7__4_), .ZN(
        npu_inst_pe_1_4_7_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_4_7_U123 ( .A(npu_inst_int_data_res_4__7__5_), .B(
        npu_inst_pe_1_4_7_add_79_carry_5_), .Z(npu_inst_pe_1_4_7_N78) );
  AND2_X1 npu_inst_pe_1_4_7_U122 ( .A1(npu_inst_pe_1_4_7_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_4__7__5_), .ZN(
        npu_inst_pe_1_4_7_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_4_7_U121 ( .A(npu_inst_int_data_res_4__7__6_), .B(
        npu_inst_pe_1_4_7_add_79_carry_6_), .Z(npu_inst_pe_1_4_7_N79) );
  AND2_X1 npu_inst_pe_1_4_7_U120 ( .A1(npu_inst_pe_1_4_7_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_4__7__6_), .ZN(
        npu_inst_pe_1_4_7_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_4_7_U119 ( .A(npu_inst_int_data_res_4__7__7_), .B(
        npu_inst_pe_1_4_7_add_79_carry_7_), .Z(npu_inst_pe_1_4_7_N80) );
  XNOR2_X1 npu_inst_pe_1_4_7_U118 ( .A(npu_inst_pe_1_4_7_sub_77_carry_2_), .B(
        npu_inst_int_data_res_4__7__2_), .ZN(npu_inst_pe_1_4_7_N67) );
  OR2_X1 npu_inst_pe_1_4_7_U117 ( .A1(npu_inst_int_data_res_4__7__2_), .A2(
        npu_inst_pe_1_4_7_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_4_7_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_4_7_U116 ( .A(npu_inst_pe_1_4_7_sub_77_carry_3_), .B(
        npu_inst_int_data_res_4__7__3_), .ZN(npu_inst_pe_1_4_7_N68) );
  OR2_X1 npu_inst_pe_1_4_7_U115 ( .A1(npu_inst_int_data_res_4__7__3_), .A2(
        npu_inst_pe_1_4_7_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_4_7_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_4_7_U114 ( .A(npu_inst_pe_1_4_7_sub_77_carry_4_), .B(
        npu_inst_int_data_res_4__7__4_), .ZN(npu_inst_pe_1_4_7_N69) );
  OR2_X1 npu_inst_pe_1_4_7_U113 ( .A1(npu_inst_int_data_res_4__7__4_), .A2(
        npu_inst_pe_1_4_7_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_4_7_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_4_7_U112 ( .A(npu_inst_pe_1_4_7_sub_77_carry_5_), .B(
        npu_inst_int_data_res_4__7__5_), .ZN(npu_inst_pe_1_4_7_N70) );
  OR2_X1 npu_inst_pe_1_4_7_U111 ( .A1(npu_inst_int_data_res_4__7__5_), .A2(
        npu_inst_pe_1_4_7_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_4_7_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_4_7_U110 ( .A(npu_inst_pe_1_4_7_sub_77_carry_6_), .B(
        npu_inst_int_data_res_4__7__6_), .ZN(npu_inst_pe_1_4_7_N71) );
  OR2_X1 npu_inst_pe_1_4_7_U109 ( .A1(npu_inst_int_data_res_4__7__6_), .A2(
        npu_inst_pe_1_4_7_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_4_7_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_4_7_U108 ( .A(npu_inst_int_data_res_4__7__7_), .B(
        npu_inst_pe_1_4_7_sub_77_carry_7_), .ZN(npu_inst_pe_1_4_7_N72) );
  INV_X1 npu_inst_pe_1_4_7_U107 ( .A(npu_inst_n59), .ZN(npu_inst_pe_1_4_7_n6)
         );
  INV_X1 npu_inst_pe_1_4_7_U106 ( .A(npu_inst_pe_1_4_7_n6), .ZN(
        npu_inst_pe_1_4_7_n5) );
  INV_X1 npu_inst_pe_1_4_7_U105 ( .A(npu_inst_n37), .ZN(npu_inst_pe_1_4_7_n2)
         );
  AOI22_X1 npu_inst_pe_1_4_7_U104 ( .A1(npu_inst_int_data_y_5__7__0_), .A2(
        npu_inst_pe_1_4_7_n58), .B1(npu_inst_pe_1_4_7_n118), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_4_7_n57) );
  INV_X1 npu_inst_pe_1_4_7_U103 ( .A(npu_inst_pe_1_4_7_n57), .ZN(
        npu_inst_pe_1_4_7_n107) );
  AOI22_X1 npu_inst_pe_1_4_7_U102 ( .A1(npu_inst_int_data_y_5__7__0_), .A2(
        npu_inst_pe_1_4_7_n54), .B1(npu_inst_pe_1_4_7_n117), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_4_7_n53) );
  INV_X1 npu_inst_pe_1_4_7_U99 ( .A(npu_inst_pe_1_4_7_n53), .ZN(
        npu_inst_pe_1_4_7_n108) );
  AOI22_X1 npu_inst_pe_1_4_7_U98 ( .A1(npu_inst_int_data_y_5__7__0_), .A2(
        npu_inst_pe_1_4_7_n50), .B1(npu_inst_pe_1_4_7_n116), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_4_7_n49) );
  INV_X1 npu_inst_pe_1_4_7_U97 ( .A(npu_inst_pe_1_4_7_n49), .ZN(
        npu_inst_pe_1_4_7_n109) );
  AOI22_X1 npu_inst_pe_1_4_7_U96 ( .A1(npu_inst_int_data_y_5__7__0_), .A2(
        npu_inst_pe_1_4_7_n46), .B1(npu_inst_pe_1_4_7_n115), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_4_7_n45) );
  INV_X1 npu_inst_pe_1_4_7_U95 ( .A(npu_inst_pe_1_4_7_n45), .ZN(
        npu_inst_pe_1_4_7_n110) );
  AOI22_X1 npu_inst_pe_1_4_7_U94 ( .A1(npu_inst_int_data_y_5__7__0_), .A2(
        npu_inst_pe_1_4_7_n42), .B1(npu_inst_pe_1_4_7_n114), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_4_7_n41) );
  INV_X1 npu_inst_pe_1_4_7_U93 ( .A(npu_inst_pe_1_4_7_n41), .ZN(
        npu_inst_pe_1_4_7_n111) );
  AOI22_X1 npu_inst_pe_1_4_7_U92 ( .A1(npu_inst_int_data_y_5__7__1_), .A2(
        npu_inst_pe_1_4_7_n58), .B1(npu_inst_pe_1_4_7_n118), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_4_7_n59) );
  INV_X1 npu_inst_pe_1_4_7_U91 ( .A(npu_inst_pe_1_4_7_n59), .ZN(
        npu_inst_pe_1_4_7_n101) );
  AOI22_X1 npu_inst_pe_1_4_7_U90 ( .A1(npu_inst_int_data_y_5__7__1_), .A2(
        npu_inst_pe_1_4_7_n54), .B1(npu_inst_pe_1_4_7_n117), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_4_7_n55) );
  INV_X1 npu_inst_pe_1_4_7_U89 ( .A(npu_inst_pe_1_4_7_n55), .ZN(
        npu_inst_pe_1_4_7_n102) );
  AOI22_X1 npu_inst_pe_1_4_7_U88 ( .A1(npu_inst_int_data_y_5__7__1_), .A2(
        npu_inst_pe_1_4_7_n50), .B1(npu_inst_pe_1_4_7_n116), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_4_7_n51) );
  INV_X1 npu_inst_pe_1_4_7_U87 ( .A(npu_inst_pe_1_4_7_n51), .ZN(
        npu_inst_pe_1_4_7_n103) );
  AOI22_X1 npu_inst_pe_1_4_7_U86 ( .A1(npu_inst_int_data_y_5__7__1_), .A2(
        npu_inst_pe_1_4_7_n46), .B1(npu_inst_pe_1_4_7_n115), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_4_7_n47) );
  INV_X1 npu_inst_pe_1_4_7_U85 ( .A(npu_inst_pe_1_4_7_n47), .ZN(
        npu_inst_pe_1_4_7_n104) );
  AOI22_X1 npu_inst_pe_1_4_7_U84 ( .A1(npu_inst_int_data_y_5__7__1_), .A2(
        npu_inst_pe_1_4_7_n42), .B1(npu_inst_pe_1_4_7_n114), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_4_7_n43) );
  INV_X1 npu_inst_pe_1_4_7_U83 ( .A(npu_inst_pe_1_4_7_n43), .ZN(
        npu_inst_pe_1_4_7_n105) );
  AOI22_X1 npu_inst_pe_1_4_7_U82 ( .A1(npu_inst_pe_1_4_7_n38), .A2(
        npu_inst_int_data_y_5__7__1_), .B1(npu_inst_pe_1_4_7_n113), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_4_7_n39) );
  INV_X1 npu_inst_pe_1_4_7_U81 ( .A(npu_inst_pe_1_4_7_n39), .ZN(
        npu_inst_pe_1_4_7_n106) );
  AND2_X1 npu_inst_pe_1_4_7_U80 ( .A1(npu_inst_pe_1_4_7_N93), .A2(npu_inst_n37), .ZN(npu_inst_int_data_y_4__7__0_) );
  AOI22_X1 npu_inst_pe_1_4_7_U79 ( .A1(npu_inst_pe_1_4_7_n38), .A2(
        npu_inst_int_data_y_5__7__0_), .B1(npu_inst_pe_1_4_7_n113), .B2(
        npu_inst_pe_1_4_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_4_7_n37) );
  INV_X1 npu_inst_pe_1_4_7_U78 ( .A(npu_inst_pe_1_4_7_n37), .ZN(
        npu_inst_pe_1_4_7_n112) );
  AND2_X1 npu_inst_pe_1_4_7_U77 ( .A1(npu_inst_n37), .A2(npu_inst_pe_1_4_7_N94), .ZN(npu_inst_int_data_y_4__7__1_) );
  AOI222_X1 npu_inst_pe_1_4_7_U76 ( .A1(npu_inst_int_data_res_5__7__0_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N73), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N65), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n84) );
  INV_X1 npu_inst_pe_1_4_7_U75 ( .A(npu_inst_pe_1_4_7_n84), .ZN(
        npu_inst_pe_1_4_7_n100) );
  AOI222_X1 npu_inst_pe_1_4_7_U74 ( .A1(npu_inst_pe_1_4_7_n1), .A2(
        npu_inst_int_data_res_5__7__7_), .B1(npu_inst_pe_1_4_7_N80), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N72), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n75) );
  INV_X1 npu_inst_pe_1_4_7_U73 ( .A(npu_inst_pe_1_4_7_n75), .ZN(
        npu_inst_pe_1_4_7_n32) );
  AOI222_X1 npu_inst_pe_1_4_7_U72 ( .A1(npu_inst_int_data_res_5__7__1_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N74), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N66), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n83) );
  INV_X1 npu_inst_pe_1_4_7_U71 ( .A(npu_inst_pe_1_4_7_n83), .ZN(
        npu_inst_pe_1_4_7_n99) );
  AOI222_X1 npu_inst_pe_1_4_7_U70 ( .A1(npu_inst_int_data_res_5__7__3_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N76), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N68), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n81) );
  INV_X1 npu_inst_pe_1_4_7_U69 ( .A(npu_inst_pe_1_4_7_n81), .ZN(
        npu_inst_pe_1_4_7_n36) );
  AOI222_X1 npu_inst_pe_1_4_7_U68 ( .A1(npu_inst_int_data_res_5__7__4_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N77), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N69), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n80) );
  INV_X1 npu_inst_pe_1_4_7_U67 ( .A(npu_inst_pe_1_4_7_n80), .ZN(
        npu_inst_pe_1_4_7_n35) );
  AOI222_X1 npu_inst_pe_1_4_7_U66 ( .A1(npu_inst_int_data_res_5__7__5_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N78), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N70), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n79) );
  INV_X1 npu_inst_pe_1_4_7_U65 ( .A(npu_inst_pe_1_4_7_n79), .ZN(
        npu_inst_pe_1_4_7_n34) );
  AOI222_X1 npu_inst_pe_1_4_7_U64 ( .A1(npu_inst_int_data_res_5__7__6_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N79), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N71), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n78) );
  INV_X1 npu_inst_pe_1_4_7_U63 ( .A(npu_inst_pe_1_4_7_n78), .ZN(
        npu_inst_pe_1_4_7_n33) );
  AND2_X1 npu_inst_pe_1_4_7_U62 ( .A1(npu_inst_int_data_x_4__7__1_), .A2(
        npu_inst_pe_1_4_7_int_q_weight_1_), .ZN(npu_inst_pe_1_4_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_4_7_U61 ( .A1(npu_inst_int_data_x_4__7__0_), .A2(
        npu_inst_pe_1_4_7_int_q_weight_1_), .ZN(npu_inst_pe_1_4_7_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_4_7_U60 ( .A(npu_inst_pe_1_4_7_int_data_1_), .ZN(
        npu_inst_pe_1_4_7_n13) );
  NAND2_X1 npu_inst_pe_1_4_7_U59 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_4_7_n60), .ZN(npu_inst_pe_1_4_7_n74) );
  OAI21_X1 npu_inst_pe_1_4_7_U58 ( .B1(npu_inst_pe_1_4_7_n63), .B2(
        npu_inst_pe_1_4_7_n60), .A(npu_inst_pe_1_4_7_n74), .ZN(
        npu_inst_pe_1_4_7_n97) );
  NAND2_X1 npu_inst_pe_1_4_7_U57 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_4_7_n60), .ZN(npu_inst_pe_1_4_7_n73) );
  OAI21_X1 npu_inst_pe_1_4_7_U56 ( .B1(npu_inst_pe_1_4_7_n61), .B2(
        npu_inst_pe_1_4_7_n60), .A(npu_inst_pe_1_4_7_n73), .ZN(
        npu_inst_pe_1_4_7_n96) );
  NAND2_X1 npu_inst_pe_1_4_7_U55 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_4_7_n56), .ZN(npu_inst_pe_1_4_7_n72) );
  OAI21_X1 npu_inst_pe_1_4_7_U54 ( .B1(npu_inst_pe_1_4_7_n63), .B2(
        npu_inst_pe_1_4_7_n56), .A(npu_inst_pe_1_4_7_n72), .ZN(
        npu_inst_pe_1_4_7_n95) );
  NAND2_X1 npu_inst_pe_1_4_7_U53 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_4_7_n56), .ZN(npu_inst_pe_1_4_7_n71) );
  OAI21_X1 npu_inst_pe_1_4_7_U52 ( .B1(npu_inst_pe_1_4_7_n61), .B2(
        npu_inst_pe_1_4_7_n56), .A(npu_inst_pe_1_4_7_n71), .ZN(
        npu_inst_pe_1_4_7_n94) );
  NAND2_X1 npu_inst_pe_1_4_7_U51 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_4_7_n52), .ZN(npu_inst_pe_1_4_7_n70) );
  OAI21_X1 npu_inst_pe_1_4_7_U50 ( .B1(npu_inst_pe_1_4_7_n63), .B2(
        npu_inst_pe_1_4_7_n52), .A(npu_inst_pe_1_4_7_n70), .ZN(
        npu_inst_pe_1_4_7_n93) );
  NAND2_X1 npu_inst_pe_1_4_7_U49 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_4_7_n52), .ZN(npu_inst_pe_1_4_7_n69) );
  OAI21_X1 npu_inst_pe_1_4_7_U48 ( .B1(npu_inst_pe_1_4_7_n61), .B2(
        npu_inst_pe_1_4_7_n52), .A(npu_inst_pe_1_4_7_n69), .ZN(
        npu_inst_pe_1_4_7_n92) );
  NAND2_X1 npu_inst_pe_1_4_7_U47 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_4_7_n48), .ZN(npu_inst_pe_1_4_7_n68) );
  OAI21_X1 npu_inst_pe_1_4_7_U46 ( .B1(npu_inst_pe_1_4_7_n63), .B2(
        npu_inst_pe_1_4_7_n48), .A(npu_inst_pe_1_4_7_n68), .ZN(
        npu_inst_pe_1_4_7_n91) );
  NAND2_X1 npu_inst_pe_1_4_7_U45 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_4_7_n48), .ZN(npu_inst_pe_1_4_7_n67) );
  OAI21_X1 npu_inst_pe_1_4_7_U44 ( .B1(npu_inst_pe_1_4_7_n61), .B2(
        npu_inst_pe_1_4_7_n48), .A(npu_inst_pe_1_4_7_n67), .ZN(
        npu_inst_pe_1_4_7_n90) );
  NAND2_X1 npu_inst_pe_1_4_7_U43 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_4_7_n44), .ZN(npu_inst_pe_1_4_7_n66) );
  OAI21_X1 npu_inst_pe_1_4_7_U42 ( .B1(npu_inst_pe_1_4_7_n63), .B2(
        npu_inst_pe_1_4_7_n44), .A(npu_inst_pe_1_4_7_n66), .ZN(
        npu_inst_pe_1_4_7_n89) );
  NAND2_X1 npu_inst_pe_1_4_7_U41 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_4_7_n44), .ZN(npu_inst_pe_1_4_7_n65) );
  OAI21_X1 npu_inst_pe_1_4_7_U40 ( .B1(npu_inst_pe_1_4_7_n61), .B2(
        npu_inst_pe_1_4_7_n44), .A(npu_inst_pe_1_4_7_n65), .ZN(
        npu_inst_pe_1_4_7_n88) );
  NAND2_X1 npu_inst_pe_1_4_7_U39 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_4_7_n40), .ZN(npu_inst_pe_1_4_7_n64) );
  OAI21_X1 npu_inst_pe_1_4_7_U38 ( .B1(npu_inst_pe_1_4_7_n63), .B2(
        npu_inst_pe_1_4_7_n40), .A(npu_inst_pe_1_4_7_n64), .ZN(
        npu_inst_pe_1_4_7_n87) );
  NAND2_X1 npu_inst_pe_1_4_7_U37 ( .A1(npu_inst_pe_1_4_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_4_7_n40), .ZN(npu_inst_pe_1_4_7_n62) );
  OAI21_X1 npu_inst_pe_1_4_7_U36 ( .B1(npu_inst_pe_1_4_7_n61), .B2(
        npu_inst_pe_1_4_7_n40), .A(npu_inst_pe_1_4_7_n62), .ZN(
        npu_inst_pe_1_4_7_n86) );
  NOR3_X1 npu_inst_pe_1_4_7_U35 ( .A1(npu_inst_pe_1_4_7_n26), .A2(npu_inst_n37), .A3(npu_inst_int_ckg[24]), .ZN(npu_inst_pe_1_4_7_n85) );
  OR2_X1 npu_inst_pe_1_4_7_U34 ( .A1(npu_inst_pe_1_4_7_n85), .A2(
        npu_inst_pe_1_4_7_n1), .ZN(npu_inst_pe_1_4_7_N84) );
  AOI222_X1 npu_inst_pe_1_4_7_U33 ( .A1(npu_inst_int_data_res_5__7__2_), .A2(
        npu_inst_pe_1_4_7_n1), .B1(npu_inst_pe_1_4_7_N75), .B2(
        npu_inst_pe_1_4_7_n76), .C1(npu_inst_pe_1_4_7_N67), .C2(
        npu_inst_pe_1_4_7_n77), .ZN(npu_inst_pe_1_4_7_n82) );
  INV_X1 npu_inst_pe_1_4_7_U32 ( .A(npu_inst_pe_1_4_7_n82), .ZN(
        npu_inst_pe_1_4_7_n98) );
  INV_X1 npu_inst_pe_1_4_7_U31 ( .A(npu_inst_pe_1_4_7_int_data_0_), .ZN(
        npu_inst_pe_1_4_7_n12) );
  INV_X1 npu_inst_pe_1_4_7_U30 ( .A(npu_inst_n51), .ZN(npu_inst_pe_1_4_7_n4)
         );
  AOI22_X1 npu_inst_pe_1_4_7_U29 ( .A1(npu_inst_n37), .A2(
        npu_inst_int_data_y_5__7__1_), .B1(npu_inst_pe_1_4_7_n2), .B2(
        int_i_data_h_npu[7]), .ZN(npu_inst_pe_1_4_7_n63) );
  AOI22_X1 npu_inst_pe_1_4_7_U28 ( .A1(npu_inst_n37), .A2(
        npu_inst_int_data_y_5__7__0_), .B1(npu_inst_pe_1_4_7_n2), .B2(
        int_i_data_h_npu[6]), .ZN(npu_inst_pe_1_4_7_n61) );
  OR3_X1 npu_inst_pe_1_4_7_U27 ( .A1(npu_inst_pe_1_4_7_n5), .A2(
        npu_inst_pe_1_4_7_n7), .A3(npu_inst_pe_1_4_7_n4), .ZN(
        npu_inst_pe_1_4_7_n56) );
  OR3_X1 npu_inst_pe_1_4_7_U26 ( .A1(npu_inst_pe_1_4_7_n4), .A2(
        npu_inst_pe_1_4_7_n7), .A3(npu_inst_pe_1_4_7_n6), .ZN(
        npu_inst_pe_1_4_7_n48) );
  INV_X1 npu_inst_pe_1_4_7_U25 ( .A(npu_inst_pe_1_4_7_n4), .ZN(
        npu_inst_pe_1_4_7_n3) );
  OR3_X1 npu_inst_pe_1_4_7_U24 ( .A1(npu_inst_pe_1_4_7_n3), .A2(
        npu_inst_pe_1_4_7_n7), .A3(npu_inst_pe_1_4_7_n6), .ZN(
        npu_inst_pe_1_4_7_n52) );
  OR3_X1 npu_inst_pe_1_4_7_U23 ( .A1(npu_inst_pe_1_4_7_n5), .A2(
        npu_inst_pe_1_4_7_n7), .A3(npu_inst_pe_1_4_7_n3), .ZN(
        npu_inst_pe_1_4_7_n60) );
  BUF_X1 npu_inst_pe_1_4_7_U22 ( .A(npu_inst_n19), .Z(npu_inst_pe_1_4_7_n1) );
  NOR2_X1 npu_inst_pe_1_4_7_U21 ( .A1(npu_inst_pe_1_4_7_n60), .A2(
        npu_inst_pe_1_4_7_n2), .ZN(npu_inst_pe_1_4_7_n58) );
  NOR2_X1 npu_inst_pe_1_4_7_U20 ( .A1(npu_inst_pe_1_4_7_n56), .A2(
        npu_inst_pe_1_4_7_n2), .ZN(npu_inst_pe_1_4_7_n54) );
  NOR2_X1 npu_inst_pe_1_4_7_U19 ( .A1(npu_inst_pe_1_4_7_n52), .A2(
        npu_inst_pe_1_4_7_n2), .ZN(npu_inst_pe_1_4_7_n50) );
  NOR2_X1 npu_inst_pe_1_4_7_U18 ( .A1(npu_inst_pe_1_4_7_n48), .A2(
        npu_inst_pe_1_4_7_n2), .ZN(npu_inst_pe_1_4_7_n46) );
  NOR2_X1 npu_inst_pe_1_4_7_U17 ( .A1(npu_inst_pe_1_4_7_n40), .A2(
        npu_inst_pe_1_4_7_n2), .ZN(npu_inst_pe_1_4_7_n38) );
  NOR2_X1 npu_inst_pe_1_4_7_U16 ( .A1(npu_inst_pe_1_4_7_n44), .A2(
        npu_inst_pe_1_4_7_n2), .ZN(npu_inst_pe_1_4_7_n42) );
  BUF_X1 npu_inst_pe_1_4_7_U15 ( .A(npu_inst_n80), .Z(npu_inst_pe_1_4_7_n7) );
  INV_X1 npu_inst_pe_1_4_7_U14 ( .A(npu_inst_n106), .ZN(npu_inst_pe_1_4_7_n11)
         );
  INV_X1 npu_inst_pe_1_4_7_U13 ( .A(npu_inst_pe_1_4_7_n38), .ZN(
        npu_inst_pe_1_4_7_n113) );
  INV_X1 npu_inst_pe_1_4_7_U12 ( .A(npu_inst_pe_1_4_7_n58), .ZN(
        npu_inst_pe_1_4_7_n118) );
  INV_X1 npu_inst_pe_1_4_7_U11 ( .A(npu_inst_pe_1_4_7_n54), .ZN(
        npu_inst_pe_1_4_7_n117) );
  INV_X1 npu_inst_pe_1_4_7_U10 ( .A(npu_inst_pe_1_4_7_n50), .ZN(
        npu_inst_pe_1_4_7_n116) );
  INV_X1 npu_inst_pe_1_4_7_U9 ( .A(npu_inst_pe_1_4_7_n46), .ZN(
        npu_inst_pe_1_4_7_n115) );
  INV_X1 npu_inst_pe_1_4_7_U8 ( .A(npu_inst_pe_1_4_7_n42), .ZN(
        npu_inst_pe_1_4_7_n114) );
  BUF_X1 npu_inst_pe_1_4_7_U7 ( .A(npu_inst_pe_1_4_7_n11), .Z(
        npu_inst_pe_1_4_7_n10) );
  BUF_X1 npu_inst_pe_1_4_7_U6 ( .A(npu_inst_pe_1_4_7_n11), .Z(
        npu_inst_pe_1_4_7_n9) );
  BUF_X1 npu_inst_pe_1_4_7_U5 ( .A(npu_inst_pe_1_4_7_n11), .Z(
        npu_inst_pe_1_4_7_n8) );
  NOR2_X1 npu_inst_pe_1_4_7_U4 ( .A1(npu_inst_pe_1_4_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_4_7_n1), .ZN(npu_inst_pe_1_4_7_n76) );
  NOR2_X1 npu_inst_pe_1_4_7_U3 ( .A1(npu_inst_pe_1_4_7_n27), .A2(
        npu_inst_pe_1_4_7_n1), .ZN(npu_inst_pe_1_4_7_n77) );
  FA_X1 npu_inst_pe_1_4_7_sub_77_U2_1 ( .A(npu_inst_int_data_res_4__7__1_), 
        .B(npu_inst_pe_1_4_7_n13), .CI(npu_inst_pe_1_4_7_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_4_7_sub_77_carry_2_), .S(npu_inst_pe_1_4_7_N66) );
  FA_X1 npu_inst_pe_1_4_7_add_79_U1_1 ( .A(npu_inst_int_data_res_4__7__1_), 
        .B(npu_inst_pe_1_4_7_int_data_1_), .CI(
        npu_inst_pe_1_4_7_add_79_carry_1_), .CO(
        npu_inst_pe_1_4_7_add_79_carry_2_), .S(npu_inst_pe_1_4_7_N74) );
  NAND3_X1 npu_inst_pe_1_4_7_U101 ( .A1(npu_inst_pe_1_4_7_n4), .A2(
        npu_inst_pe_1_4_7_n6), .A3(npu_inst_pe_1_4_7_n7), .ZN(
        npu_inst_pe_1_4_7_n44) );
  NAND3_X1 npu_inst_pe_1_4_7_U100 ( .A1(npu_inst_pe_1_4_7_n3), .A2(
        npu_inst_pe_1_4_7_n6), .A3(npu_inst_pe_1_4_7_n7), .ZN(
        npu_inst_pe_1_4_7_n40) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_4_7_n33), .CK(
        npu_inst_pe_1_4_7_net3581), .RN(npu_inst_pe_1_4_7_n8), .Q(
        npu_inst_int_data_res_4__7__6_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_4_7_n34), .CK(
        npu_inst_pe_1_4_7_net3581), .RN(npu_inst_pe_1_4_7_n8), .Q(
        npu_inst_int_data_res_4__7__5_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_4_7_n35), .CK(
        npu_inst_pe_1_4_7_net3581), .RN(npu_inst_pe_1_4_7_n8), .Q(
        npu_inst_int_data_res_4__7__4_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_4_7_n36), .CK(
        npu_inst_pe_1_4_7_net3581), .RN(npu_inst_pe_1_4_7_n8), .Q(
        npu_inst_int_data_res_4__7__3_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_4_7_n98), .CK(
        npu_inst_pe_1_4_7_net3581), .RN(npu_inst_pe_1_4_7_n8), .Q(
        npu_inst_int_data_res_4__7__2_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_4_7_n99), .CK(
        npu_inst_pe_1_4_7_net3581), .RN(npu_inst_pe_1_4_7_n8), .Q(
        npu_inst_int_data_res_4__7__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_4_7_n32), .CK(
        npu_inst_pe_1_4_7_net3581), .RN(npu_inst_pe_1_4_7_n8), .Q(
        npu_inst_int_data_res_4__7__7_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_4_7_n100), 
        .CK(npu_inst_pe_1_4_7_net3581), .RN(npu_inst_pe_1_4_7_n8), .Q(
        npu_inst_int_data_res_4__7__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_weight_reg_0_ ( .D(npu_inst_n92), .CK(
        npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n8), .Q(
        npu_inst_pe_1_4_7_int_q_weight_0_), .QN(npu_inst_pe_1_4_7_n27) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_weight_reg_1_ ( .D(npu_inst_n98), .CK(
        npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n8), .Q(
        npu_inst_pe_1_4_7_int_q_weight_1_), .QN(npu_inst_pe_1_4_7_n26) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_4_7_n112), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n8), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_4_7_n106), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n8), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_4_7_n111), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_4_7_n105), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_4_7_n110), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_4_7_n104), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_4_7_n109), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_4_7_n103), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_4_7_n108), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_4_7_n102), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_4_7_n107), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_4_7_n101), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_4_7_n86), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_4_7_n87), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n9), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_4_7_n88), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_4_7_n89), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_4_7_n90), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_4_7_n91), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_4_7_n92), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_4_7_n93), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_4_7_n94), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_4_7_n95), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_4_7_n96), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_4_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_4_7_n97), 
        .CK(npu_inst_pe_1_4_7_net3587), .RN(npu_inst_pe_1_4_7_n10), .Q(
        npu_inst_pe_1_4_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_4_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_4_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_4_7_net3581) );
  CLKGATETST_X1 npu_inst_pe_1_4_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n45), .SE(1'b0), .GCK(npu_inst_pe_1_4_7_net3587) );
  MUX2_X1 npu_inst_pe_1_5_0_U152 ( .A(npu_inst_pe_1_5_0_n30), .B(
        npu_inst_pe_1_5_0_n25), .S(npu_inst_pe_1_5_0_n6), .Z(
        npu_inst_pe_1_5_0_N93) );
  MUX2_X1 npu_inst_pe_1_5_0_U151 ( .A(npu_inst_pe_1_5_0_n29), .B(
        npu_inst_pe_1_5_0_n28), .S(npu_inst_n58), .Z(npu_inst_pe_1_5_0_n30) );
  MUX2_X1 npu_inst_pe_1_5_0_U150 ( .A(npu_inst_pe_1_5_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_0_n3), .Z(
        npu_inst_pe_1_5_0_n29) );
  MUX2_X1 npu_inst_pe_1_5_0_U149 ( .A(npu_inst_pe_1_5_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_0_n3), .Z(
        npu_inst_pe_1_5_0_n28) );
  MUX2_X1 npu_inst_pe_1_5_0_U148 ( .A(npu_inst_pe_1_5_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_0_n3), .Z(
        npu_inst_pe_1_5_0_n25) );
  MUX2_X1 npu_inst_pe_1_5_0_U147 ( .A(npu_inst_pe_1_5_0_n24), .B(
        npu_inst_pe_1_5_0_n21), .S(npu_inst_pe_1_5_0_n6), .Z(
        npu_inst_pe_1_5_0_N94) );
  MUX2_X1 npu_inst_pe_1_5_0_U146 ( .A(npu_inst_pe_1_5_0_n23), .B(
        npu_inst_pe_1_5_0_n22), .S(npu_inst_n58), .Z(npu_inst_pe_1_5_0_n24) );
  MUX2_X1 npu_inst_pe_1_5_0_U145 ( .A(npu_inst_pe_1_5_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_0_n3), .Z(
        npu_inst_pe_1_5_0_n23) );
  MUX2_X1 npu_inst_pe_1_5_0_U144 ( .A(npu_inst_pe_1_5_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_0_n3), .Z(
        npu_inst_pe_1_5_0_n22) );
  MUX2_X1 npu_inst_pe_1_5_0_U143 ( .A(npu_inst_pe_1_5_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_0_n3), .Z(
        npu_inst_pe_1_5_0_n21) );
  MUX2_X1 npu_inst_pe_1_5_0_U142 ( .A(npu_inst_pe_1_5_0_n20), .B(
        npu_inst_pe_1_5_0_n17), .S(npu_inst_pe_1_5_0_n6), .Z(
        npu_inst_pe_1_5_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_5_0_U141 ( .A(npu_inst_pe_1_5_0_n19), .B(
        npu_inst_pe_1_5_0_n18), .S(npu_inst_n58), .Z(npu_inst_pe_1_5_0_n20) );
  MUX2_X1 npu_inst_pe_1_5_0_U140 ( .A(npu_inst_pe_1_5_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_0_n3), .Z(
        npu_inst_pe_1_5_0_n19) );
  MUX2_X1 npu_inst_pe_1_5_0_U139 ( .A(npu_inst_pe_1_5_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_0_n3), .Z(
        npu_inst_pe_1_5_0_n18) );
  MUX2_X1 npu_inst_pe_1_5_0_U138 ( .A(npu_inst_pe_1_5_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_0_n3), .Z(
        npu_inst_pe_1_5_0_n17) );
  MUX2_X1 npu_inst_pe_1_5_0_U137 ( .A(npu_inst_pe_1_5_0_n16), .B(
        npu_inst_pe_1_5_0_n13), .S(npu_inst_pe_1_5_0_n6), .Z(
        npu_inst_pe_1_5_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_5_0_U136 ( .A(npu_inst_pe_1_5_0_n15), .B(
        npu_inst_pe_1_5_0_n14), .S(npu_inst_n58), .Z(npu_inst_pe_1_5_0_n16) );
  MUX2_X1 npu_inst_pe_1_5_0_U135 ( .A(npu_inst_pe_1_5_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_0_n3), .Z(
        npu_inst_pe_1_5_0_n15) );
  MUX2_X1 npu_inst_pe_1_5_0_U134 ( .A(npu_inst_pe_1_5_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_0_n3), .Z(
        npu_inst_pe_1_5_0_n14) );
  MUX2_X1 npu_inst_pe_1_5_0_U133 ( .A(npu_inst_pe_1_5_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_0_n3), .Z(
        npu_inst_pe_1_5_0_n13) );
  XOR2_X1 npu_inst_pe_1_5_0_U132 ( .A(npu_inst_pe_1_5_0_int_data_0_), .B(
        npu_inst_int_data_res_5__0__0_), .Z(npu_inst_pe_1_5_0_N73) );
  AND2_X1 npu_inst_pe_1_5_0_U131 ( .A1(npu_inst_int_data_res_5__0__0_), .A2(
        npu_inst_pe_1_5_0_int_data_0_), .ZN(npu_inst_pe_1_5_0_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_0_U130 ( .A(npu_inst_int_data_res_5__0__0_), .B(
        npu_inst_pe_1_5_0_n11), .ZN(npu_inst_pe_1_5_0_N65) );
  OR2_X1 npu_inst_pe_1_5_0_U129 ( .A1(npu_inst_pe_1_5_0_n11), .A2(
        npu_inst_int_data_res_5__0__0_), .ZN(npu_inst_pe_1_5_0_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_0_U128 ( .A(npu_inst_int_data_res_5__0__2_), .B(
        npu_inst_pe_1_5_0_add_79_carry_2_), .Z(npu_inst_pe_1_5_0_N75) );
  AND2_X1 npu_inst_pe_1_5_0_U127 ( .A1(npu_inst_pe_1_5_0_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_5__0__2_), .ZN(
        npu_inst_pe_1_5_0_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_0_U126 ( .A(npu_inst_int_data_res_5__0__3_), .B(
        npu_inst_pe_1_5_0_add_79_carry_3_), .Z(npu_inst_pe_1_5_0_N76) );
  AND2_X1 npu_inst_pe_1_5_0_U125 ( .A1(npu_inst_pe_1_5_0_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_5__0__3_), .ZN(
        npu_inst_pe_1_5_0_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_0_U124 ( .A(npu_inst_int_data_res_5__0__4_), .B(
        npu_inst_pe_1_5_0_add_79_carry_4_), .Z(npu_inst_pe_1_5_0_N77) );
  AND2_X1 npu_inst_pe_1_5_0_U123 ( .A1(npu_inst_pe_1_5_0_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_5__0__4_), .ZN(
        npu_inst_pe_1_5_0_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_0_U122 ( .A(npu_inst_int_data_res_5__0__5_), .B(
        npu_inst_pe_1_5_0_add_79_carry_5_), .Z(npu_inst_pe_1_5_0_N78) );
  AND2_X1 npu_inst_pe_1_5_0_U121 ( .A1(npu_inst_pe_1_5_0_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_5__0__5_), .ZN(
        npu_inst_pe_1_5_0_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_0_U120 ( .A(npu_inst_int_data_res_5__0__6_), .B(
        npu_inst_pe_1_5_0_add_79_carry_6_), .Z(npu_inst_pe_1_5_0_N79) );
  AND2_X1 npu_inst_pe_1_5_0_U119 ( .A1(npu_inst_pe_1_5_0_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_5__0__6_), .ZN(
        npu_inst_pe_1_5_0_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_0_U118 ( .A(npu_inst_int_data_res_5__0__7_), .B(
        npu_inst_pe_1_5_0_add_79_carry_7_), .Z(npu_inst_pe_1_5_0_N80) );
  XNOR2_X1 npu_inst_pe_1_5_0_U117 ( .A(npu_inst_pe_1_5_0_sub_77_carry_2_), .B(
        npu_inst_int_data_res_5__0__2_), .ZN(npu_inst_pe_1_5_0_N67) );
  OR2_X1 npu_inst_pe_1_5_0_U116 ( .A1(npu_inst_int_data_res_5__0__2_), .A2(
        npu_inst_pe_1_5_0_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_5_0_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_0_U115 ( .A(npu_inst_pe_1_5_0_sub_77_carry_3_), .B(
        npu_inst_int_data_res_5__0__3_), .ZN(npu_inst_pe_1_5_0_N68) );
  OR2_X1 npu_inst_pe_1_5_0_U114 ( .A1(npu_inst_int_data_res_5__0__3_), .A2(
        npu_inst_pe_1_5_0_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_5_0_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_0_U113 ( .A(npu_inst_pe_1_5_0_sub_77_carry_4_), .B(
        npu_inst_int_data_res_5__0__4_), .ZN(npu_inst_pe_1_5_0_N69) );
  OR2_X1 npu_inst_pe_1_5_0_U112 ( .A1(npu_inst_int_data_res_5__0__4_), .A2(
        npu_inst_pe_1_5_0_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_5_0_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_0_U111 ( .A(npu_inst_pe_1_5_0_sub_77_carry_5_), .B(
        npu_inst_int_data_res_5__0__5_), .ZN(npu_inst_pe_1_5_0_N70) );
  OR2_X1 npu_inst_pe_1_5_0_U110 ( .A1(npu_inst_int_data_res_5__0__5_), .A2(
        npu_inst_pe_1_5_0_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_5_0_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_0_U109 ( .A(npu_inst_pe_1_5_0_sub_77_carry_6_), .B(
        npu_inst_int_data_res_5__0__6_), .ZN(npu_inst_pe_1_5_0_N71) );
  OR2_X1 npu_inst_pe_1_5_0_U108 ( .A1(npu_inst_int_data_res_5__0__6_), .A2(
        npu_inst_pe_1_5_0_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_5_0_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_0_U107 ( .A(npu_inst_int_data_res_5__0__7_), .B(
        npu_inst_pe_1_5_0_sub_77_carry_7_), .ZN(npu_inst_pe_1_5_0_N72) );
  INV_X1 npu_inst_pe_1_5_0_U106 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_5_0_n5)
         );
  INV_X1 npu_inst_pe_1_5_0_U105 ( .A(npu_inst_n37), .ZN(npu_inst_pe_1_5_0_n2)
         );
  AOI22_X1 npu_inst_pe_1_5_0_U104 ( .A1(npu_inst_int_data_y_6__0__0_), .A2(
        npu_inst_pe_1_5_0_n58), .B1(npu_inst_pe_1_5_0_n117), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_0_n57) );
  INV_X1 npu_inst_pe_1_5_0_U103 ( .A(npu_inst_pe_1_5_0_n57), .ZN(
        npu_inst_pe_1_5_0_n106) );
  AOI22_X1 npu_inst_pe_1_5_0_U102 ( .A1(npu_inst_int_data_y_6__0__0_), .A2(
        npu_inst_pe_1_5_0_n54), .B1(npu_inst_pe_1_5_0_n116), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_0_n53) );
  INV_X1 npu_inst_pe_1_5_0_U99 ( .A(npu_inst_pe_1_5_0_n53), .ZN(
        npu_inst_pe_1_5_0_n107) );
  AOI22_X1 npu_inst_pe_1_5_0_U98 ( .A1(npu_inst_int_data_y_6__0__0_), .A2(
        npu_inst_pe_1_5_0_n50), .B1(npu_inst_pe_1_5_0_n115), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_0_n49) );
  INV_X1 npu_inst_pe_1_5_0_U97 ( .A(npu_inst_pe_1_5_0_n49), .ZN(
        npu_inst_pe_1_5_0_n108) );
  AOI22_X1 npu_inst_pe_1_5_0_U96 ( .A1(npu_inst_int_data_y_6__0__0_), .A2(
        npu_inst_pe_1_5_0_n46), .B1(npu_inst_pe_1_5_0_n114), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_0_n45) );
  INV_X1 npu_inst_pe_1_5_0_U95 ( .A(npu_inst_pe_1_5_0_n45), .ZN(
        npu_inst_pe_1_5_0_n109) );
  AOI22_X1 npu_inst_pe_1_5_0_U94 ( .A1(npu_inst_int_data_y_6__0__0_), .A2(
        npu_inst_pe_1_5_0_n42), .B1(npu_inst_pe_1_5_0_n113), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_0_n41) );
  INV_X1 npu_inst_pe_1_5_0_U93 ( .A(npu_inst_pe_1_5_0_n41), .ZN(
        npu_inst_pe_1_5_0_n110) );
  AOI22_X1 npu_inst_pe_1_5_0_U92 ( .A1(npu_inst_int_data_y_6__0__1_), .A2(
        npu_inst_pe_1_5_0_n58), .B1(npu_inst_pe_1_5_0_n117), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_0_n59) );
  INV_X1 npu_inst_pe_1_5_0_U91 ( .A(npu_inst_pe_1_5_0_n59), .ZN(
        npu_inst_pe_1_5_0_n100) );
  AOI22_X1 npu_inst_pe_1_5_0_U90 ( .A1(npu_inst_int_data_y_6__0__1_), .A2(
        npu_inst_pe_1_5_0_n54), .B1(npu_inst_pe_1_5_0_n116), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_0_n55) );
  INV_X1 npu_inst_pe_1_5_0_U89 ( .A(npu_inst_pe_1_5_0_n55), .ZN(
        npu_inst_pe_1_5_0_n101) );
  AOI22_X1 npu_inst_pe_1_5_0_U88 ( .A1(npu_inst_int_data_y_6__0__1_), .A2(
        npu_inst_pe_1_5_0_n50), .B1(npu_inst_pe_1_5_0_n115), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_0_n51) );
  INV_X1 npu_inst_pe_1_5_0_U87 ( .A(npu_inst_pe_1_5_0_n51), .ZN(
        npu_inst_pe_1_5_0_n102) );
  AOI22_X1 npu_inst_pe_1_5_0_U86 ( .A1(npu_inst_int_data_y_6__0__1_), .A2(
        npu_inst_pe_1_5_0_n46), .B1(npu_inst_pe_1_5_0_n114), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_0_n47) );
  INV_X1 npu_inst_pe_1_5_0_U85 ( .A(npu_inst_pe_1_5_0_n47), .ZN(
        npu_inst_pe_1_5_0_n103) );
  AOI22_X1 npu_inst_pe_1_5_0_U84 ( .A1(npu_inst_int_data_y_6__0__1_), .A2(
        npu_inst_pe_1_5_0_n42), .B1(npu_inst_pe_1_5_0_n113), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_0_n43) );
  INV_X1 npu_inst_pe_1_5_0_U83 ( .A(npu_inst_pe_1_5_0_n43), .ZN(
        npu_inst_pe_1_5_0_n104) );
  AOI22_X1 npu_inst_pe_1_5_0_U82 ( .A1(npu_inst_pe_1_5_0_n38), .A2(
        npu_inst_int_data_y_6__0__1_), .B1(npu_inst_pe_1_5_0_n112), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_0_n39) );
  INV_X1 npu_inst_pe_1_5_0_U81 ( .A(npu_inst_pe_1_5_0_n39), .ZN(
        npu_inst_pe_1_5_0_n105) );
  AND2_X1 npu_inst_pe_1_5_0_U80 ( .A1(npu_inst_pe_1_5_0_N93), .A2(npu_inst_n37), .ZN(npu_inst_int_data_y_5__0__0_) );
  NAND2_X1 npu_inst_pe_1_5_0_U79 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_0_n60), .ZN(npu_inst_pe_1_5_0_n74) );
  OAI21_X1 npu_inst_pe_1_5_0_U78 ( .B1(npu_inst_pe_1_5_0_n63), .B2(
        npu_inst_pe_1_5_0_n60), .A(npu_inst_pe_1_5_0_n74), .ZN(
        npu_inst_pe_1_5_0_n97) );
  NAND2_X1 npu_inst_pe_1_5_0_U77 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_0_n60), .ZN(npu_inst_pe_1_5_0_n73) );
  OAI21_X1 npu_inst_pe_1_5_0_U76 ( .B1(npu_inst_pe_1_5_0_n61), .B2(
        npu_inst_pe_1_5_0_n60), .A(npu_inst_pe_1_5_0_n73), .ZN(
        npu_inst_pe_1_5_0_n96) );
  NAND2_X1 npu_inst_pe_1_5_0_U75 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_0_n56), .ZN(npu_inst_pe_1_5_0_n72) );
  OAI21_X1 npu_inst_pe_1_5_0_U74 ( .B1(npu_inst_pe_1_5_0_n63), .B2(
        npu_inst_pe_1_5_0_n56), .A(npu_inst_pe_1_5_0_n72), .ZN(
        npu_inst_pe_1_5_0_n95) );
  NAND2_X1 npu_inst_pe_1_5_0_U73 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_0_n56), .ZN(npu_inst_pe_1_5_0_n71) );
  OAI21_X1 npu_inst_pe_1_5_0_U72 ( .B1(npu_inst_pe_1_5_0_n61), .B2(
        npu_inst_pe_1_5_0_n56), .A(npu_inst_pe_1_5_0_n71), .ZN(
        npu_inst_pe_1_5_0_n94) );
  NAND2_X1 npu_inst_pe_1_5_0_U71 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_0_n52), .ZN(npu_inst_pe_1_5_0_n70) );
  OAI21_X1 npu_inst_pe_1_5_0_U70 ( .B1(npu_inst_pe_1_5_0_n63), .B2(
        npu_inst_pe_1_5_0_n52), .A(npu_inst_pe_1_5_0_n70), .ZN(
        npu_inst_pe_1_5_0_n93) );
  NAND2_X1 npu_inst_pe_1_5_0_U69 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_0_n52), .ZN(npu_inst_pe_1_5_0_n69) );
  OAI21_X1 npu_inst_pe_1_5_0_U68 ( .B1(npu_inst_pe_1_5_0_n61), .B2(
        npu_inst_pe_1_5_0_n52), .A(npu_inst_pe_1_5_0_n69), .ZN(
        npu_inst_pe_1_5_0_n92) );
  NAND2_X1 npu_inst_pe_1_5_0_U67 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_0_n48), .ZN(npu_inst_pe_1_5_0_n68) );
  OAI21_X1 npu_inst_pe_1_5_0_U66 ( .B1(npu_inst_pe_1_5_0_n63), .B2(
        npu_inst_pe_1_5_0_n48), .A(npu_inst_pe_1_5_0_n68), .ZN(
        npu_inst_pe_1_5_0_n91) );
  NAND2_X1 npu_inst_pe_1_5_0_U65 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_0_n48), .ZN(npu_inst_pe_1_5_0_n67) );
  OAI21_X1 npu_inst_pe_1_5_0_U64 ( .B1(npu_inst_pe_1_5_0_n61), .B2(
        npu_inst_pe_1_5_0_n48), .A(npu_inst_pe_1_5_0_n67), .ZN(
        npu_inst_pe_1_5_0_n90) );
  NAND2_X1 npu_inst_pe_1_5_0_U63 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_0_n44), .ZN(npu_inst_pe_1_5_0_n66) );
  OAI21_X1 npu_inst_pe_1_5_0_U62 ( .B1(npu_inst_pe_1_5_0_n63), .B2(
        npu_inst_pe_1_5_0_n44), .A(npu_inst_pe_1_5_0_n66), .ZN(
        npu_inst_pe_1_5_0_n89) );
  NAND2_X1 npu_inst_pe_1_5_0_U61 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_0_n44), .ZN(npu_inst_pe_1_5_0_n65) );
  OAI21_X1 npu_inst_pe_1_5_0_U60 ( .B1(npu_inst_pe_1_5_0_n61), .B2(
        npu_inst_pe_1_5_0_n44), .A(npu_inst_pe_1_5_0_n65), .ZN(
        npu_inst_pe_1_5_0_n88) );
  NAND2_X1 npu_inst_pe_1_5_0_U59 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_0_n40), .ZN(npu_inst_pe_1_5_0_n64) );
  OAI21_X1 npu_inst_pe_1_5_0_U58 ( .B1(npu_inst_pe_1_5_0_n63), .B2(
        npu_inst_pe_1_5_0_n40), .A(npu_inst_pe_1_5_0_n64), .ZN(
        npu_inst_pe_1_5_0_n87) );
  NAND2_X1 npu_inst_pe_1_5_0_U57 ( .A1(npu_inst_pe_1_5_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_0_n40), .ZN(npu_inst_pe_1_5_0_n62) );
  OAI21_X1 npu_inst_pe_1_5_0_U56 ( .B1(npu_inst_pe_1_5_0_n61), .B2(
        npu_inst_pe_1_5_0_n40), .A(npu_inst_pe_1_5_0_n62), .ZN(
        npu_inst_pe_1_5_0_n86) );
  AOI22_X1 npu_inst_pe_1_5_0_U55 ( .A1(npu_inst_pe_1_5_0_n38), .A2(
        npu_inst_int_data_y_6__0__0_), .B1(npu_inst_pe_1_5_0_n112), .B2(
        npu_inst_pe_1_5_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_0_n37) );
  INV_X1 npu_inst_pe_1_5_0_U54 ( .A(npu_inst_pe_1_5_0_n37), .ZN(
        npu_inst_pe_1_5_0_n111) );
  AND2_X1 npu_inst_pe_1_5_0_U53 ( .A1(npu_inst_n37), .A2(npu_inst_pe_1_5_0_N94), .ZN(npu_inst_int_data_y_5__0__1_) );
  AOI222_X1 npu_inst_pe_1_5_0_U52 ( .A1(npu_inst_int_data_res_6__0__0_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N73), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N65), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n84) );
  INV_X1 npu_inst_pe_1_5_0_U51 ( .A(npu_inst_pe_1_5_0_n84), .ZN(
        npu_inst_pe_1_5_0_n99) );
  AOI222_X1 npu_inst_pe_1_5_0_U50 ( .A1(npu_inst_pe_1_5_0_n1), .A2(
        npu_inst_int_data_res_6__0__7_), .B1(npu_inst_pe_1_5_0_N80), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N72), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n75) );
  INV_X1 npu_inst_pe_1_5_0_U49 ( .A(npu_inst_pe_1_5_0_n75), .ZN(
        npu_inst_pe_1_5_0_n31) );
  AOI222_X1 npu_inst_pe_1_5_0_U48 ( .A1(npu_inst_int_data_res_6__0__1_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N74), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N66), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n83) );
  INV_X1 npu_inst_pe_1_5_0_U47 ( .A(npu_inst_pe_1_5_0_n83), .ZN(
        npu_inst_pe_1_5_0_n98) );
  AOI222_X1 npu_inst_pe_1_5_0_U46 ( .A1(npu_inst_int_data_res_6__0__3_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N76), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N68), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n81) );
  INV_X1 npu_inst_pe_1_5_0_U45 ( .A(npu_inst_pe_1_5_0_n81), .ZN(
        npu_inst_pe_1_5_0_n35) );
  AOI222_X1 npu_inst_pe_1_5_0_U44 ( .A1(npu_inst_int_data_res_6__0__4_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N77), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N69), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n80) );
  INV_X1 npu_inst_pe_1_5_0_U43 ( .A(npu_inst_pe_1_5_0_n80), .ZN(
        npu_inst_pe_1_5_0_n34) );
  AOI222_X1 npu_inst_pe_1_5_0_U42 ( .A1(npu_inst_int_data_res_6__0__5_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N78), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N70), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n79) );
  INV_X1 npu_inst_pe_1_5_0_U41 ( .A(npu_inst_pe_1_5_0_n79), .ZN(
        npu_inst_pe_1_5_0_n33) );
  AOI222_X1 npu_inst_pe_1_5_0_U40 ( .A1(npu_inst_int_data_res_6__0__6_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N79), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N71), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n78) );
  INV_X1 npu_inst_pe_1_5_0_U39 ( .A(npu_inst_pe_1_5_0_n78), .ZN(
        npu_inst_pe_1_5_0_n32) );
  NOR3_X1 npu_inst_pe_1_5_0_U38 ( .A1(npu_inst_pe_1_5_0_n26), .A2(npu_inst_n37), .A3(npu_inst_int_ckg[23]), .ZN(npu_inst_pe_1_5_0_n85) );
  OR2_X1 npu_inst_pe_1_5_0_U37 ( .A1(npu_inst_pe_1_5_0_n85), .A2(
        npu_inst_pe_1_5_0_n1), .ZN(npu_inst_pe_1_5_0_N84) );
  AND2_X1 npu_inst_pe_1_5_0_U36 ( .A1(npu_inst_pe_1_5_0_o_data_h_1_), .A2(
        npu_inst_pe_1_5_0_int_q_weight_1_), .ZN(npu_inst_pe_1_5_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_0_U35 ( .A1(npu_inst_pe_1_5_0_o_data_h_0_), .A2(
        npu_inst_pe_1_5_0_int_q_weight_1_), .ZN(npu_inst_pe_1_5_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_5_0_U34 ( .A(npu_inst_pe_1_5_0_int_data_1_), .ZN(
        npu_inst_pe_1_5_0_n12) );
  AOI222_X1 npu_inst_pe_1_5_0_U33 ( .A1(npu_inst_int_data_res_6__0__2_), .A2(
        npu_inst_pe_1_5_0_n1), .B1(npu_inst_pe_1_5_0_N75), .B2(
        npu_inst_pe_1_5_0_n76), .C1(npu_inst_pe_1_5_0_N67), .C2(
        npu_inst_pe_1_5_0_n77), .ZN(npu_inst_pe_1_5_0_n82) );
  INV_X1 npu_inst_pe_1_5_0_U32 ( .A(npu_inst_pe_1_5_0_n82), .ZN(
        npu_inst_pe_1_5_0_n36) );
  AOI22_X1 npu_inst_pe_1_5_0_U31 ( .A1(npu_inst_n37), .A2(
        npu_inst_int_data_y_6__0__1_), .B1(npu_inst_pe_1_5_0_n2), .B2(
        npu_inst_int_data_x_5__1__1_), .ZN(npu_inst_pe_1_5_0_n63) );
  AOI22_X1 npu_inst_pe_1_5_0_U30 ( .A1(npu_inst_n37), .A2(
        npu_inst_int_data_y_6__0__0_), .B1(npu_inst_pe_1_5_0_n2), .B2(
        npu_inst_int_data_x_5__1__0_), .ZN(npu_inst_pe_1_5_0_n61) );
  INV_X1 npu_inst_pe_1_5_0_U29 ( .A(npu_inst_pe_1_5_0_int_data_0_), .ZN(
        npu_inst_pe_1_5_0_n11) );
  INV_X1 npu_inst_pe_1_5_0_U28 ( .A(npu_inst_n50), .ZN(npu_inst_pe_1_5_0_n4)
         );
  OR3_X1 npu_inst_pe_1_5_0_U27 ( .A1(npu_inst_n58), .A2(npu_inst_pe_1_5_0_n6), 
        .A3(npu_inst_pe_1_5_0_n4), .ZN(npu_inst_pe_1_5_0_n56) );
  OR3_X1 npu_inst_pe_1_5_0_U26 ( .A1(npu_inst_pe_1_5_0_n4), .A2(
        npu_inst_pe_1_5_0_n6), .A3(npu_inst_pe_1_5_0_n5), .ZN(
        npu_inst_pe_1_5_0_n48) );
  INV_X1 npu_inst_pe_1_5_0_U25 ( .A(npu_inst_pe_1_5_0_n4), .ZN(
        npu_inst_pe_1_5_0_n3) );
  OR3_X1 npu_inst_pe_1_5_0_U24 ( .A1(npu_inst_pe_1_5_0_n3), .A2(
        npu_inst_pe_1_5_0_n6), .A3(npu_inst_pe_1_5_0_n5), .ZN(
        npu_inst_pe_1_5_0_n52) );
  OR3_X1 npu_inst_pe_1_5_0_U23 ( .A1(npu_inst_n58), .A2(npu_inst_pe_1_5_0_n6), 
        .A3(npu_inst_pe_1_5_0_n3), .ZN(npu_inst_pe_1_5_0_n60) );
  BUF_X1 npu_inst_pe_1_5_0_U22 ( .A(npu_inst_n18), .Z(npu_inst_pe_1_5_0_n1) );
  NOR2_X1 npu_inst_pe_1_5_0_U21 ( .A1(npu_inst_pe_1_5_0_n60), .A2(
        npu_inst_pe_1_5_0_n2), .ZN(npu_inst_pe_1_5_0_n58) );
  NOR2_X1 npu_inst_pe_1_5_0_U20 ( .A1(npu_inst_pe_1_5_0_n56), .A2(
        npu_inst_pe_1_5_0_n2), .ZN(npu_inst_pe_1_5_0_n54) );
  NOR2_X1 npu_inst_pe_1_5_0_U19 ( .A1(npu_inst_pe_1_5_0_n52), .A2(
        npu_inst_pe_1_5_0_n2), .ZN(npu_inst_pe_1_5_0_n50) );
  NOR2_X1 npu_inst_pe_1_5_0_U18 ( .A1(npu_inst_pe_1_5_0_n48), .A2(
        npu_inst_pe_1_5_0_n2), .ZN(npu_inst_pe_1_5_0_n46) );
  NOR2_X1 npu_inst_pe_1_5_0_U17 ( .A1(npu_inst_pe_1_5_0_n40), .A2(
        npu_inst_pe_1_5_0_n2), .ZN(npu_inst_pe_1_5_0_n38) );
  NOR2_X1 npu_inst_pe_1_5_0_U16 ( .A1(npu_inst_pe_1_5_0_n44), .A2(
        npu_inst_pe_1_5_0_n2), .ZN(npu_inst_pe_1_5_0_n42) );
  BUF_X1 npu_inst_pe_1_5_0_U15 ( .A(npu_inst_n79), .Z(npu_inst_pe_1_5_0_n6) );
  INV_X1 npu_inst_pe_1_5_0_U14 ( .A(npu_inst_n105), .ZN(npu_inst_pe_1_5_0_n10)
         );
  INV_X1 npu_inst_pe_1_5_0_U13 ( .A(npu_inst_pe_1_5_0_n38), .ZN(
        npu_inst_pe_1_5_0_n112) );
  INV_X1 npu_inst_pe_1_5_0_U12 ( .A(npu_inst_pe_1_5_0_n58), .ZN(
        npu_inst_pe_1_5_0_n117) );
  INV_X1 npu_inst_pe_1_5_0_U11 ( .A(npu_inst_pe_1_5_0_n54), .ZN(
        npu_inst_pe_1_5_0_n116) );
  INV_X1 npu_inst_pe_1_5_0_U10 ( .A(npu_inst_pe_1_5_0_n50), .ZN(
        npu_inst_pe_1_5_0_n115) );
  INV_X1 npu_inst_pe_1_5_0_U9 ( .A(npu_inst_pe_1_5_0_n46), .ZN(
        npu_inst_pe_1_5_0_n114) );
  INV_X1 npu_inst_pe_1_5_0_U8 ( .A(npu_inst_pe_1_5_0_n42), .ZN(
        npu_inst_pe_1_5_0_n113) );
  BUF_X1 npu_inst_pe_1_5_0_U7 ( .A(npu_inst_pe_1_5_0_n10), .Z(
        npu_inst_pe_1_5_0_n9) );
  BUF_X1 npu_inst_pe_1_5_0_U6 ( .A(npu_inst_pe_1_5_0_n10), .Z(
        npu_inst_pe_1_5_0_n8) );
  BUF_X1 npu_inst_pe_1_5_0_U5 ( .A(npu_inst_pe_1_5_0_n10), .Z(
        npu_inst_pe_1_5_0_n7) );
  NOR2_X1 npu_inst_pe_1_5_0_U4 ( .A1(npu_inst_pe_1_5_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_0_n1), .ZN(npu_inst_pe_1_5_0_n76) );
  NOR2_X1 npu_inst_pe_1_5_0_U3 ( .A1(npu_inst_pe_1_5_0_n27), .A2(
        npu_inst_pe_1_5_0_n1), .ZN(npu_inst_pe_1_5_0_n77) );
  FA_X1 npu_inst_pe_1_5_0_sub_77_U2_1 ( .A(npu_inst_int_data_res_5__0__1_), 
        .B(npu_inst_pe_1_5_0_n12), .CI(npu_inst_pe_1_5_0_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_5_0_sub_77_carry_2_), .S(npu_inst_pe_1_5_0_N66) );
  FA_X1 npu_inst_pe_1_5_0_add_79_U1_1 ( .A(npu_inst_int_data_res_5__0__1_), 
        .B(npu_inst_pe_1_5_0_int_data_1_), .CI(
        npu_inst_pe_1_5_0_add_79_carry_1_), .CO(
        npu_inst_pe_1_5_0_add_79_carry_2_), .S(npu_inst_pe_1_5_0_N74) );
  NAND3_X1 npu_inst_pe_1_5_0_U101 ( .A1(npu_inst_pe_1_5_0_n4), .A2(
        npu_inst_pe_1_5_0_n5), .A3(npu_inst_pe_1_5_0_n6), .ZN(
        npu_inst_pe_1_5_0_n44) );
  NAND3_X1 npu_inst_pe_1_5_0_U100 ( .A1(npu_inst_pe_1_5_0_n3), .A2(
        npu_inst_pe_1_5_0_n5), .A3(npu_inst_pe_1_5_0_n6), .ZN(
        npu_inst_pe_1_5_0_n40) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_0_n32), .CK(
        npu_inst_pe_1_5_0_net3558), .RN(npu_inst_pe_1_5_0_n7), .Q(
        npu_inst_int_data_res_5__0__6_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_0_n33), .CK(
        npu_inst_pe_1_5_0_net3558), .RN(npu_inst_pe_1_5_0_n7), .Q(
        npu_inst_int_data_res_5__0__5_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_0_n34), .CK(
        npu_inst_pe_1_5_0_net3558), .RN(npu_inst_pe_1_5_0_n7), .Q(
        npu_inst_int_data_res_5__0__4_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_0_n35), .CK(
        npu_inst_pe_1_5_0_net3558), .RN(npu_inst_pe_1_5_0_n7), .Q(
        npu_inst_int_data_res_5__0__3_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_0_n36), .CK(
        npu_inst_pe_1_5_0_net3558), .RN(npu_inst_pe_1_5_0_n7), .Q(
        npu_inst_int_data_res_5__0__2_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_0_n98), .CK(
        npu_inst_pe_1_5_0_net3558), .RN(npu_inst_pe_1_5_0_n7), .Q(
        npu_inst_int_data_res_5__0__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_0_n31), .CK(
        npu_inst_pe_1_5_0_net3558), .RN(npu_inst_pe_1_5_0_n7), .Q(
        npu_inst_int_data_res_5__0__7_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_0_n99), .CK(
        npu_inst_pe_1_5_0_net3558), .RN(npu_inst_pe_1_5_0_n7), .Q(
        npu_inst_int_data_res_5__0__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_weight_reg_0_ ( .D(npu_inst_n91), .CK(
        npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n7), .Q(
        npu_inst_pe_1_5_0_int_q_weight_0_), .QN(npu_inst_pe_1_5_0_n27) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_weight_reg_1_ ( .D(npu_inst_n97), .CK(
        npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n7), .Q(
        npu_inst_pe_1_5_0_int_q_weight_1_), .QN(npu_inst_pe_1_5_0_n26) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_0_n111), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n7), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_0_n105), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n7), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_0_n110), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_0_n104), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_0_n109), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_0_n103), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_0_n108), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_0_n102), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_0_n107), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_0_n101), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_0_n106), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_0_n100), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_0_n86), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_0_n87), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n8), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_0_n88), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_0_n89), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_0_n90), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_0_n91), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_0_n92), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_0_n93), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_0_n94), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_0_n95), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_0_n96), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_0_n97), 
        .CK(npu_inst_pe_1_5_0_net3564), .RN(npu_inst_pe_1_5_0_n9), .Q(
        npu_inst_pe_1_5_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_0_net3558) );
  CLKGATETST_X1 npu_inst_pe_1_5_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n45), .SE(1'b0), .GCK(npu_inst_pe_1_5_0_net3564) );
  MUX2_X1 npu_inst_pe_1_5_1_U153 ( .A(npu_inst_pe_1_5_1_n31), .B(
        npu_inst_pe_1_5_1_n28), .S(npu_inst_pe_1_5_1_n7), .Z(
        npu_inst_pe_1_5_1_N93) );
  MUX2_X1 npu_inst_pe_1_5_1_U152 ( .A(npu_inst_pe_1_5_1_n30), .B(
        npu_inst_pe_1_5_1_n29), .S(npu_inst_pe_1_5_1_n5), .Z(
        npu_inst_pe_1_5_1_n31) );
  MUX2_X1 npu_inst_pe_1_5_1_U151 ( .A(npu_inst_pe_1_5_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_1_n3), .Z(
        npu_inst_pe_1_5_1_n30) );
  MUX2_X1 npu_inst_pe_1_5_1_U150 ( .A(npu_inst_pe_1_5_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_1_n3), .Z(
        npu_inst_pe_1_5_1_n29) );
  MUX2_X1 npu_inst_pe_1_5_1_U149 ( .A(npu_inst_pe_1_5_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_1_n3), .Z(
        npu_inst_pe_1_5_1_n28) );
  MUX2_X1 npu_inst_pe_1_5_1_U148 ( .A(npu_inst_pe_1_5_1_n25), .B(
        npu_inst_pe_1_5_1_n22), .S(npu_inst_pe_1_5_1_n7), .Z(
        npu_inst_pe_1_5_1_N94) );
  MUX2_X1 npu_inst_pe_1_5_1_U147 ( .A(npu_inst_pe_1_5_1_n24), .B(
        npu_inst_pe_1_5_1_n23), .S(npu_inst_pe_1_5_1_n5), .Z(
        npu_inst_pe_1_5_1_n25) );
  MUX2_X1 npu_inst_pe_1_5_1_U146 ( .A(npu_inst_pe_1_5_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_1_n3), .Z(
        npu_inst_pe_1_5_1_n24) );
  MUX2_X1 npu_inst_pe_1_5_1_U145 ( .A(npu_inst_pe_1_5_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_1_n3), .Z(
        npu_inst_pe_1_5_1_n23) );
  MUX2_X1 npu_inst_pe_1_5_1_U144 ( .A(npu_inst_pe_1_5_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_1_n3), .Z(
        npu_inst_pe_1_5_1_n22) );
  MUX2_X1 npu_inst_pe_1_5_1_U143 ( .A(npu_inst_pe_1_5_1_n21), .B(
        npu_inst_pe_1_5_1_n18), .S(npu_inst_pe_1_5_1_n7), .Z(
        npu_inst_int_data_x_5__1__1_) );
  MUX2_X1 npu_inst_pe_1_5_1_U142 ( .A(npu_inst_pe_1_5_1_n20), .B(
        npu_inst_pe_1_5_1_n19), .S(npu_inst_pe_1_5_1_n5), .Z(
        npu_inst_pe_1_5_1_n21) );
  MUX2_X1 npu_inst_pe_1_5_1_U141 ( .A(npu_inst_pe_1_5_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_1_n3), .Z(
        npu_inst_pe_1_5_1_n20) );
  MUX2_X1 npu_inst_pe_1_5_1_U140 ( .A(npu_inst_pe_1_5_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_1_n3), .Z(
        npu_inst_pe_1_5_1_n19) );
  MUX2_X1 npu_inst_pe_1_5_1_U139 ( .A(npu_inst_pe_1_5_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_1_n3), .Z(
        npu_inst_pe_1_5_1_n18) );
  MUX2_X1 npu_inst_pe_1_5_1_U138 ( .A(npu_inst_pe_1_5_1_n17), .B(
        npu_inst_pe_1_5_1_n14), .S(npu_inst_pe_1_5_1_n7), .Z(
        npu_inst_int_data_x_5__1__0_) );
  MUX2_X1 npu_inst_pe_1_5_1_U137 ( .A(npu_inst_pe_1_5_1_n16), .B(
        npu_inst_pe_1_5_1_n15), .S(npu_inst_pe_1_5_1_n5), .Z(
        npu_inst_pe_1_5_1_n17) );
  MUX2_X1 npu_inst_pe_1_5_1_U136 ( .A(npu_inst_pe_1_5_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_1_n3), .Z(
        npu_inst_pe_1_5_1_n16) );
  MUX2_X1 npu_inst_pe_1_5_1_U135 ( .A(npu_inst_pe_1_5_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_1_n3), .Z(
        npu_inst_pe_1_5_1_n15) );
  MUX2_X1 npu_inst_pe_1_5_1_U134 ( .A(npu_inst_pe_1_5_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_1_n3), .Z(
        npu_inst_pe_1_5_1_n14) );
  XOR2_X1 npu_inst_pe_1_5_1_U133 ( .A(npu_inst_pe_1_5_1_int_data_0_), .B(
        npu_inst_int_data_res_5__1__0_), .Z(npu_inst_pe_1_5_1_N73) );
  AND2_X1 npu_inst_pe_1_5_1_U132 ( .A1(npu_inst_int_data_res_5__1__0_), .A2(
        npu_inst_pe_1_5_1_int_data_0_), .ZN(npu_inst_pe_1_5_1_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_1_U131 ( .A(npu_inst_int_data_res_5__1__0_), .B(
        npu_inst_pe_1_5_1_n12), .ZN(npu_inst_pe_1_5_1_N65) );
  OR2_X1 npu_inst_pe_1_5_1_U130 ( .A1(npu_inst_pe_1_5_1_n12), .A2(
        npu_inst_int_data_res_5__1__0_), .ZN(npu_inst_pe_1_5_1_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_1_U129 ( .A(npu_inst_int_data_res_5__1__2_), .B(
        npu_inst_pe_1_5_1_add_79_carry_2_), .Z(npu_inst_pe_1_5_1_N75) );
  AND2_X1 npu_inst_pe_1_5_1_U128 ( .A1(npu_inst_pe_1_5_1_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_5__1__2_), .ZN(
        npu_inst_pe_1_5_1_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_1_U127 ( .A(npu_inst_int_data_res_5__1__3_), .B(
        npu_inst_pe_1_5_1_add_79_carry_3_), .Z(npu_inst_pe_1_5_1_N76) );
  AND2_X1 npu_inst_pe_1_5_1_U126 ( .A1(npu_inst_pe_1_5_1_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_5__1__3_), .ZN(
        npu_inst_pe_1_5_1_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_1_U125 ( .A(npu_inst_int_data_res_5__1__4_), .B(
        npu_inst_pe_1_5_1_add_79_carry_4_), .Z(npu_inst_pe_1_5_1_N77) );
  AND2_X1 npu_inst_pe_1_5_1_U124 ( .A1(npu_inst_pe_1_5_1_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_5__1__4_), .ZN(
        npu_inst_pe_1_5_1_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_1_U123 ( .A(npu_inst_int_data_res_5__1__5_), .B(
        npu_inst_pe_1_5_1_add_79_carry_5_), .Z(npu_inst_pe_1_5_1_N78) );
  AND2_X1 npu_inst_pe_1_5_1_U122 ( .A1(npu_inst_pe_1_5_1_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_5__1__5_), .ZN(
        npu_inst_pe_1_5_1_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_1_U121 ( .A(npu_inst_int_data_res_5__1__6_), .B(
        npu_inst_pe_1_5_1_add_79_carry_6_), .Z(npu_inst_pe_1_5_1_N79) );
  AND2_X1 npu_inst_pe_1_5_1_U120 ( .A1(npu_inst_pe_1_5_1_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_5__1__6_), .ZN(
        npu_inst_pe_1_5_1_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_1_U119 ( .A(npu_inst_int_data_res_5__1__7_), .B(
        npu_inst_pe_1_5_1_add_79_carry_7_), .Z(npu_inst_pe_1_5_1_N80) );
  XNOR2_X1 npu_inst_pe_1_5_1_U118 ( .A(npu_inst_pe_1_5_1_sub_77_carry_2_), .B(
        npu_inst_int_data_res_5__1__2_), .ZN(npu_inst_pe_1_5_1_N67) );
  OR2_X1 npu_inst_pe_1_5_1_U117 ( .A1(npu_inst_int_data_res_5__1__2_), .A2(
        npu_inst_pe_1_5_1_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_5_1_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_1_U116 ( .A(npu_inst_pe_1_5_1_sub_77_carry_3_), .B(
        npu_inst_int_data_res_5__1__3_), .ZN(npu_inst_pe_1_5_1_N68) );
  OR2_X1 npu_inst_pe_1_5_1_U115 ( .A1(npu_inst_int_data_res_5__1__3_), .A2(
        npu_inst_pe_1_5_1_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_5_1_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_1_U114 ( .A(npu_inst_pe_1_5_1_sub_77_carry_4_), .B(
        npu_inst_int_data_res_5__1__4_), .ZN(npu_inst_pe_1_5_1_N69) );
  OR2_X1 npu_inst_pe_1_5_1_U113 ( .A1(npu_inst_int_data_res_5__1__4_), .A2(
        npu_inst_pe_1_5_1_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_5_1_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_1_U112 ( .A(npu_inst_pe_1_5_1_sub_77_carry_5_), .B(
        npu_inst_int_data_res_5__1__5_), .ZN(npu_inst_pe_1_5_1_N70) );
  OR2_X1 npu_inst_pe_1_5_1_U111 ( .A1(npu_inst_int_data_res_5__1__5_), .A2(
        npu_inst_pe_1_5_1_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_5_1_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_1_U110 ( .A(npu_inst_pe_1_5_1_sub_77_carry_6_), .B(
        npu_inst_int_data_res_5__1__6_), .ZN(npu_inst_pe_1_5_1_N71) );
  OR2_X1 npu_inst_pe_1_5_1_U109 ( .A1(npu_inst_int_data_res_5__1__6_), .A2(
        npu_inst_pe_1_5_1_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_5_1_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_1_U108 ( .A(npu_inst_int_data_res_5__1__7_), .B(
        npu_inst_pe_1_5_1_sub_77_carry_7_), .ZN(npu_inst_pe_1_5_1_N72) );
  INV_X1 npu_inst_pe_1_5_1_U107 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_5_1_n6)
         );
  INV_X1 npu_inst_pe_1_5_1_U106 ( .A(npu_inst_pe_1_5_1_n6), .ZN(
        npu_inst_pe_1_5_1_n5) );
  INV_X1 npu_inst_pe_1_5_1_U105 ( .A(npu_inst_n37), .ZN(npu_inst_pe_1_5_1_n2)
         );
  AOI22_X1 npu_inst_pe_1_5_1_U104 ( .A1(npu_inst_int_data_y_6__1__0_), .A2(
        npu_inst_pe_1_5_1_n58), .B1(npu_inst_pe_1_5_1_n118), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_1_n57) );
  INV_X1 npu_inst_pe_1_5_1_U103 ( .A(npu_inst_pe_1_5_1_n57), .ZN(
        npu_inst_pe_1_5_1_n107) );
  AOI22_X1 npu_inst_pe_1_5_1_U102 ( .A1(npu_inst_int_data_y_6__1__0_), .A2(
        npu_inst_pe_1_5_1_n54), .B1(npu_inst_pe_1_5_1_n117), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_1_n53) );
  INV_X1 npu_inst_pe_1_5_1_U99 ( .A(npu_inst_pe_1_5_1_n53), .ZN(
        npu_inst_pe_1_5_1_n108) );
  AOI22_X1 npu_inst_pe_1_5_1_U98 ( .A1(npu_inst_int_data_y_6__1__0_), .A2(
        npu_inst_pe_1_5_1_n50), .B1(npu_inst_pe_1_5_1_n116), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_1_n49) );
  INV_X1 npu_inst_pe_1_5_1_U97 ( .A(npu_inst_pe_1_5_1_n49), .ZN(
        npu_inst_pe_1_5_1_n109) );
  AOI22_X1 npu_inst_pe_1_5_1_U96 ( .A1(npu_inst_int_data_y_6__1__0_), .A2(
        npu_inst_pe_1_5_1_n46), .B1(npu_inst_pe_1_5_1_n115), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_1_n45) );
  INV_X1 npu_inst_pe_1_5_1_U95 ( .A(npu_inst_pe_1_5_1_n45), .ZN(
        npu_inst_pe_1_5_1_n110) );
  AOI22_X1 npu_inst_pe_1_5_1_U94 ( .A1(npu_inst_int_data_y_6__1__0_), .A2(
        npu_inst_pe_1_5_1_n42), .B1(npu_inst_pe_1_5_1_n114), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_1_n41) );
  INV_X1 npu_inst_pe_1_5_1_U93 ( .A(npu_inst_pe_1_5_1_n41), .ZN(
        npu_inst_pe_1_5_1_n111) );
  AOI22_X1 npu_inst_pe_1_5_1_U92 ( .A1(npu_inst_int_data_y_6__1__1_), .A2(
        npu_inst_pe_1_5_1_n58), .B1(npu_inst_pe_1_5_1_n118), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_1_n59) );
  INV_X1 npu_inst_pe_1_5_1_U91 ( .A(npu_inst_pe_1_5_1_n59), .ZN(
        npu_inst_pe_1_5_1_n101) );
  AOI22_X1 npu_inst_pe_1_5_1_U90 ( .A1(npu_inst_int_data_y_6__1__1_), .A2(
        npu_inst_pe_1_5_1_n54), .B1(npu_inst_pe_1_5_1_n117), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_1_n55) );
  INV_X1 npu_inst_pe_1_5_1_U89 ( .A(npu_inst_pe_1_5_1_n55), .ZN(
        npu_inst_pe_1_5_1_n102) );
  AOI22_X1 npu_inst_pe_1_5_1_U88 ( .A1(npu_inst_int_data_y_6__1__1_), .A2(
        npu_inst_pe_1_5_1_n50), .B1(npu_inst_pe_1_5_1_n116), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_1_n51) );
  INV_X1 npu_inst_pe_1_5_1_U87 ( .A(npu_inst_pe_1_5_1_n51), .ZN(
        npu_inst_pe_1_5_1_n103) );
  AOI22_X1 npu_inst_pe_1_5_1_U86 ( .A1(npu_inst_int_data_y_6__1__1_), .A2(
        npu_inst_pe_1_5_1_n46), .B1(npu_inst_pe_1_5_1_n115), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_1_n47) );
  INV_X1 npu_inst_pe_1_5_1_U85 ( .A(npu_inst_pe_1_5_1_n47), .ZN(
        npu_inst_pe_1_5_1_n104) );
  AOI22_X1 npu_inst_pe_1_5_1_U84 ( .A1(npu_inst_int_data_y_6__1__1_), .A2(
        npu_inst_pe_1_5_1_n42), .B1(npu_inst_pe_1_5_1_n114), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_1_n43) );
  INV_X1 npu_inst_pe_1_5_1_U83 ( .A(npu_inst_pe_1_5_1_n43), .ZN(
        npu_inst_pe_1_5_1_n105) );
  AOI22_X1 npu_inst_pe_1_5_1_U82 ( .A1(npu_inst_pe_1_5_1_n38), .A2(
        npu_inst_int_data_y_6__1__1_), .B1(npu_inst_pe_1_5_1_n113), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_1_n39) );
  INV_X1 npu_inst_pe_1_5_1_U81 ( .A(npu_inst_pe_1_5_1_n39), .ZN(
        npu_inst_pe_1_5_1_n106) );
  AND2_X1 npu_inst_pe_1_5_1_U80 ( .A1(npu_inst_pe_1_5_1_N93), .A2(npu_inst_n37), .ZN(npu_inst_int_data_y_5__1__0_) );
  NAND2_X1 npu_inst_pe_1_5_1_U79 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_1_n60), .ZN(npu_inst_pe_1_5_1_n74) );
  OAI21_X1 npu_inst_pe_1_5_1_U78 ( .B1(npu_inst_pe_1_5_1_n63), .B2(
        npu_inst_pe_1_5_1_n60), .A(npu_inst_pe_1_5_1_n74), .ZN(
        npu_inst_pe_1_5_1_n97) );
  NAND2_X1 npu_inst_pe_1_5_1_U77 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_1_n60), .ZN(npu_inst_pe_1_5_1_n73) );
  OAI21_X1 npu_inst_pe_1_5_1_U76 ( .B1(npu_inst_pe_1_5_1_n61), .B2(
        npu_inst_pe_1_5_1_n60), .A(npu_inst_pe_1_5_1_n73), .ZN(
        npu_inst_pe_1_5_1_n96) );
  NAND2_X1 npu_inst_pe_1_5_1_U75 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_1_n56), .ZN(npu_inst_pe_1_5_1_n72) );
  OAI21_X1 npu_inst_pe_1_5_1_U74 ( .B1(npu_inst_pe_1_5_1_n63), .B2(
        npu_inst_pe_1_5_1_n56), .A(npu_inst_pe_1_5_1_n72), .ZN(
        npu_inst_pe_1_5_1_n95) );
  NAND2_X1 npu_inst_pe_1_5_1_U73 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_1_n56), .ZN(npu_inst_pe_1_5_1_n71) );
  OAI21_X1 npu_inst_pe_1_5_1_U72 ( .B1(npu_inst_pe_1_5_1_n61), .B2(
        npu_inst_pe_1_5_1_n56), .A(npu_inst_pe_1_5_1_n71), .ZN(
        npu_inst_pe_1_5_1_n94) );
  NAND2_X1 npu_inst_pe_1_5_1_U71 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_1_n52), .ZN(npu_inst_pe_1_5_1_n70) );
  OAI21_X1 npu_inst_pe_1_5_1_U70 ( .B1(npu_inst_pe_1_5_1_n63), .B2(
        npu_inst_pe_1_5_1_n52), .A(npu_inst_pe_1_5_1_n70), .ZN(
        npu_inst_pe_1_5_1_n93) );
  NAND2_X1 npu_inst_pe_1_5_1_U69 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_1_n52), .ZN(npu_inst_pe_1_5_1_n69) );
  OAI21_X1 npu_inst_pe_1_5_1_U68 ( .B1(npu_inst_pe_1_5_1_n61), .B2(
        npu_inst_pe_1_5_1_n52), .A(npu_inst_pe_1_5_1_n69), .ZN(
        npu_inst_pe_1_5_1_n92) );
  NAND2_X1 npu_inst_pe_1_5_1_U67 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_1_n48), .ZN(npu_inst_pe_1_5_1_n68) );
  OAI21_X1 npu_inst_pe_1_5_1_U66 ( .B1(npu_inst_pe_1_5_1_n63), .B2(
        npu_inst_pe_1_5_1_n48), .A(npu_inst_pe_1_5_1_n68), .ZN(
        npu_inst_pe_1_5_1_n91) );
  NAND2_X1 npu_inst_pe_1_5_1_U65 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_1_n48), .ZN(npu_inst_pe_1_5_1_n67) );
  OAI21_X1 npu_inst_pe_1_5_1_U64 ( .B1(npu_inst_pe_1_5_1_n61), .B2(
        npu_inst_pe_1_5_1_n48), .A(npu_inst_pe_1_5_1_n67), .ZN(
        npu_inst_pe_1_5_1_n90) );
  NAND2_X1 npu_inst_pe_1_5_1_U63 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_1_n44), .ZN(npu_inst_pe_1_5_1_n66) );
  OAI21_X1 npu_inst_pe_1_5_1_U62 ( .B1(npu_inst_pe_1_5_1_n63), .B2(
        npu_inst_pe_1_5_1_n44), .A(npu_inst_pe_1_5_1_n66), .ZN(
        npu_inst_pe_1_5_1_n89) );
  NAND2_X1 npu_inst_pe_1_5_1_U61 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_1_n44), .ZN(npu_inst_pe_1_5_1_n65) );
  OAI21_X1 npu_inst_pe_1_5_1_U60 ( .B1(npu_inst_pe_1_5_1_n61), .B2(
        npu_inst_pe_1_5_1_n44), .A(npu_inst_pe_1_5_1_n65), .ZN(
        npu_inst_pe_1_5_1_n88) );
  NAND2_X1 npu_inst_pe_1_5_1_U59 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_1_n40), .ZN(npu_inst_pe_1_5_1_n64) );
  OAI21_X1 npu_inst_pe_1_5_1_U58 ( .B1(npu_inst_pe_1_5_1_n63), .B2(
        npu_inst_pe_1_5_1_n40), .A(npu_inst_pe_1_5_1_n64), .ZN(
        npu_inst_pe_1_5_1_n87) );
  NAND2_X1 npu_inst_pe_1_5_1_U57 ( .A1(npu_inst_pe_1_5_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_1_n40), .ZN(npu_inst_pe_1_5_1_n62) );
  OAI21_X1 npu_inst_pe_1_5_1_U56 ( .B1(npu_inst_pe_1_5_1_n61), .B2(
        npu_inst_pe_1_5_1_n40), .A(npu_inst_pe_1_5_1_n62), .ZN(
        npu_inst_pe_1_5_1_n86) );
  AOI22_X1 npu_inst_pe_1_5_1_U55 ( .A1(npu_inst_pe_1_5_1_n38), .A2(
        npu_inst_int_data_y_6__1__0_), .B1(npu_inst_pe_1_5_1_n113), .B2(
        npu_inst_pe_1_5_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_1_n37) );
  INV_X1 npu_inst_pe_1_5_1_U54 ( .A(npu_inst_pe_1_5_1_n37), .ZN(
        npu_inst_pe_1_5_1_n112) );
  AND2_X1 npu_inst_pe_1_5_1_U53 ( .A1(npu_inst_n37), .A2(npu_inst_pe_1_5_1_N94), .ZN(npu_inst_int_data_y_5__1__1_) );
  AOI222_X1 npu_inst_pe_1_5_1_U52 ( .A1(npu_inst_int_data_res_6__1__0_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N73), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N65), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n84) );
  INV_X1 npu_inst_pe_1_5_1_U51 ( .A(npu_inst_pe_1_5_1_n84), .ZN(
        npu_inst_pe_1_5_1_n100) );
  AOI222_X1 npu_inst_pe_1_5_1_U50 ( .A1(npu_inst_pe_1_5_1_n1), .A2(
        npu_inst_int_data_res_6__1__7_), .B1(npu_inst_pe_1_5_1_N80), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N72), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n75) );
  INV_X1 npu_inst_pe_1_5_1_U49 ( .A(npu_inst_pe_1_5_1_n75), .ZN(
        npu_inst_pe_1_5_1_n32) );
  AOI222_X1 npu_inst_pe_1_5_1_U48 ( .A1(npu_inst_int_data_res_6__1__1_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N74), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N66), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n83) );
  INV_X1 npu_inst_pe_1_5_1_U47 ( .A(npu_inst_pe_1_5_1_n83), .ZN(
        npu_inst_pe_1_5_1_n99) );
  AOI222_X1 npu_inst_pe_1_5_1_U46 ( .A1(npu_inst_int_data_res_6__1__3_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N76), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N68), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n81) );
  INV_X1 npu_inst_pe_1_5_1_U45 ( .A(npu_inst_pe_1_5_1_n81), .ZN(
        npu_inst_pe_1_5_1_n36) );
  AOI222_X1 npu_inst_pe_1_5_1_U44 ( .A1(npu_inst_int_data_res_6__1__4_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N77), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N69), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n80) );
  INV_X1 npu_inst_pe_1_5_1_U43 ( .A(npu_inst_pe_1_5_1_n80), .ZN(
        npu_inst_pe_1_5_1_n35) );
  AOI222_X1 npu_inst_pe_1_5_1_U42 ( .A1(npu_inst_int_data_res_6__1__5_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N78), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N70), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n79) );
  INV_X1 npu_inst_pe_1_5_1_U41 ( .A(npu_inst_pe_1_5_1_n79), .ZN(
        npu_inst_pe_1_5_1_n34) );
  AOI222_X1 npu_inst_pe_1_5_1_U40 ( .A1(npu_inst_int_data_res_6__1__6_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N79), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N71), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n78) );
  INV_X1 npu_inst_pe_1_5_1_U39 ( .A(npu_inst_pe_1_5_1_n78), .ZN(
        npu_inst_pe_1_5_1_n33) );
  NOR3_X1 npu_inst_pe_1_5_1_U38 ( .A1(npu_inst_pe_1_5_1_n26), .A2(npu_inst_n37), .A3(npu_inst_int_ckg[22]), .ZN(npu_inst_pe_1_5_1_n85) );
  OR2_X1 npu_inst_pe_1_5_1_U37 ( .A1(npu_inst_pe_1_5_1_n85), .A2(
        npu_inst_pe_1_5_1_n1), .ZN(npu_inst_pe_1_5_1_N84) );
  AND2_X1 npu_inst_pe_1_5_1_U36 ( .A1(npu_inst_int_data_x_5__1__1_), .A2(
        npu_inst_pe_1_5_1_int_q_weight_1_), .ZN(npu_inst_pe_1_5_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_1_U35 ( .A1(npu_inst_int_data_x_5__1__0_), .A2(
        npu_inst_pe_1_5_1_int_q_weight_1_), .ZN(npu_inst_pe_1_5_1_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_5_1_U34 ( .A(npu_inst_pe_1_5_1_int_data_1_), .ZN(
        npu_inst_pe_1_5_1_n13) );
  AOI222_X1 npu_inst_pe_1_5_1_U33 ( .A1(npu_inst_int_data_res_6__1__2_), .A2(
        npu_inst_pe_1_5_1_n1), .B1(npu_inst_pe_1_5_1_N75), .B2(
        npu_inst_pe_1_5_1_n76), .C1(npu_inst_pe_1_5_1_N67), .C2(
        npu_inst_pe_1_5_1_n77), .ZN(npu_inst_pe_1_5_1_n82) );
  INV_X1 npu_inst_pe_1_5_1_U32 ( .A(npu_inst_pe_1_5_1_n82), .ZN(
        npu_inst_pe_1_5_1_n98) );
  AOI22_X1 npu_inst_pe_1_5_1_U31 ( .A1(npu_inst_n37), .A2(
        npu_inst_int_data_y_6__1__1_), .B1(npu_inst_pe_1_5_1_n2), .B2(
        npu_inst_int_data_x_5__2__1_), .ZN(npu_inst_pe_1_5_1_n63) );
  AOI22_X1 npu_inst_pe_1_5_1_U30 ( .A1(npu_inst_n37), .A2(
        npu_inst_int_data_y_6__1__0_), .B1(npu_inst_pe_1_5_1_n2), .B2(
        npu_inst_int_data_x_5__2__0_), .ZN(npu_inst_pe_1_5_1_n61) );
  INV_X1 npu_inst_pe_1_5_1_U29 ( .A(npu_inst_pe_1_5_1_int_data_0_), .ZN(
        npu_inst_pe_1_5_1_n12) );
  INV_X1 npu_inst_pe_1_5_1_U28 ( .A(npu_inst_n50), .ZN(npu_inst_pe_1_5_1_n4)
         );
  OR3_X1 npu_inst_pe_1_5_1_U27 ( .A1(npu_inst_pe_1_5_1_n5), .A2(
        npu_inst_pe_1_5_1_n7), .A3(npu_inst_pe_1_5_1_n4), .ZN(
        npu_inst_pe_1_5_1_n56) );
  OR3_X1 npu_inst_pe_1_5_1_U26 ( .A1(npu_inst_pe_1_5_1_n4), .A2(
        npu_inst_pe_1_5_1_n7), .A3(npu_inst_pe_1_5_1_n6), .ZN(
        npu_inst_pe_1_5_1_n48) );
  INV_X1 npu_inst_pe_1_5_1_U25 ( .A(npu_inst_pe_1_5_1_n4), .ZN(
        npu_inst_pe_1_5_1_n3) );
  OR3_X1 npu_inst_pe_1_5_1_U24 ( .A1(npu_inst_pe_1_5_1_n3), .A2(
        npu_inst_pe_1_5_1_n7), .A3(npu_inst_pe_1_5_1_n6), .ZN(
        npu_inst_pe_1_5_1_n52) );
  OR3_X1 npu_inst_pe_1_5_1_U23 ( .A1(npu_inst_pe_1_5_1_n5), .A2(
        npu_inst_pe_1_5_1_n7), .A3(npu_inst_pe_1_5_1_n3), .ZN(
        npu_inst_pe_1_5_1_n60) );
  BUF_X1 npu_inst_pe_1_5_1_U22 ( .A(npu_inst_n18), .Z(npu_inst_pe_1_5_1_n1) );
  NOR2_X1 npu_inst_pe_1_5_1_U21 ( .A1(npu_inst_pe_1_5_1_n60), .A2(
        npu_inst_pe_1_5_1_n2), .ZN(npu_inst_pe_1_5_1_n58) );
  NOR2_X1 npu_inst_pe_1_5_1_U20 ( .A1(npu_inst_pe_1_5_1_n56), .A2(
        npu_inst_pe_1_5_1_n2), .ZN(npu_inst_pe_1_5_1_n54) );
  NOR2_X1 npu_inst_pe_1_5_1_U19 ( .A1(npu_inst_pe_1_5_1_n52), .A2(
        npu_inst_pe_1_5_1_n2), .ZN(npu_inst_pe_1_5_1_n50) );
  NOR2_X1 npu_inst_pe_1_5_1_U18 ( .A1(npu_inst_pe_1_5_1_n48), .A2(
        npu_inst_pe_1_5_1_n2), .ZN(npu_inst_pe_1_5_1_n46) );
  NOR2_X1 npu_inst_pe_1_5_1_U17 ( .A1(npu_inst_pe_1_5_1_n40), .A2(
        npu_inst_pe_1_5_1_n2), .ZN(npu_inst_pe_1_5_1_n38) );
  NOR2_X1 npu_inst_pe_1_5_1_U16 ( .A1(npu_inst_pe_1_5_1_n44), .A2(
        npu_inst_pe_1_5_1_n2), .ZN(npu_inst_pe_1_5_1_n42) );
  BUF_X1 npu_inst_pe_1_5_1_U15 ( .A(npu_inst_n79), .Z(npu_inst_pe_1_5_1_n7) );
  INV_X1 npu_inst_pe_1_5_1_U14 ( .A(npu_inst_n105), .ZN(npu_inst_pe_1_5_1_n11)
         );
  INV_X1 npu_inst_pe_1_5_1_U13 ( .A(npu_inst_pe_1_5_1_n38), .ZN(
        npu_inst_pe_1_5_1_n113) );
  INV_X1 npu_inst_pe_1_5_1_U12 ( .A(npu_inst_pe_1_5_1_n58), .ZN(
        npu_inst_pe_1_5_1_n118) );
  INV_X1 npu_inst_pe_1_5_1_U11 ( .A(npu_inst_pe_1_5_1_n54), .ZN(
        npu_inst_pe_1_5_1_n117) );
  INV_X1 npu_inst_pe_1_5_1_U10 ( .A(npu_inst_pe_1_5_1_n50), .ZN(
        npu_inst_pe_1_5_1_n116) );
  INV_X1 npu_inst_pe_1_5_1_U9 ( .A(npu_inst_pe_1_5_1_n46), .ZN(
        npu_inst_pe_1_5_1_n115) );
  INV_X1 npu_inst_pe_1_5_1_U8 ( .A(npu_inst_pe_1_5_1_n42), .ZN(
        npu_inst_pe_1_5_1_n114) );
  BUF_X1 npu_inst_pe_1_5_1_U7 ( .A(npu_inst_pe_1_5_1_n11), .Z(
        npu_inst_pe_1_5_1_n10) );
  BUF_X1 npu_inst_pe_1_5_1_U6 ( .A(npu_inst_pe_1_5_1_n11), .Z(
        npu_inst_pe_1_5_1_n9) );
  BUF_X1 npu_inst_pe_1_5_1_U5 ( .A(npu_inst_pe_1_5_1_n11), .Z(
        npu_inst_pe_1_5_1_n8) );
  NOR2_X1 npu_inst_pe_1_5_1_U4 ( .A1(npu_inst_pe_1_5_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_1_n1), .ZN(npu_inst_pe_1_5_1_n76) );
  NOR2_X1 npu_inst_pe_1_5_1_U3 ( .A1(npu_inst_pe_1_5_1_n27), .A2(
        npu_inst_pe_1_5_1_n1), .ZN(npu_inst_pe_1_5_1_n77) );
  FA_X1 npu_inst_pe_1_5_1_sub_77_U2_1 ( .A(npu_inst_int_data_res_5__1__1_), 
        .B(npu_inst_pe_1_5_1_n13), .CI(npu_inst_pe_1_5_1_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_5_1_sub_77_carry_2_), .S(npu_inst_pe_1_5_1_N66) );
  FA_X1 npu_inst_pe_1_5_1_add_79_U1_1 ( .A(npu_inst_int_data_res_5__1__1_), 
        .B(npu_inst_pe_1_5_1_int_data_1_), .CI(
        npu_inst_pe_1_5_1_add_79_carry_1_), .CO(
        npu_inst_pe_1_5_1_add_79_carry_2_), .S(npu_inst_pe_1_5_1_N74) );
  NAND3_X1 npu_inst_pe_1_5_1_U101 ( .A1(npu_inst_pe_1_5_1_n4), .A2(
        npu_inst_pe_1_5_1_n6), .A3(npu_inst_pe_1_5_1_n7), .ZN(
        npu_inst_pe_1_5_1_n44) );
  NAND3_X1 npu_inst_pe_1_5_1_U100 ( .A1(npu_inst_pe_1_5_1_n3), .A2(
        npu_inst_pe_1_5_1_n6), .A3(npu_inst_pe_1_5_1_n7), .ZN(
        npu_inst_pe_1_5_1_n40) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_1_n33), .CK(
        npu_inst_pe_1_5_1_net3535), .RN(npu_inst_pe_1_5_1_n8), .Q(
        npu_inst_int_data_res_5__1__6_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_1_n34), .CK(
        npu_inst_pe_1_5_1_net3535), .RN(npu_inst_pe_1_5_1_n8), .Q(
        npu_inst_int_data_res_5__1__5_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_1_n35), .CK(
        npu_inst_pe_1_5_1_net3535), .RN(npu_inst_pe_1_5_1_n8), .Q(
        npu_inst_int_data_res_5__1__4_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_1_n36), .CK(
        npu_inst_pe_1_5_1_net3535), .RN(npu_inst_pe_1_5_1_n8), .Q(
        npu_inst_int_data_res_5__1__3_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_1_n98), .CK(
        npu_inst_pe_1_5_1_net3535), .RN(npu_inst_pe_1_5_1_n8), .Q(
        npu_inst_int_data_res_5__1__2_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_1_n99), .CK(
        npu_inst_pe_1_5_1_net3535), .RN(npu_inst_pe_1_5_1_n8), .Q(
        npu_inst_int_data_res_5__1__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_1_n32), .CK(
        npu_inst_pe_1_5_1_net3535), .RN(npu_inst_pe_1_5_1_n8), .Q(
        npu_inst_int_data_res_5__1__7_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_1_n100), 
        .CK(npu_inst_pe_1_5_1_net3535), .RN(npu_inst_pe_1_5_1_n8), .Q(
        npu_inst_int_data_res_5__1__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_weight_reg_0_ ( .D(npu_inst_n91), .CK(
        npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n8), .Q(
        npu_inst_pe_1_5_1_int_q_weight_0_), .QN(npu_inst_pe_1_5_1_n27) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_weight_reg_1_ ( .D(npu_inst_n97), .CK(
        npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n8), .Q(
        npu_inst_pe_1_5_1_int_q_weight_1_), .QN(npu_inst_pe_1_5_1_n26) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_1_n112), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n8), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_1_n106), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n8), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_1_n111), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_1_n105), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_1_n110), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_1_n104), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_1_n109), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_1_n103), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_1_n108), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_1_n102), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_1_n107), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_1_n101), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_1_n86), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_1_n87), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n9), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_1_n88), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_1_n89), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_1_n90), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_1_n91), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_1_n92), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_1_n93), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_1_n94), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_1_n95), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_1_n96), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_1_n97), 
        .CK(npu_inst_pe_1_5_1_net3541), .RN(npu_inst_pe_1_5_1_n10), .Q(
        npu_inst_pe_1_5_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_1_net3535) );
  CLKGATETST_X1 npu_inst_pe_1_5_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n45), .SE(1'b0), .GCK(npu_inst_pe_1_5_1_net3541) );
  MUX2_X1 npu_inst_pe_1_5_2_U153 ( .A(npu_inst_pe_1_5_2_n31), .B(
        npu_inst_pe_1_5_2_n28), .S(npu_inst_pe_1_5_2_n7), .Z(
        npu_inst_pe_1_5_2_N93) );
  MUX2_X1 npu_inst_pe_1_5_2_U152 ( .A(npu_inst_pe_1_5_2_n30), .B(
        npu_inst_pe_1_5_2_n29), .S(npu_inst_pe_1_5_2_n5), .Z(
        npu_inst_pe_1_5_2_n31) );
  MUX2_X1 npu_inst_pe_1_5_2_U151 ( .A(npu_inst_pe_1_5_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_2_n3), .Z(
        npu_inst_pe_1_5_2_n30) );
  MUX2_X1 npu_inst_pe_1_5_2_U150 ( .A(npu_inst_pe_1_5_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_2_n3), .Z(
        npu_inst_pe_1_5_2_n29) );
  MUX2_X1 npu_inst_pe_1_5_2_U149 ( .A(npu_inst_pe_1_5_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_2_n3), .Z(
        npu_inst_pe_1_5_2_n28) );
  MUX2_X1 npu_inst_pe_1_5_2_U148 ( .A(npu_inst_pe_1_5_2_n25), .B(
        npu_inst_pe_1_5_2_n22), .S(npu_inst_pe_1_5_2_n7), .Z(
        npu_inst_pe_1_5_2_N94) );
  MUX2_X1 npu_inst_pe_1_5_2_U147 ( .A(npu_inst_pe_1_5_2_n24), .B(
        npu_inst_pe_1_5_2_n23), .S(npu_inst_pe_1_5_2_n5), .Z(
        npu_inst_pe_1_5_2_n25) );
  MUX2_X1 npu_inst_pe_1_5_2_U146 ( .A(npu_inst_pe_1_5_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_2_n3), .Z(
        npu_inst_pe_1_5_2_n24) );
  MUX2_X1 npu_inst_pe_1_5_2_U145 ( .A(npu_inst_pe_1_5_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_2_n3), .Z(
        npu_inst_pe_1_5_2_n23) );
  MUX2_X1 npu_inst_pe_1_5_2_U144 ( .A(npu_inst_pe_1_5_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_2_n3), .Z(
        npu_inst_pe_1_5_2_n22) );
  MUX2_X1 npu_inst_pe_1_5_2_U143 ( .A(npu_inst_pe_1_5_2_n21), .B(
        npu_inst_pe_1_5_2_n18), .S(npu_inst_pe_1_5_2_n7), .Z(
        npu_inst_int_data_x_5__2__1_) );
  MUX2_X1 npu_inst_pe_1_5_2_U142 ( .A(npu_inst_pe_1_5_2_n20), .B(
        npu_inst_pe_1_5_2_n19), .S(npu_inst_pe_1_5_2_n5), .Z(
        npu_inst_pe_1_5_2_n21) );
  MUX2_X1 npu_inst_pe_1_5_2_U141 ( .A(npu_inst_pe_1_5_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_2_n3), .Z(
        npu_inst_pe_1_5_2_n20) );
  MUX2_X1 npu_inst_pe_1_5_2_U140 ( .A(npu_inst_pe_1_5_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_2_n3), .Z(
        npu_inst_pe_1_5_2_n19) );
  MUX2_X1 npu_inst_pe_1_5_2_U139 ( .A(npu_inst_pe_1_5_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_2_n3), .Z(
        npu_inst_pe_1_5_2_n18) );
  MUX2_X1 npu_inst_pe_1_5_2_U138 ( .A(npu_inst_pe_1_5_2_n17), .B(
        npu_inst_pe_1_5_2_n14), .S(npu_inst_pe_1_5_2_n7), .Z(
        npu_inst_int_data_x_5__2__0_) );
  MUX2_X1 npu_inst_pe_1_5_2_U137 ( .A(npu_inst_pe_1_5_2_n16), .B(
        npu_inst_pe_1_5_2_n15), .S(npu_inst_pe_1_5_2_n5), .Z(
        npu_inst_pe_1_5_2_n17) );
  MUX2_X1 npu_inst_pe_1_5_2_U136 ( .A(npu_inst_pe_1_5_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_2_n3), .Z(
        npu_inst_pe_1_5_2_n16) );
  MUX2_X1 npu_inst_pe_1_5_2_U135 ( .A(npu_inst_pe_1_5_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_2_n3), .Z(
        npu_inst_pe_1_5_2_n15) );
  MUX2_X1 npu_inst_pe_1_5_2_U134 ( .A(npu_inst_pe_1_5_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_2_n3), .Z(
        npu_inst_pe_1_5_2_n14) );
  XOR2_X1 npu_inst_pe_1_5_2_U133 ( .A(npu_inst_pe_1_5_2_int_data_0_), .B(
        npu_inst_int_data_res_5__2__0_), .Z(npu_inst_pe_1_5_2_N73) );
  AND2_X1 npu_inst_pe_1_5_2_U132 ( .A1(npu_inst_int_data_res_5__2__0_), .A2(
        npu_inst_pe_1_5_2_int_data_0_), .ZN(npu_inst_pe_1_5_2_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_2_U131 ( .A(npu_inst_int_data_res_5__2__0_), .B(
        npu_inst_pe_1_5_2_n12), .ZN(npu_inst_pe_1_5_2_N65) );
  OR2_X1 npu_inst_pe_1_5_2_U130 ( .A1(npu_inst_pe_1_5_2_n12), .A2(
        npu_inst_int_data_res_5__2__0_), .ZN(npu_inst_pe_1_5_2_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_2_U129 ( .A(npu_inst_int_data_res_5__2__2_), .B(
        npu_inst_pe_1_5_2_add_79_carry_2_), .Z(npu_inst_pe_1_5_2_N75) );
  AND2_X1 npu_inst_pe_1_5_2_U128 ( .A1(npu_inst_pe_1_5_2_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_5__2__2_), .ZN(
        npu_inst_pe_1_5_2_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_2_U127 ( .A(npu_inst_int_data_res_5__2__3_), .B(
        npu_inst_pe_1_5_2_add_79_carry_3_), .Z(npu_inst_pe_1_5_2_N76) );
  AND2_X1 npu_inst_pe_1_5_2_U126 ( .A1(npu_inst_pe_1_5_2_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_5__2__3_), .ZN(
        npu_inst_pe_1_5_2_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_2_U125 ( .A(npu_inst_int_data_res_5__2__4_), .B(
        npu_inst_pe_1_5_2_add_79_carry_4_), .Z(npu_inst_pe_1_5_2_N77) );
  AND2_X1 npu_inst_pe_1_5_2_U124 ( .A1(npu_inst_pe_1_5_2_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_5__2__4_), .ZN(
        npu_inst_pe_1_5_2_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_2_U123 ( .A(npu_inst_int_data_res_5__2__5_), .B(
        npu_inst_pe_1_5_2_add_79_carry_5_), .Z(npu_inst_pe_1_5_2_N78) );
  AND2_X1 npu_inst_pe_1_5_2_U122 ( .A1(npu_inst_pe_1_5_2_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_5__2__5_), .ZN(
        npu_inst_pe_1_5_2_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_2_U121 ( .A(npu_inst_int_data_res_5__2__6_), .B(
        npu_inst_pe_1_5_2_add_79_carry_6_), .Z(npu_inst_pe_1_5_2_N79) );
  AND2_X1 npu_inst_pe_1_5_2_U120 ( .A1(npu_inst_pe_1_5_2_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_5__2__6_), .ZN(
        npu_inst_pe_1_5_2_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_2_U119 ( .A(npu_inst_int_data_res_5__2__7_), .B(
        npu_inst_pe_1_5_2_add_79_carry_7_), .Z(npu_inst_pe_1_5_2_N80) );
  XNOR2_X1 npu_inst_pe_1_5_2_U118 ( .A(npu_inst_pe_1_5_2_sub_77_carry_2_), .B(
        npu_inst_int_data_res_5__2__2_), .ZN(npu_inst_pe_1_5_2_N67) );
  OR2_X1 npu_inst_pe_1_5_2_U117 ( .A1(npu_inst_int_data_res_5__2__2_), .A2(
        npu_inst_pe_1_5_2_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_5_2_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_2_U116 ( .A(npu_inst_pe_1_5_2_sub_77_carry_3_), .B(
        npu_inst_int_data_res_5__2__3_), .ZN(npu_inst_pe_1_5_2_N68) );
  OR2_X1 npu_inst_pe_1_5_2_U115 ( .A1(npu_inst_int_data_res_5__2__3_), .A2(
        npu_inst_pe_1_5_2_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_5_2_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_2_U114 ( .A(npu_inst_pe_1_5_2_sub_77_carry_4_), .B(
        npu_inst_int_data_res_5__2__4_), .ZN(npu_inst_pe_1_5_2_N69) );
  OR2_X1 npu_inst_pe_1_5_2_U113 ( .A1(npu_inst_int_data_res_5__2__4_), .A2(
        npu_inst_pe_1_5_2_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_5_2_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_2_U112 ( .A(npu_inst_pe_1_5_2_sub_77_carry_5_), .B(
        npu_inst_int_data_res_5__2__5_), .ZN(npu_inst_pe_1_5_2_N70) );
  OR2_X1 npu_inst_pe_1_5_2_U111 ( .A1(npu_inst_int_data_res_5__2__5_), .A2(
        npu_inst_pe_1_5_2_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_5_2_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_2_U110 ( .A(npu_inst_pe_1_5_2_sub_77_carry_6_), .B(
        npu_inst_int_data_res_5__2__6_), .ZN(npu_inst_pe_1_5_2_N71) );
  OR2_X1 npu_inst_pe_1_5_2_U109 ( .A1(npu_inst_int_data_res_5__2__6_), .A2(
        npu_inst_pe_1_5_2_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_5_2_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_2_U108 ( .A(npu_inst_int_data_res_5__2__7_), .B(
        npu_inst_pe_1_5_2_sub_77_carry_7_), .ZN(npu_inst_pe_1_5_2_N72) );
  INV_X1 npu_inst_pe_1_5_2_U107 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_5_2_n6)
         );
  INV_X1 npu_inst_pe_1_5_2_U106 ( .A(npu_inst_pe_1_5_2_n6), .ZN(
        npu_inst_pe_1_5_2_n5) );
  INV_X1 npu_inst_pe_1_5_2_U105 ( .A(npu_inst_n37), .ZN(npu_inst_pe_1_5_2_n2)
         );
  AOI22_X1 npu_inst_pe_1_5_2_U104 ( .A1(npu_inst_int_data_y_6__2__0_), .A2(
        npu_inst_pe_1_5_2_n58), .B1(npu_inst_pe_1_5_2_n118), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_2_n57) );
  INV_X1 npu_inst_pe_1_5_2_U103 ( .A(npu_inst_pe_1_5_2_n57), .ZN(
        npu_inst_pe_1_5_2_n107) );
  AOI22_X1 npu_inst_pe_1_5_2_U102 ( .A1(npu_inst_int_data_y_6__2__0_), .A2(
        npu_inst_pe_1_5_2_n54), .B1(npu_inst_pe_1_5_2_n117), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_2_n53) );
  INV_X1 npu_inst_pe_1_5_2_U99 ( .A(npu_inst_pe_1_5_2_n53), .ZN(
        npu_inst_pe_1_5_2_n108) );
  AOI22_X1 npu_inst_pe_1_5_2_U98 ( .A1(npu_inst_int_data_y_6__2__0_), .A2(
        npu_inst_pe_1_5_2_n50), .B1(npu_inst_pe_1_5_2_n116), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_2_n49) );
  INV_X1 npu_inst_pe_1_5_2_U97 ( .A(npu_inst_pe_1_5_2_n49), .ZN(
        npu_inst_pe_1_5_2_n109) );
  AOI22_X1 npu_inst_pe_1_5_2_U96 ( .A1(npu_inst_int_data_y_6__2__0_), .A2(
        npu_inst_pe_1_5_2_n46), .B1(npu_inst_pe_1_5_2_n115), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_2_n45) );
  INV_X1 npu_inst_pe_1_5_2_U95 ( .A(npu_inst_pe_1_5_2_n45), .ZN(
        npu_inst_pe_1_5_2_n110) );
  AOI22_X1 npu_inst_pe_1_5_2_U94 ( .A1(npu_inst_int_data_y_6__2__0_), .A2(
        npu_inst_pe_1_5_2_n42), .B1(npu_inst_pe_1_5_2_n114), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_2_n41) );
  INV_X1 npu_inst_pe_1_5_2_U93 ( .A(npu_inst_pe_1_5_2_n41), .ZN(
        npu_inst_pe_1_5_2_n111) );
  AOI22_X1 npu_inst_pe_1_5_2_U92 ( .A1(npu_inst_int_data_y_6__2__1_), .A2(
        npu_inst_pe_1_5_2_n58), .B1(npu_inst_pe_1_5_2_n118), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_2_n59) );
  INV_X1 npu_inst_pe_1_5_2_U91 ( .A(npu_inst_pe_1_5_2_n59), .ZN(
        npu_inst_pe_1_5_2_n101) );
  AOI22_X1 npu_inst_pe_1_5_2_U90 ( .A1(npu_inst_int_data_y_6__2__1_), .A2(
        npu_inst_pe_1_5_2_n54), .B1(npu_inst_pe_1_5_2_n117), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_2_n55) );
  INV_X1 npu_inst_pe_1_5_2_U89 ( .A(npu_inst_pe_1_5_2_n55), .ZN(
        npu_inst_pe_1_5_2_n102) );
  AOI22_X1 npu_inst_pe_1_5_2_U88 ( .A1(npu_inst_int_data_y_6__2__1_), .A2(
        npu_inst_pe_1_5_2_n50), .B1(npu_inst_pe_1_5_2_n116), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_2_n51) );
  INV_X1 npu_inst_pe_1_5_2_U87 ( .A(npu_inst_pe_1_5_2_n51), .ZN(
        npu_inst_pe_1_5_2_n103) );
  AOI22_X1 npu_inst_pe_1_5_2_U86 ( .A1(npu_inst_int_data_y_6__2__1_), .A2(
        npu_inst_pe_1_5_2_n46), .B1(npu_inst_pe_1_5_2_n115), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_2_n47) );
  INV_X1 npu_inst_pe_1_5_2_U85 ( .A(npu_inst_pe_1_5_2_n47), .ZN(
        npu_inst_pe_1_5_2_n104) );
  AOI22_X1 npu_inst_pe_1_5_2_U84 ( .A1(npu_inst_int_data_y_6__2__1_), .A2(
        npu_inst_pe_1_5_2_n42), .B1(npu_inst_pe_1_5_2_n114), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_2_n43) );
  INV_X1 npu_inst_pe_1_5_2_U83 ( .A(npu_inst_pe_1_5_2_n43), .ZN(
        npu_inst_pe_1_5_2_n105) );
  AOI22_X1 npu_inst_pe_1_5_2_U82 ( .A1(npu_inst_pe_1_5_2_n38), .A2(
        npu_inst_int_data_y_6__2__1_), .B1(npu_inst_pe_1_5_2_n113), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_2_n39) );
  INV_X1 npu_inst_pe_1_5_2_U81 ( .A(npu_inst_pe_1_5_2_n39), .ZN(
        npu_inst_pe_1_5_2_n106) );
  AND2_X1 npu_inst_pe_1_5_2_U80 ( .A1(npu_inst_pe_1_5_2_N93), .A2(npu_inst_n37), .ZN(npu_inst_int_data_y_5__2__0_) );
  NAND2_X1 npu_inst_pe_1_5_2_U79 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_2_n60), .ZN(npu_inst_pe_1_5_2_n74) );
  OAI21_X1 npu_inst_pe_1_5_2_U78 ( .B1(npu_inst_pe_1_5_2_n63), .B2(
        npu_inst_pe_1_5_2_n60), .A(npu_inst_pe_1_5_2_n74), .ZN(
        npu_inst_pe_1_5_2_n97) );
  NAND2_X1 npu_inst_pe_1_5_2_U77 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_2_n60), .ZN(npu_inst_pe_1_5_2_n73) );
  OAI21_X1 npu_inst_pe_1_5_2_U76 ( .B1(npu_inst_pe_1_5_2_n61), .B2(
        npu_inst_pe_1_5_2_n60), .A(npu_inst_pe_1_5_2_n73), .ZN(
        npu_inst_pe_1_5_2_n96) );
  NAND2_X1 npu_inst_pe_1_5_2_U75 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_2_n56), .ZN(npu_inst_pe_1_5_2_n72) );
  OAI21_X1 npu_inst_pe_1_5_2_U74 ( .B1(npu_inst_pe_1_5_2_n63), .B2(
        npu_inst_pe_1_5_2_n56), .A(npu_inst_pe_1_5_2_n72), .ZN(
        npu_inst_pe_1_5_2_n95) );
  NAND2_X1 npu_inst_pe_1_5_2_U73 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_2_n56), .ZN(npu_inst_pe_1_5_2_n71) );
  OAI21_X1 npu_inst_pe_1_5_2_U72 ( .B1(npu_inst_pe_1_5_2_n61), .B2(
        npu_inst_pe_1_5_2_n56), .A(npu_inst_pe_1_5_2_n71), .ZN(
        npu_inst_pe_1_5_2_n94) );
  NAND2_X1 npu_inst_pe_1_5_2_U71 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_2_n52), .ZN(npu_inst_pe_1_5_2_n70) );
  OAI21_X1 npu_inst_pe_1_5_2_U70 ( .B1(npu_inst_pe_1_5_2_n63), .B2(
        npu_inst_pe_1_5_2_n52), .A(npu_inst_pe_1_5_2_n70), .ZN(
        npu_inst_pe_1_5_2_n93) );
  NAND2_X1 npu_inst_pe_1_5_2_U69 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_2_n52), .ZN(npu_inst_pe_1_5_2_n69) );
  OAI21_X1 npu_inst_pe_1_5_2_U68 ( .B1(npu_inst_pe_1_5_2_n61), .B2(
        npu_inst_pe_1_5_2_n52), .A(npu_inst_pe_1_5_2_n69), .ZN(
        npu_inst_pe_1_5_2_n92) );
  NAND2_X1 npu_inst_pe_1_5_2_U67 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_2_n48), .ZN(npu_inst_pe_1_5_2_n68) );
  OAI21_X1 npu_inst_pe_1_5_2_U66 ( .B1(npu_inst_pe_1_5_2_n63), .B2(
        npu_inst_pe_1_5_2_n48), .A(npu_inst_pe_1_5_2_n68), .ZN(
        npu_inst_pe_1_5_2_n91) );
  NAND2_X1 npu_inst_pe_1_5_2_U65 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_2_n48), .ZN(npu_inst_pe_1_5_2_n67) );
  OAI21_X1 npu_inst_pe_1_5_2_U64 ( .B1(npu_inst_pe_1_5_2_n61), .B2(
        npu_inst_pe_1_5_2_n48), .A(npu_inst_pe_1_5_2_n67), .ZN(
        npu_inst_pe_1_5_2_n90) );
  NAND2_X1 npu_inst_pe_1_5_2_U63 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_2_n44), .ZN(npu_inst_pe_1_5_2_n66) );
  OAI21_X1 npu_inst_pe_1_5_2_U62 ( .B1(npu_inst_pe_1_5_2_n63), .B2(
        npu_inst_pe_1_5_2_n44), .A(npu_inst_pe_1_5_2_n66), .ZN(
        npu_inst_pe_1_5_2_n89) );
  NAND2_X1 npu_inst_pe_1_5_2_U61 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_2_n44), .ZN(npu_inst_pe_1_5_2_n65) );
  OAI21_X1 npu_inst_pe_1_5_2_U60 ( .B1(npu_inst_pe_1_5_2_n61), .B2(
        npu_inst_pe_1_5_2_n44), .A(npu_inst_pe_1_5_2_n65), .ZN(
        npu_inst_pe_1_5_2_n88) );
  NAND2_X1 npu_inst_pe_1_5_2_U59 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_2_n40), .ZN(npu_inst_pe_1_5_2_n64) );
  OAI21_X1 npu_inst_pe_1_5_2_U58 ( .B1(npu_inst_pe_1_5_2_n63), .B2(
        npu_inst_pe_1_5_2_n40), .A(npu_inst_pe_1_5_2_n64), .ZN(
        npu_inst_pe_1_5_2_n87) );
  NAND2_X1 npu_inst_pe_1_5_2_U57 ( .A1(npu_inst_pe_1_5_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_2_n40), .ZN(npu_inst_pe_1_5_2_n62) );
  OAI21_X1 npu_inst_pe_1_5_2_U56 ( .B1(npu_inst_pe_1_5_2_n61), .B2(
        npu_inst_pe_1_5_2_n40), .A(npu_inst_pe_1_5_2_n62), .ZN(
        npu_inst_pe_1_5_2_n86) );
  AOI22_X1 npu_inst_pe_1_5_2_U55 ( .A1(npu_inst_pe_1_5_2_n38), .A2(
        npu_inst_int_data_y_6__2__0_), .B1(npu_inst_pe_1_5_2_n113), .B2(
        npu_inst_pe_1_5_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_2_n37) );
  INV_X1 npu_inst_pe_1_5_2_U54 ( .A(npu_inst_pe_1_5_2_n37), .ZN(
        npu_inst_pe_1_5_2_n112) );
  AND2_X1 npu_inst_pe_1_5_2_U53 ( .A1(npu_inst_n37), .A2(npu_inst_pe_1_5_2_N94), .ZN(npu_inst_int_data_y_5__2__1_) );
  AOI222_X1 npu_inst_pe_1_5_2_U52 ( .A1(npu_inst_int_data_res_6__2__0_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N73), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N65), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n84) );
  INV_X1 npu_inst_pe_1_5_2_U51 ( .A(npu_inst_pe_1_5_2_n84), .ZN(
        npu_inst_pe_1_5_2_n100) );
  AOI222_X1 npu_inst_pe_1_5_2_U50 ( .A1(npu_inst_pe_1_5_2_n1), .A2(
        npu_inst_int_data_res_6__2__7_), .B1(npu_inst_pe_1_5_2_N80), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N72), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n75) );
  INV_X1 npu_inst_pe_1_5_2_U49 ( .A(npu_inst_pe_1_5_2_n75), .ZN(
        npu_inst_pe_1_5_2_n32) );
  AOI222_X1 npu_inst_pe_1_5_2_U48 ( .A1(npu_inst_int_data_res_6__2__1_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N74), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N66), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n83) );
  INV_X1 npu_inst_pe_1_5_2_U47 ( .A(npu_inst_pe_1_5_2_n83), .ZN(
        npu_inst_pe_1_5_2_n99) );
  AOI222_X1 npu_inst_pe_1_5_2_U46 ( .A1(npu_inst_int_data_res_6__2__3_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N76), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N68), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n81) );
  INV_X1 npu_inst_pe_1_5_2_U45 ( .A(npu_inst_pe_1_5_2_n81), .ZN(
        npu_inst_pe_1_5_2_n36) );
  AOI222_X1 npu_inst_pe_1_5_2_U44 ( .A1(npu_inst_int_data_res_6__2__4_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N77), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N69), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n80) );
  INV_X1 npu_inst_pe_1_5_2_U43 ( .A(npu_inst_pe_1_5_2_n80), .ZN(
        npu_inst_pe_1_5_2_n35) );
  AOI222_X1 npu_inst_pe_1_5_2_U42 ( .A1(npu_inst_int_data_res_6__2__5_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N78), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N70), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n79) );
  INV_X1 npu_inst_pe_1_5_2_U41 ( .A(npu_inst_pe_1_5_2_n79), .ZN(
        npu_inst_pe_1_5_2_n34) );
  AOI222_X1 npu_inst_pe_1_5_2_U40 ( .A1(npu_inst_int_data_res_6__2__6_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N79), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N71), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n78) );
  INV_X1 npu_inst_pe_1_5_2_U39 ( .A(npu_inst_pe_1_5_2_n78), .ZN(
        npu_inst_pe_1_5_2_n33) );
  NOR3_X1 npu_inst_pe_1_5_2_U38 ( .A1(npu_inst_pe_1_5_2_n26), .A2(npu_inst_n37), .A3(npu_inst_int_ckg[21]), .ZN(npu_inst_pe_1_5_2_n85) );
  OR2_X1 npu_inst_pe_1_5_2_U37 ( .A1(npu_inst_pe_1_5_2_n85), .A2(
        npu_inst_pe_1_5_2_n1), .ZN(npu_inst_pe_1_5_2_N84) );
  AND2_X1 npu_inst_pe_1_5_2_U36 ( .A1(npu_inst_int_data_x_5__2__1_), .A2(
        npu_inst_pe_1_5_2_int_q_weight_1_), .ZN(npu_inst_pe_1_5_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_2_U35 ( .A1(npu_inst_int_data_x_5__2__0_), .A2(
        npu_inst_pe_1_5_2_int_q_weight_1_), .ZN(npu_inst_pe_1_5_2_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_5_2_U34 ( .A(npu_inst_pe_1_5_2_int_data_1_), .ZN(
        npu_inst_pe_1_5_2_n13) );
  AOI222_X1 npu_inst_pe_1_5_2_U33 ( .A1(npu_inst_int_data_res_6__2__2_), .A2(
        npu_inst_pe_1_5_2_n1), .B1(npu_inst_pe_1_5_2_N75), .B2(
        npu_inst_pe_1_5_2_n76), .C1(npu_inst_pe_1_5_2_N67), .C2(
        npu_inst_pe_1_5_2_n77), .ZN(npu_inst_pe_1_5_2_n82) );
  INV_X1 npu_inst_pe_1_5_2_U32 ( .A(npu_inst_pe_1_5_2_n82), .ZN(
        npu_inst_pe_1_5_2_n98) );
  AOI22_X1 npu_inst_pe_1_5_2_U31 ( .A1(npu_inst_n37), .A2(
        npu_inst_int_data_y_6__2__1_), .B1(npu_inst_pe_1_5_2_n2), .B2(
        npu_inst_int_data_x_5__3__1_), .ZN(npu_inst_pe_1_5_2_n63) );
  AOI22_X1 npu_inst_pe_1_5_2_U30 ( .A1(npu_inst_n37), .A2(
        npu_inst_int_data_y_6__2__0_), .B1(npu_inst_pe_1_5_2_n2), .B2(
        npu_inst_int_data_x_5__3__0_), .ZN(npu_inst_pe_1_5_2_n61) );
  INV_X1 npu_inst_pe_1_5_2_U29 ( .A(npu_inst_pe_1_5_2_int_data_0_), .ZN(
        npu_inst_pe_1_5_2_n12) );
  INV_X1 npu_inst_pe_1_5_2_U28 ( .A(npu_inst_n50), .ZN(npu_inst_pe_1_5_2_n4)
         );
  OR3_X1 npu_inst_pe_1_5_2_U27 ( .A1(npu_inst_pe_1_5_2_n5), .A2(
        npu_inst_pe_1_5_2_n7), .A3(npu_inst_pe_1_5_2_n4), .ZN(
        npu_inst_pe_1_5_2_n56) );
  OR3_X1 npu_inst_pe_1_5_2_U26 ( .A1(npu_inst_pe_1_5_2_n4), .A2(
        npu_inst_pe_1_5_2_n7), .A3(npu_inst_pe_1_5_2_n6), .ZN(
        npu_inst_pe_1_5_2_n48) );
  INV_X1 npu_inst_pe_1_5_2_U25 ( .A(npu_inst_pe_1_5_2_n4), .ZN(
        npu_inst_pe_1_5_2_n3) );
  OR3_X1 npu_inst_pe_1_5_2_U24 ( .A1(npu_inst_pe_1_5_2_n3), .A2(
        npu_inst_pe_1_5_2_n7), .A3(npu_inst_pe_1_5_2_n6), .ZN(
        npu_inst_pe_1_5_2_n52) );
  OR3_X1 npu_inst_pe_1_5_2_U23 ( .A1(npu_inst_pe_1_5_2_n5), .A2(
        npu_inst_pe_1_5_2_n7), .A3(npu_inst_pe_1_5_2_n3), .ZN(
        npu_inst_pe_1_5_2_n60) );
  BUF_X1 npu_inst_pe_1_5_2_U22 ( .A(npu_inst_n18), .Z(npu_inst_pe_1_5_2_n1) );
  NOR2_X1 npu_inst_pe_1_5_2_U21 ( .A1(npu_inst_pe_1_5_2_n60), .A2(
        npu_inst_pe_1_5_2_n2), .ZN(npu_inst_pe_1_5_2_n58) );
  NOR2_X1 npu_inst_pe_1_5_2_U20 ( .A1(npu_inst_pe_1_5_2_n56), .A2(
        npu_inst_pe_1_5_2_n2), .ZN(npu_inst_pe_1_5_2_n54) );
  NOR2_X1 npu_inst_pe_1_5_2_U19 ( .A1(npu_inst_pe_1_5_2_n52), .A2(
        npu_inst_pe_1_5_2_n2), .ZN(npu_inst_pe_1_5_2_n50) );
  NOR2_X1 npu_inst_pe_1_5_2_U18 ( .A1(npu_inst_pe_1_5_2_n48), .A2(
        npu_inst_pe_1_5_2_n2), .ZN(npu_inst_pe_1_5_2_n46) );
  NOR2_X1 npu_inst_pe_1_5_2_U17 ( .A1(npu_inst_pe_1_5_2_n40), .A2(
        npu_inst_pe_1_5_2_n2), .ZN(npu_inst_pe_1_5_2_n38) );
  NOR2_X1 npu_inst_pe_1_5_2_U16 ( .A1(npu_inst_pe_1_5_2_n44), .A2(
        npu_inst_pe_1_5_2_n2), .ZN(npu_inst_pe_1_5_2_n42) );
  BUF_X1 npu_inst_pe_1_5_2_U15 ( .A(npu_inst_n79), .Z(npu_inst_pe_1_5_2_n7) );
  INV_X1 npu_inst_pe_1_5_2_U14 ( .A(npu_inst_n105), .ZN(npu_inst_pe_1_5_2_n11)
         );
  INV_X1 npu_inst_pe_1_5_2_U13 ( .A(npu_inst_pe_1_5_2_n38), .ZN(
        npu_inst_pe_1_5_2_n113) );
  INV_X1 npu_inst_pe_1_5_2_U12 ( .A(npu_inst_pe_1_5_2_n58), .ZN(
        npu_inst_pe_1_5_2_n118) );
  INV_X1 npu_inst_pe_1_5_2_U11 ( .A(npu_inst_pe_1_5_2_n54), .ZN(
        npu_inst_pe_1_5_2_n117) );
  INV_X1 npu_inst_pe_1_5_2_U10 ( .A(npu_inst_pe_1_5_2_n50), .ZN(
        npu_inst_pe_1_5_2_n116) );
  INV_X1 npu_inst_pe_1_5_2_U9 ( .A(npu_inst_pe_1_5_2_n46), .ZN(
        npu_inst_pe_1_5_2_n115) );
  INV_X1 npu_inst_pe_1_5_2_U8 ( .A(npu_inst_pe_1_5_2_n42), .ZN(
        npu_inst_pe_1_5_2_n114) );
  BUF_X1 npu_inst_pe_1_5_2_U7 ( .A(npu_inst_pe_1_5_2_n11), .Z(
        npu_inst_pe_1_5_2_n10) );
  BUF_X1 npu_inst_pe_1_5_2_U6 ( .A(npu_inst_pe_1_5_2_n11), .Z(
        npu_inst_pe_1_5_2_n9) );
  BUF_X1 npu_inst_pe_1_5_2_U5 ( .A(npu_inst_pe_1_5_2_n11), .Z(
        npu_inst_pe_1_5_2_n8) );
  NOR2_X1 npu_inst_pe_1_5_2_U4 ( .A1(npu_inst_pe_1_5_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_2_n1), .ZN(npu_inst_pe_1_5_2_n76) );
  NOR2_X1 npu_inst_pe_1_5_2_U3 ( .A1(npu_inst_pe_1_5_2_n27), .A2(
        npu_inst_pe_1_5_2_n1), .ZN(npu_inst_pe_1_5_2_n77) );
  FA_X1 npu_inst_pe_1_5_2_sub_77_U2_1 ( .A(npu_inst_int_data_res_5__2__1_), 
        .B(npu_inst_pe_1_5_2_n13), .CI(npu_inst_pe_1_5_2_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_5_2_sub_77_carry_2_), .S(npu_inst_pe_1_5_2_N66) );
  FA_X1 npu_inst_pe_1_5_2_add_79_U1_1 ( .A(npu_inst_int_data_res_5__2__1_), 
        .B(npu_inst_pe_1_5_2_int_data_1_), .CI(
        npu_inst_pe_1_5_2_add_79_carry_1_), .CO(
        npu_inst_pe_1_5_2_add_79_carry_2_), .S(npu_inst_pe_1_5_2_N74) );
  NAND3_X1 npu_inst_pe_1_5_2_U101 ( .A1(npu_inst_pe_1_5_2_n4), .A2(
        npu_inst_pe_1_5_2_n6), .A3(npu_inst_pe_1_5_2_n7), .ZN(
        npu_inst_pe_1_5_2_n44) );
  NAND3_X1 npu_inst_pe_1_5_2_U100 ( .A1(npu_inst_pe_1_5_2_n3), .A2(
        npu_inst_pe_1_5_2_n6), .A3(npu_inst_pe_1_5_2_n7), .ZN(
        npu_inst_pe_1_5_2_n40) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_2_n33), .CK(
        npu_inst_pe_1_5_2_net3512), .RN(npu_inst_pe_1_5_2_n8), .Q(
        npu_inst_int_data_res_5__2__6_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_2_n34), .CK(
        npu_inst_pe_1_5_2_net3512), .RN(npu_inst_pe_1_5_2_n8), .Q(
        npu_inst_int_data_res_5__2__5_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_2_n35), .CK(
        npu_inst_pe_1_5_2_net3512), .RN(npu_inst_pe_1_5_2_n8), .Q(
        npu_inst_int_data_res_5__2__4_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_2_n36), .CK(
        npu_inst_pe_1_5_2_net3512), .RN(npu_inst_pe_1_5_2_n8), .Q(
        npu_inst_int_data_res_5__2__3_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_2_n98), .CK(
        npu_inst_pe_1_5_2_net3512), .RN(npu_inst_pe_1_5_2_n8), .Q(
        npu_inst_int_data_res_5__2__2_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_2_n99), .CK(
        npu_inst_pe_1_5_2_net3512), .RN(npu_inst_pe_1_5_2_n8), .Q(
        npu_inst_int_data_res_5__2__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_2_n32), .CK(
        npu_inst_pe_1_5_2_net3512), .RN(npu_inst_pe_1_5_2_n8), .Q(
        npu_inst_int_data_res_5__2__7_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_2_n100), 
        .CK(npu_inst_pe_1_5_2_net3512), .RN(npu_inst_pe_1_5_2_n8), .Q(
        npu_inst_int_data_res_5__2__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_weight_reg_0_ ( .D(npu_inst_n91), .CK(
        npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n8), .Q(
        npu_inst_pe_1_5_2_int_q_weight_0_), .QN(npu_inst_pe_1_5_2_n27) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_weight_reg_1_ ( .D(npu_inst_n97), .CK(
        npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n8), .Q(
        npu_inst_pe_1_5_2_int_q_weight_1_), .QN(npu_inst_pe_1_5_2_n26) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_2_n112), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n8), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_2_n106), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n8), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_2_n111), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_2_n105), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_2_n110), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_2_n104), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_2_n109), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_2_n103), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_2_n108), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_2_n102), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_2_n107), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_2_n101), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_2_n86), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_2_n87), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n9), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_2_n88), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_2_n89), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_2_n90), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_2_n91), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_2_n92), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_2_n93), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_2_n94), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_2_n95), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_2_n96), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_2_n97), 
        .CK(npu_inst_pe_1_5_2_net3518), .RN(npu_inst_pe_1_5_2_n10), .Q(
        npu_inst_pe_1_5_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_2_net3512) );
  CLKGATETST_X1 npu_inst_pe_1_5_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n44), .SE(1'b0), .GCK(npu_inst_pe_1_5_2_net3518) );
  MUX2_X1 npu_inst_pe_1_5_3_U153 ( .A(npu_inst_pe_1_5_3_n31), .B(
        npu_inst_pe_1_5_3_n28), .S(npu_inst_pe_1_5_3_n7), .Z(
        npu_inst_pe_1_5_3_N93) );
  MUX2_X1 npu_inst_pe_1_5_3_U152 ( .A(npu_inst_pe_1_5_3_n30), .B(
        npu_inst_pe_1_5_3_n29), .S(npu_inst_pe_1_5_3_n5), .Z(
        npu_inst_pe_1_5_3_n31) );
  MUX2_X1 npu_inst_pe_1_5_3_U151 ( .A(npu_inst_pe_1_5_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_3_n3), .Z(
        npu_inst_pe_1_5_3_n30) );
  MUX2_X1 npu_inst_pe_1_5_3_U150 ( .A(npu_inst_pe_1_5_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_3_n3), .Z(
        npu_inst_pe_1_5_3_n29) );
  MUX2_X1 npu_inst_pe_1_5_3_U149 ( .A(npu_inst_pe_1_5_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_3_n3), .Z(
        npu_inst_pe_1_5_3_n28) );
  MUX2_X1 npu_inst_pe_1_5_3_U148 ( .A(npu_inst_pe_1_5_3_n25), .B(
        npu_inst_pe_1_5_3_n22), .S(npu_inst_pe_1_5_3_n7), .Z(
        npu_inst_pe_1_5_3_N94) );
  MUX2_X1 npu_inst_pe_1_5_3_U147 ( .A(npu_inst_pe_1_5_3_n24), .B(
        npu_inst_pe_1_5_3_n23), .S(npu_inst_pe_1_5_3_n5), .Z(
        npu_inst_pe_1_5_3_n25) );
  MUX2_X1 npu_inst_pe_1_5_3_U146 ( .A(npu_inst_pe_1_5_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_3_n3), .Z(
        npu_inst_pe_1_5_3_n24) );
  MUX2_X1 npu_inst_pe_1_5_3_U145 ( .A(npu_inst_pe_1_5_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_3_n3), .Z(
        npu_inst_pe_1_5_3_n23) );
  MUX2_X1 npu_inst_pe_1_5_3_U144 ( .A(npu_inst_pe_1_5_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_3_n3), .Z(
        npu_inst_pe_1_5_3_n22) );
  MUX2_X1 npu_inst_pe_1_5_3_U143 ( .A(npu_inst_pe_1_5_3_n21), .B(
        npu_inst_pe_1_5_3_n18), .S(npu_inst_pe_1_5_3_n7), .Z(
        npu_inst_int_data_x_5__3__1_) );
  MUX2_X1 npu_inst_pe_1_5_3_U142 ( .A(npu_inst_pe_1_5_3_n20), .B(
        npu_inst_pe_1_5_3_n19), .S(npu_inst_pe_1_5_3_n5), .Z(
        npu_inst_pe_1_5_3_n21) );
  MUX2_X1 npu_inst_pe_1_5_3_U141 ( .A(npu_inst_pe_1_5_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_3_n3), .Z(
        npu_inst_pe_1_5_3_n20) );
  MUX2_X1 npu_inst_pe_1_5_3_U140 ( .A(npu_inst_pe_1_5_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_3_n3), .Z(
        npu_inst_pe_1_5_3_n19) );
  MUX2_X1 npu_inst_pe_1_5_3_U139 ( .A(npu_inst_pe_1_5_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_3_n3), .Z(
        npu_inst_pe_1_5_3_n18) );
  MUX2_X1 npu_inst_pe_1_5_3_U138 ( .A(npu_inst_pe_1_5_3_n17), .B(
        npu_inst_pe_1_5_3_n14), .S(npu_inst_pe_1_5_3_n7), .Z(
        npu_inst_int_data_x_5__3__0_) );
  MUX2_X1 npu_inst_pe_1_5_3_U137 ( .A(npu_inst_pe_1_5_3_n16), .B(
        npu_inst_pe_1_5_3_n15), .S(npu_inst_pe_1_5_3_n5), .Z(
        npu_inst_pe_1_5_3_n17) );
  MUX2_X1 npu_inst_pe_1_5_3_U136 ( .A(npu_inst_pe_1_5_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_3_n3), .Z(
        npu_inst_pe_1_5_3_n16) );
  MUX2_X1 npu_inst_pe_1_5_3_U135 ( .A(npu_inst_pe_1_5_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_3_n3), .Z(
        npu_inst_pe_1_5_3_n15) );
  MUX2_X1 npu_inst_pe_1_5_3_U134 ( .A(npu_inst_pe_1_5_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_3_n3), .Z(
        npu_inst_pe_1_5_3_n14) );
  XOR2_X1 npu_inst_pe_1_5_3_U133 ( .A(npu_inst_pe_1_5_3_int_data_0_), .B(
        npu_inst_int_data_res_5__3__0_), .Z(npu_inst_pe_1_5_3_N73) );
  AND2_X1 npu_inst_pe_1_5_3_U132 ( .A1(npu_inst_int_data_res_5__3__0_), .A2(
        npu_inst_pe_1_5_3_int_data_0_), .ZN(npu_inst_pe_1_5_3_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_3_U131 ( .A(npu_inst_int_data_res_5__3__0_), .B(
        npu_inst_pe_1_5_3_n12), .ZN(npu_inst_pe_1_5_3_N65) );
  OR2_X1 npu_inst_pe_1_5_3_U130 ( .A1(npu_inst_pe_1_5_3_n12), .A2(
        npu_inst_int_data_res_5__3__0_), .ZN(npu_inst_pe_1_5_3_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_3_U129 ( .A(npu_inst_int_data_res_5__3__2_), .B(
        npu_inst_pe_1_5_3_add_79_carry_2_), .Z(npu_inst_pe_1_5_3_N75) );
  AND2_X1 npu_inst_pe_1_5_3_U128 ( .A1(npu_inst_pe_1_5_3_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_5__3__2_), .ZN(
        npu_inst_pe_1_5_3_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_3_U127 ( .A(npu_inst_int_data_res_5__3__3_), .B(
        npu_inst_pe_1_5_3_add_79_carry_3_), .Z(npu_inst_pe_1_5_3_N76) );
  AND2_X1 npu_inst_pe_1_5_3_U126 ( .A1(npu_inst_pe_1_5_3_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_5__3__3_), .ZN(
        npu_inst_pe_1_5_3_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_3_U125 ( .A(npu_inst_int_data_res_5__3__4_), .B(
        npu_inst_pe_1_5_3_add_79_carry_4_), .Z(npu_inst_pe_1_5_3_N77) );
  AND2_X1 npu_inst_pe_1_5_3_U124 ( .A1(npu_inst_pe_1_5_3_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_5__3__4_), .ZN(
        npu_inst_pe_1_5_3_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_3_U123 ( .A(npu_inst_int_data_res_5__3__5_), .B(
        npu_inst_pe_1_5_3_add_79_carry_5_), .Z(npu_inst_pe_1_5_3_N78) );
  AND2_X1 npu_inst_pe_1_5_3_U122 ( .A1(npu_inst_pe_1_5_3_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_5__3__5_), .ZN(
        npu_inst_pe_1_5_3_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_3_U121 ( .A(npu_inst_int_data_res_5__3__6_), .B(
        npu_inst_pe_1_5_3_add_79_carry_6_), .Z(npu_inst_pe_1_5_3_N79) );
  AND2_X1 npu_inst_pe_1_5_3_U120 ( .A1(npu_inst_pe_1_5_3_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_5__3__6_), .ZN(
        npu_inst_pe_1_5_3_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_3_U119 ( .A(npu_inst_int_data_res_5__3__7_), .B(
        npu_inst_pe_1_5_3_add_79_carry_7_), .Z(npu_inst_pe_1_5_3_N80) );
  XNOR2_X1 npu_inst_pe_1_5_3_U118 ( .A(npu_inst_pe_1_5_3_sub_77_carry_2_), .B(
        npu_inst_int_data_res_5__3__2_), .ZN(npu_inst_pe_1_5_3_N67) );
  OR2_X1 npu_inst_pe_1_5_3_U117 ( .A1(npu_inst_int_data_res_5__3__2_), .A2(
        npu_inst_pe_1_5_3_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_5_3_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_3_U116 ( .A(npu_inst_pe_1_5_3_sub_77_carry_3_), .B(
        npu_inst_int_data_res_5__3__3_), .ZN(npu_inst_pe_1_5_3_N68) );
  OR2_X1 npu_inst_pe_1_5_3_U115 ( .A1(npu_inst_int_data_res_5__3__3_), .A2(
        npu_inst_pe_1_5_3_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_5_3_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_3_U114 ( .A(npu_inst_pe_1_5_3_sub_77_carry_4_), .B(
        npu_inst_int_data_res_5__3__4_), .ZN(npu_inst_pe_1_5_3_N69) );
  OR2_X1 npu_inst_pe_1_5_3_U113 ( .A1(npu_inst_int_data_res_5__3__4_), .A2(
        npu_inst_pe_1_5_3_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_5_3_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_3_U112 ( .A(npu_inst_pe_1_5_3_sub_77_carry_5_), .B(
        npu_inst_int_data_res_5__3__5_), .ZN(npu_inst_pe_1_5_3_N70) );
  OR2_X1 npu_inst_pe_1_5_3_U111 ( .A1(npu_inst_int_data_res_5__3__5_), .A2(
        npu_inst_pe_1_5_3_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_5_3_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_3_U110 ( .A(npu_inst_pe_1_5_3_sub_77_carry_6_), .B(
        npu_inst_int_data_res_5__3__6_), .ZN(npu_inst_pe_1_5_3_N71) );
  OR2_X1 npu_inst_pe_1_5_3_U109 ( .A1(npu_inst_int_data_res_5__3__6_), .A2(
        npu_inst_pe_1_5_3_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_5_3_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_3_U108 ( .A(npu_inst_int_data_res_5__3__7_), .B(
        npu_inst_pe_1_5_3_sub_77_carry_7_), .ZN(npu_inst_pe_1_5_3_N72) );
  INV_X1 npu_inst_pe_1_5_3_U107 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_5_3_n6)
         );
  INV_X1 npu_inst_pe_1_5_3_U106 ( .A(npu_inst_pe_1_5_3_n6), .ZN(
        npu_inst_pe_1_5_3_n5) );
  INV_X1 npu_inst_pe_1_5_3_U105 ( .A(npu_inst_n36), .ZN(npu_inst_pe_1_5_3_n2)
         );
  AOI22_X1 npu_inst_pe_1_5_3_U104 ( .A1(npu_inst_int_data_y_6__3__0_), .A2(
        npu_inst_pe_1_5_3_n58), .B1(npu_inst_pe_1_5_3_n118), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_3_n57) );
  INV_X1 npu_inst_pe_1_5_3_U103 ( .A(npu_inst_pe_1_5_3_n57), .ZN(
        npu_inst_pe_1_5_3_n107) );
  AOI22_X1 npu_inst_pe_1_5_3_U102 ( .A1(npu_inst_int_data_y_6__3__0_), .A2(
        npu_inst_pe_1_5_3_n54), .B1(npu_inst_pe_1_5_3_n117), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_3_n53) );
  INV_X1 npu_inst_pe_1_5_3_U99 ( .A(npu_inst_pe_1_5_3_n53), .ZN(
        npu_inst_pe_1_5_3_n108) );
  AOI22_X1 npu_inst_pe_1_5_3_U98 ( .A1(npu_inst_int_data_y_6__3__0_), .A2(
        npu_inst_pe_1_5_3_n50), .B1(npu_inst_pe_1_5_3_n116), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_3_n49) );
  INV_X1 npu_inst_pe_1_5_3_U97 ( .A(npu_inst_pe_1_5_3_n49), .ZN(
        npu_inst_pe_1_5_3_n109) );
  AOI22_X1 npu_inst_pe_1_5_3_U96 ( .A1(npu_inst_int_data_y_6__3__0_), .A2(
        npu_inst_pe_1_5_3_n46), .B1(npu_inst_pe_1_5_3_n115), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_3_n45) );
  INV_X1 npu_inst_pe_1_5_3_U95 ( .A(npu_inst_pe_1_5_3_n45), .ZN(
        npu_inst_pe_1_5_3_n110) );
  AOI22_X1 npu_inst_pe_1_5_3_U94 ( .A1(npu_inst_int_data_y_6__3__0_), .A2(
        npu_inst_pe_1_5_3_n42), .B1(npu_inst_pe_1_5_3_n114), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_3_n41) );
  INV_X1 npu_inst_pe_1_5_3_U93 ( .A(npu_inst_pe_1_5_3_n41), .ZN(
        npu_inst_pe_1_5_3_n111) );
  AOI22_X1 npu_inst_pe_1_5_3_U92 ( .A1(npu_inst_int_data_y_6__3__1_), .A2(
        npu_inst_pe_1_5_3_n58), .B1(npu_inst_pe_1_5_3_n118), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_3_n59) );
  INV_X1 npu_inst_pe_1_5_3_U91 ( .A(npu_inst_pe_1_5_3_n59), .ZN(
        npu_inst_pe_1_5_3_n101) );
  AOI22_X1 npu_inst_pe_1_5_3_U90 ( .A1(npu_inst_int_data_y_6__3__1_), .A2(
        npu_inst_pe_1_5_3_n54), .B1(npu_inst_pe_1_5_3_n117), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_3_n55) );
  INV_X1 npu_inst_pe_1_5_3_U89 ( .A(npu_inst_pe_1_5_3_n55), .ZN(
        npu_inst_pe_1_5_3_n102) );
  AOI22_X1 npu_inst_pe_1_5_3_U88 ( .A1(npu_inst_int_data_y_6__3__1_), .A2(
        npu_inst_pe_1_5_3_n50), .B1(npu_inst_pe_1_5_3_n116), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_3_n51) );
  INV_X1 npu_inst_pe_1_5_3_U87 ( .A(npu_inst_pe_1_5_3_n51), .ZN(
        npu_inst_pe_1_5_3_n103) );
  AOI22_X1 npu_inst_pe_1_5_3_U86 ( .A1(npu_inst_int_data_y_6__3__1_), .A2(
        npu_inst_pe_1_5_3_n46), .B1(npu_inst_pe_1_5_3_n115), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_3_n47) );
  INV_X1 npu_inst_pe_1_5_3_U85 ( .A(npu_inst_pe_1_5_3_n47), .ZN(
        npu_inst_pe_1_5_3_n104) );
  AOI22_X1 npu_inst_pe_1_5_3_U84 ( .A1(npu_inst_int_data_y_6__3__1_), .A2(
        npu_inst_pe_1_5_3_n42), .B1(npu_inst_pe_1_5_3_n114), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_3_n43) );
  INV_X1 npu_inst_pe_1_5_3_U83 ( .A(npu_inst_pe_1_5_3_n43), .ZN(
        npu_inst_pe_1_5_3_n105) );
  AOI22_X1 npu_inst_pe_1_5_3_U82 ( .A1(npu_inst_pe_1_5_3_n38), .A2(
        npu_inst_int_data_y_6__3__1_), .B1(npu_inst_pe_1_5_3_n113), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_3_n39) );
  INV_X1 npu_inst_pe_1_5_3_U81 ( .A(npu_inst_pe_1_5_3_n39), .ZN(
        npu_inst_pe_1_5_3_n106) );
  AND2_X1 npu_inst_pe_1_5_3_U80 ( .A1(npu_inst_pe_1_5_3_N93), .A2(npu_inst_n36), .ZN(npu_inst_int_data_y_5__3__0_) );
  NAND2_X1 npu_inst_pe_1_5_3_U79 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_3_n60), .ZN(npu_inst_pe_1_5_3_n74) );
  OAI21_X1 npu_inst_pe_1_5_3_U78 ( .B1(npu_inst_pe_1_5_3_n63), .B2(
        npu_inst_pe_1_5_3_n60), .A(npu_inst_pe_1_5_3_n74), .ZN(
        npu_inst_pe_1_5_3_n97) );
  NAND2_X1 npu_inst_pe_1_5_3_U77 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_3_n60), .ZN(npu_inst_pe_1_5_3_n73) );
  OAI21_X1 npu_inst_pe_1_5_3_U76 ( .B1(npu_inst_pe_1_5_3_n61), .B2(
        npu_inst_pe_1_5_3_n60), .A(npu_inst_pe_1_5_3_n73), .ZN(
        npu_inst_pe_1_5_3_n96) );
  NAND2_X1 npu_inst_pe_1_5_3_U75 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_3_n56), .ZN(npu_inst_pe_1_5_3_n72) );
  OAI21_X1 npu_inst_pe_1_5_3_U74 ( .B1(npu_inst_pe_1_5_3_n63), .B2(
        npu_inst_pe_1_5_3_n56), .A(npu_inst_pe_1_5_3_n72), .ZN(
        npu_inst_pe_1_5_3_n95) );
  NAND2_X1 npu_inst_pe_1_5_3_U73 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_3_n56), .ZN(npu_inst_pe_1_5_3_n71) );
  OAI21_X1 npu_inst_pe_1_5_3_U72 ( .B1(npu_inst_pe_1_5_3_n61), .B2(
        npu_inst_pe_1_5_3_n56), .A(npu_inst_pe_1_5_3_n71), .ZN(
        npu_inst_pe_1_5_3_n94) );
  NAND2_X1 npu_inst_pe_1_5_3_U71 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_3_n52), .ZN(npu_inst_pe_1_5_3_n70) );
  OAI21_X1 npu_inst_pe_1_5_3_U70 ( .B1(npu_inst_pe_1_5_3_n63), .B2(
        npu_inst_pe_1_5_3_n52), .A(npu_inst_pe_1_5_3_n70), .ZN(
        npu_inst_pe_1_5_3_n93) );
  NAND2_X1 npu_inst_pe_1_5_3_U69 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_3_n52), .ZN(npu_inst_pe_1_5_3_n69) );
  OAI21_X1 npu_inst_pe_1_5_3_U68 ( .B1(npu_inst_pe_1_5_3_n61), .B2(
        npu_inst_pe_1_5_3_n52), .A(npu_inst_pe_1_5_3_n69), .ZN(
        npu_inst_pe_1_5_3_n92) );
  NAND2_X1 npu_inst_pe_1_5_3_U67 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_3_n48), .ZN(npu_inst_pe_1_5_3_n68) );
  OAI21_X1 npu_inst_pe_1_5_3_U66 ( .B1(npu_inst_pe_1_5_3_n63), .B2(
        npu_inst_pe_1_5_3_n48), .A(npu_inst_pe_1_5_3_n68), .ZN(
        npu_inst_pe_1_5_3_n91) );
  NAND2_X1 npu_inst_pe_1_5_3_U65 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_3_n48), .ZN(npu_inst_pe_1_5_3_n67) );
  OAI21_X1 npu_inst_pe_1_5_3_U64 ( .B1(npu_inst_pe_1_5_3_n61), .B2(
        npu_inst_pe_1_5_3_n48), .A(npu_inst_pe_1_5_3_n67), .ZN(
        npu_inst_pe_1_5_3_n90) );
  NAND2_X1 npu_inst_pe_1_5_3_U63 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_3_n44), .ZN(npu_inst_pe_1_5_3_n66) );
  OAI21_X1 npu_inst_pe_1_5_3_U62 ( .B1(npu_inst_pe_1_5_3_n63), .B2(
        npu_inst_pe_1_5_3_n44), .A(npu_inst_pe_1_5_3_n66), .ZN(
        npu_inst_pe_1_5_3_n89) );
  NAND2_X1 npu_inst_pe_1_5_3_U61 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_3_n44), .ZN(npu_inst_pe_1_5_3_n65) );
  OAI21_X1 npu_inst_pe_1_5_3_U60 ( .B1(npu_inst_pe_1_5_3_n61), .B2(
        npu_inst_pe_1_5_3_n44), .A(npu_inst_pe_1_5_3_n65), .ZN(
        npu_inst_pe_1_5_3_n88) );
  NAND2_X1 npu_inst_pe_1_5_3_U59 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_3_n40), .ZN(npu_inst_pe_1_5_3_n64) );
  OAI21_X1 npu_inst_pe_1_5_3_U58 ( .B1(npu_inst_pe_1_5_3_n63), .B2(
        npu_inst_pe_1_5_3_n40), .A(npu_inst_pe_1_5_3_n64), .ZN(
        npu_inst_pe_1_5_3_n87) );
  NAND2_X1 npu_inst_pe_1_5_3_U57 ( .A1(npu_inst_pe_1_5_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_3_n40), .ZN(npu_inst_pe_1_5_3_n62) );
  OAI21_X1 npu_inst_pe_1_5_3_U56 ( .B1(npu_inst_pe_1_5_3_n61), .B2(
        npu_inst_pe_1_5_3_n40), .A(npu_inst_pe_1_5_3_n62), .ZN(
        npu_inst_pe_1_5_3_n86) );
  AOI22_X1 npu_inst_pe_1_5_3_U55 ( .A1(npu_inst_pe_1_5_3_n38), .A2(
        npu_inst_int_data_y_6__3__0_), .B1(npu_inst_pe_1_5_3_n113), .B2(
        npu_inst_pe_1_5_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_3_n37) );
  INV_X1 npu_inst_pe_1_5_3_U54 ( .A(npu_inst_pe_1_5_3_n37), .ZN(
        npu_inst_pe_1_5_3_n112) );
  AND2_X1 npu_inst_pe_1_5_3_U53 ( .A1(npu_inst_n36), .A2(npu_inst_pe_1_5_3_N94), .ZN(npu_inst_int_data_y_5__3__1_) );
  AOI222_X1 npu_inst_pe_1_5_3_U52 ( .A1(npu_inst_int_data_res_6__3__0_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N73), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N65), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n84) );
  INV_X1 npu_inst_pe_1_5_3_U51 ( .A(npu_inst_pe_1_5_3_n84), .ZN(
        npu_inst_pe_1_5_3_n100) );
  AOI222_X1 npu_inst_pe_1_5_3_U50 ( .A1(npu_inst_pe_1_5_3_n1), .A2(
        npu_inst_int_data_res_6__3__7_), .B1(npu_inst_pe_1_5_3_N80), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N72), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n75) );
  INV_X1 npu_inst_pe_1_5_3_U49 ( .A(npu_inst_pe_1_5_3_n75), .ZN(
        npu_inst_pe_1_5_3_n32) );
  AOI222_X1 npu_inst_pe_1_5_3_U48 ( .A1(npu_inst_int_data_res_6__3__1_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N74), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N66), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n83) );
  INV_X1 npu_inst_pe_1_5_3_U47 ( .A(npu_inst_pe_1_5_3_n83), .ZN(
        npu_inst_pe_1_5_3_n99) );
  AOI222_X1 npu_inst_pe_1_5_3_U46 ( .A1(npu_inst_int_data_res_6__3__3_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N76), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N68), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n81) );
  INV_X1 npu_inst_pe_1_5_3_U45 ( .A(npu_inst_pe_1_5_3_n81), .ZN(
        npu_inst_pe_1_5_3_n36) );
  AOI222_X1 npu_inst_pe_1_5_3_U44 ( .A1(npu_inst_int_data_res_6__3__4_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N77), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N69), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n80) );
  INV_X1 npu_inst_pe_1_5_3_U43 ( .A(npu_inst_pe_1_5_3_n80), .ZN(
        npu_inst_pe_1_5_3_n35) );
  AOI222_X1 npu_inst_pe_1_5_3_U42 ( .A1(npu_inst_int_data_res_6__3__5_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N78), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N70), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n79) );
  INV_X1 npu_inst_pe_1_5_3_U41 ( .A(npu_inst_pe_1_5_3_n79), .ZN(
        npu_inst_pe_1_5_3_n34) );
  AOI222_X1 npu_inst_pe_1_5_3_U40 ( .A1(npu_inst_int_data_res_6__3__6_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N79), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N71), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n78) );
  INV_X1 npu_inst_pe_1_5_3_U39 ( .A(npu_inst_pe_1_5_3_n78), .ZN(
        npu_inst_pe_1_5_3_n33) );
  NOR3_X1 npu_inst_pe_1_5_3_U38 ( .A1(npu_inst_pe_1_5_3_n26), .A2(npu_inst_n36), .A3(npu_inst_int_ckg[20]), .ZN(npu_inst_pe_1_5_3_n85) );
  OR2_X1 npu_inst_pe_1_5_3_U37 ( .A1(npu_inst_pe_1_5_3_n85), .A2(
        npu_inst_pe_1_5_3_n1), .ZN(npu_inst_pe_1_5_3_N84) );
  AND2_X1 npu_inst_pe_1_5_3_U36 ( .A1(npu_inst_int_data_x_5__3__1_), .A2(
        npu_inst_pe_1_5_3_int_q_weight_1_), .ZN(npu_inst_pe_1_5_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_3_U35 ( .A1(npu_inst_int_data_x_5__3__0_), .A2(
        npu_inst_pe_1_5_3_int_q_weight_1_), .ZN(npu_inst_pe_1_5_3_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_5_3_U34 ( .A(npu_inst_pe_1_5_3_int_data_1_), .ZN(
        npu_inst_pe_1_5_3_n13) );
  AOI222_X1 npu_inst_pe_1_5_3_U33 ( .A1(npu_inst_int_data_res_6__3__2_), .A2(
        npu_inst_pe_1_5_3_n1), .B1(npu_inst_pe_1_5_3_N75), .B2(
        npu_inst_pe_1_5_3_n76), .C1(npu_inst_pe_1_5_3_N67), .C2(
        npu_inst_pe_1_5_3_n77), .ZN(npu_inst_pe_1_5_3_n82) );
  INV_X1 npu_inst_pe_1_5_3_U32 ( .A(npu_inst_pe_1_5_3_n82), .ZN(
        npu_inst_pe_1_5_3_n98) );
  AOI22_X1 npu_inst_pe_1_5_3_U31 ( .A1(npu_inst_n36), .A2(
        npu_inst_int_data_y_6__3__1_), .B1(npu_inst_pe_1_5_3_n2), .B2(
        npu_inst_int_data_x_5__4__1_), .ZN(npu_inst_pe_1_5_3_n63) );
  AOI22_X1 npu_inst_pe_1_5_3_U30 ( .A1(npu_inst_n36), .A2(
        npu_inst_int_data_y_6__3__0_), .B1(npu_inst_pe_1_5_3_n2), .B2(
        npu_inst_int_data_x_5__4__0_), .ZN(npu_inst_pe_1_5_3_n61) );
  INV_X1 npu_inst_pe_1_5_3_U29 ( .A(npu_inst_pe_1_5_3_int_data_0_), .ZN(
        npu_inst_pe_1_5_3_n12) );
  INV_X1 npu_inst_pe_1_5_3_U28 ( .A(npu_inst_n50), .ZN(npu_inst_pe_1_5_3_n4)
         );
  OR3_X1 npu_inst_pe_1_5_3_U27 ( .A1(npu_inst_pe_1_5_3_n5), .A2(
        npu_inst_pe_1_5_3_n7), .A3(npu_inst_pe_1_5_3_n4), .ZN(
        npu_inst_pe_1_5_3_n56) );
  OR3_X1 npu_inst_pe_1_5_3_U26 ( .A1(npu_inst_pe_1_5_3_n4), .A2(
        npu_inst_pe_1_5_3_n7), .A3(npu_inst_pe_1_5_3_n6), .ZN(
        npu_inst_pe_1_5_3_n48) );
  INV_X1 npu_inst_pe_1_5_3_U25 ( .A(npu_inst_pe_1_5_3_n4), .ZN(
        npu_inst_pe_1_5_3_n3) );
  OR3_X1 npu_inst_pe_1_5_3_U24 ( .A1(npu_inst_pe_1_5_3_n3), .A2(
        npu_inst_pe_1_5_3_n7), .A3(npu_inst_pe_1_5_3_n6), .ZN(
        npu_inst_pe_1_5_3_n52) );
  OR3_X1 npu_inst_pe_1_5_3_U23 ( .A1(npu_inst_pe_1_5_3_n5), .A2(
        npu_inst_pe_1_5_3_n7), .A3(npu_inst_pe_1_5_3_n3), .ZN(
        npu_inst_pe_1_5_3_n60) );
  BUF_X1 npu_inst_pe_1_5_3_U22 ( .A(npu_inst_n17), .Z(npu_inst_pe_1_5_3_n1) );
  NOR2_X1 npu_inst_pe_1_5_3_U21 ( .A1(npu_inst_pe_1_5_3_n60), .A2(
        npu_inst_pe_1_5_3_n2), .ZN(npu_inst_pe_1_5_3_n58) );
  NOR2_X1 npu_inst_pe_1_5_3_U20 ( .A1(npu_inst_pe_1_5_3_n56), .A2(
        npu_inst_pe_1_5_3_n2), .ZN(npu_inst_pe_1_5_3_n54) );
  NOR2_X1 npu_inst_pe_1_5_3_U19 ( .A1(npu_inst_pe_1_5_3_n52), .A2(
        npu_inst_pe_1_5_3_n2), .ZN(npu_inst_pe_1_5_3_n50) );
  NOR2_X1 npu_inst_pe_1_5_3_U18 ( .A1(npu_inst_pe_1_5_3_n48), .A2(
        npu_inst_pe_1_5_3_n2), .ZN(npu_inst_pe_1_5_3_n46) );
  NOR2_X1 npu_inst_pe_1_5_3_U17 ( .A1(npu_inst_pe_1_5_3_n40), .A2(
        npu_inst_pe_1_5_3_n2), .ZN(npu_inst_pe_1_5_3_n38) );
  NOR2_X1 npu_inst_pe_1_5_3_U16 ( .A1(npu_inst_pe_1_5_3_n44), .A2(
        npu_inst_pe_1_5_3_n2), .ZN(npu_inst_pe_1_5_3_n42) );
  BUF_X1 npu_inst_pe_1_5_3_U15 ( .A(npu_inst_n79), .Z(npu_inst_pe_1_5_3_n7) );
  INV_X1 npu_inst_pe_1_5_3_U14 ( .A(npu_inst_n105), .ZN(npu_inst_pe_1_5_3_n11)
         );
  INV_X1 npu_inst_pe_1_5_3_U13 ( .A(npu_inst_pe_1_5_3_n38), .ZN(
        npu_inst_pe_1_5_3_n113) );
  INV_X1 npu_inst_pe_1_5_3_U12 ( .A(npu_inst_pe_1_5_3_n58), .ZN(
        npu_inst_pe_1_5_3_n118) );
  INV_X1 npu_inst_pe_1_5_3_U11 ( .A(npu_inst_pe_1_5_3_n54), .ZN(
        npu_inst_pe_1_5_3_n117) );
  INV_X1 npu_inst_pe_1_5_3_U10 ( .A(npu_inst_pe_1_5_3_n50), .ZN(
        npu_inst_pe_1_5_3_n116) );
  INV_X1 npu_inst_pe_1_5_3_U9 ( .A(npu_inst_pe_1_5_3_n46), .ZN(
        npu_inst_pe_1_5_3_n115) );
  INV_X1 npu_inst_pe_1_5_3_U8 ( .A(npu_inst_pe_1_5_3_n42), .ZN(
        npu_inst_pe_1_5_3_n114) );
  BUF_X1 npu_inst_pe_1_5_3_U7 ( .A(npu_inst_pe_1_5_3_n11), .Z(
        npu_inst_pe_1_5_3_n10) );
  BUF_X1 npu_inst_pe_1_5_3_U6 ( .A(npu_inst_pe_1_5_3_n11), .Z(
        npu_inst_pe_1_5_3_n9) );
  BUF_X1 npu_inst_pe_1_5_3_U5 ( .A(npu_inst_pe_1_5_3_n11), .Z(
        npu_inst_pe_1_5_3_n8) );
  NOR2_X1 npu_inst_pe_1_5_3_U4 ( .A1(npu_inst_pe_1_5_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_3_n1), .ZN(npu_inst_pe_1_5_3_n76) );
  NOR2_X1 npu_inst_pe_1_5_3_U3 ( .A1(npu_inst_pe_1_5_3_n27), .A2(
        npu_inst_pe_1_5_3_n1), .ZN(npu_inst_pe_1_5_3_n77) );
  FA_X1 npu_inst_pe_1_5_3_sub_77_U2_1 ( .A(npu_inst_int_data_res_5__3__1_), 
        .B(npu_inst_pe_1_5_3_n13), .CI(npu_inst_pe_1_5_3_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_5_3_sub_77_carry_2_), .S(npu_inst_pe_1_5_3_N66) );
  FA_X1 npu_inst_pe_1_5_3_add_79_U1_1 ( .A(npu_inst_int_data_res_5__3__1_), 
        .B(npu_inst_pe_1_5_3_int_data_1_), .CI(
        npu_inst_pe_1_5_3_add_79_carry_1_), .CO(
        npu_inst_pe_1_5_3_add_79_carry_2_), .S(npu_inst_pe_1_5_3_N74) );
  NAND3_X1 npu_inst_pe_1_5_3_U101 ( .A1(npu_inst_pe_1_5_3_n4), .A2(
        npu_inst_pe_1_5_3_n6), .A3(npu_inst_pe_1_5_3_n7), .ZN(
        npu_inst_pe_1_5_3_n44) );
  NAND3_X1 npu_inst_pe_1_5_3_U100 ( .A1(npu_inst_pe_1_5_3_n3), .A2(
        npu_inst_pe_1_5_3_n6), .A3(npu_inst_pe_1_5_3_n7), .ZN(
        npu_inst_pe_1_5_3_n40) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_3_n33), .CK(
        npu_inst_pe_1_5_3_net3489), .RN(npu_inst_pe_1_5_3_n8), .Q(
        npu_inst_int_data_res_5__3__6_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_3_n34), .CK(
        npu_inst_pe_1_5_3_net3489), .RN(npu_inst_pe_1_5_3_n8), .Q(
        npu_inst_int_data_res_5__3__5_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_3_n35), .CK(
        npu_inst_pe_1_5_3_net3489), .RN(npu_inst_pe_1_5_3_n8), .Q(
        npu_inst_int_data_res_5__3__4_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_3_n36), .CK(
        npu_inst_pe_1_5_3_net3489), .RN(npu_inst_pe_1_5_3_n8), .Q(
        npu_inst_int_data_res_5__3__3_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_3_n98), .CK(
        npu_inst_pe_1_5_3_net3489), .RN(npu_inst_pe_1_5_3_n8), .Q(
        npu_inst_int_data_res_5__3__2_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_3_n99), .CK(
        npu_inst_pe_1_5_3_net3489), .RN(npu_inst_pe_1_5_3_n8), .Q(
        npu_inst_int_data_res_5__3__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_3_n32), .CK(
        npu_inst_pe_1_5_3_net3489), .RN(npu_inst_pe_1_5_3_n8), .Q(
        npu_inst_int_data_res_5__3__7_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_3_n100), 
        .CK(npu_inst_pe_1_5_3_net3489), .RN(npu_inst_pe_1_5_3_n8), .Q(
        npu_inst_int_data_res_5__3__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_weight_reg_0_ ( .D(npu_inst_n91), .CK(
        npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n8), .Q(
        npu_inst_pe_1_5_3_int_q_weight_0_), .QN(npu_inst_pe_1_5_3_n27) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_weight_reg_1_ ( .D(npu_inst_n97), .CK(
        npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n8), .Q(
        npu_inst_pe_1_5_3_int_q_weight_1_), .QN(npu_inst_pe_1_5_3_n26) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_3_n112), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n8), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_3_n106), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n8), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_3_n111), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_3_n105), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_3_n110), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_3_n104), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_3_n109), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_3_n103), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_3_n108), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_3_n102), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_3_n107), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_3_n101), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_3_n86), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_3_n87), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n9), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_3_n88), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_3_n89), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_3_n90), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_3_n91), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_3_n92), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_3_n93), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_3_n94), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_3_n95), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_3_n96), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_3_n97), 
        .CK(npu_inst_pe_1_5_3_net3495), .RN(npu_inst_pe_1_5_3_n10), .Q(
        npu_inst_pe_1_5_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_3_net3489) );
  CLKGATETST_X1 npu_inst_pe_1_5_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n44), .SE(1'b0), .GCK(npu_inst_pe_1_5_3_net3495) );
  MUX2_X1 npu_inst_pe_1_5_4_U153 ( .A(npu_inst_pe_1_5_4_n31), .B(
        npu_inst_pe_1_5_4_n28), .S(npu_inst_pe_1_5_4_n7), .Z(
        npu_inst_pe_1_5_4_N93) );
  MUX2_X1 npu_inst_pe_1_5_4_U152 ( .A(npu_inst_pe_1_5_4_n30), .B(
        npu_inst_pe_1_5_4_n29), .S(npu_inst_pe_1_5_4_n5), .Z(
        npu_inst_pe_1_5_4_n31) );
  MUX2_X1 npu_inst_pe_1_5_4_U151 ( .A(npu_inst_pe_1_5_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_4_n3), .Z(
        npu_inst_pe_1_5_4_n30) );
  MUX2_X1 npu_inst_pe_1_5_4_U150 ( .A(npu_inst_pe_1_5_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_4_n3), .Z(
        npu_inst_pe_1_5_4_n29) );
  MUX2_X1 npu_inst_pe_1_5_4_U149 ( .A(npu_inst_pe_1_5_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_4_n3), .Z(
        npu_inst_pe_1_5_4_n28) );
  MUX2_X1 npu_inst_pe_1_5_4_U148 ( .A(npu_inst_pe_1_5_4_n25), .B(
        npu_inst_pe_1_5_4_n22), .S(npu_inst_pe_1_5_4_n7), .Z(
        npu_inst_pe_1_5_4_N94) );
  MUX2_X1 npu_inst_pe_1_5_4_U147 ( .A(npu_inst_pe_1_5_4_n24), .B(
        npu_inst_pe_1_5_4_n23), .S(npu_inst_pe_1_5_4_n5), .Z(
        npu_inst_pe_1_5_4_n25) );
  MUX2_X1 npu_inst_pe_1_5_4_U146 ( .A(npu_inst_pe_1_5_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_4_n3), .Z(
        npu_inst_pe_1_5_4_n24) );
  MUX2_X1 npu_inst_pe_1_5_4_U145 ( .A(npu_inst_pe_1_5_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_4_n3), .Z(
        npu_inst_pe_1_5_4_n23) );
  MUX2_X1 npu_inst_pe_1_5_4_U144 ( .A(npu_inst_pe_1_5_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_4_n3), .Z(
        npu_inst_pe_1_5_4_n22) );
  MUX2_X1 npu_inst_pe_1_5_4_U143 ( .A(npu_inst_pe_1_5_4_n21), .B(
        npu_inst_pe_1_5_4_n18), .S(npu_inst_pe_1_5_4_n7), .Z(
        npu_inst_int_data_x_5__4__1_) );
  MUX2_X1 npu_inst_pe_1_5_4_U142 ( .A(npu_inst_pe_1_5_4_n20), .B(
        npu_inst_pe_1_5_4_n19), .S(npu_inst_pe_1_5_4_n5), .Z(
        npu_inst_pe_1_5_4_n21) );
  MUX2_X1 npu_inst_pe_1_5_4_U141 ( .A(npu_inst_pe_1_5_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_4_n3), .Z(
        npu_inst_pe_1_5_4_n20) );
  MUX2_X1 npu_inst_pe_1_5_4_U140 ( .A(npu_inst_pe_1_5_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_4_n3), .Z(
        npu_inst_pe_1_5_4_n19) );
  MUX2_X1 npu_inst_pe_1_5_4_U139 ( .A(npu_inst_pe_1_5_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_4_n3), .Z(
        npu_inst_pe_1_5_4_n18) );
  MUX2_X1 npu_inst_pe_1_5_4_U138 ( .A(npu_inst_pe_1_5_4_n17), .B(
        npu_inst_pe_1_5_4_n14), .S(npu_inst_pe_1_5_4_n7), .Z(
        npu_inst_int_data_x_5__4__0_) );
  MUX2_X1 npu_inst_pe_1_5_4_U137 ( .A(npu_inst_pe_1_5_4_n16), .B(
        npu_inst_pe_1_5_4_n15), .S(npu_inst_pe_1_5_4_n5), .Z(
        npu_inst_pe_1_5_4_n17) );
  MUX2_X1 npu_inst_pe_1_5_4_U136 ( .A(npu_inst_pe_1_5_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_4_n3), .Z(
        npu_inst_pe_1_5_4_n16) );
  MUX2_X1 npu_inst_pe_1_5_4_U135 ( .A(npu_inst_pe_1_5_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_4_n3), .Z(
        npu_inst_pe_1_5_4_n15) );
  MUX2_X1 npu_inst_pe_1_5_4_U134 ( .A(npu_inst_pe_1_5_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_4_n3), .Z(
        npu_inst_pe_1_5_4_n14) );
  XOR2_X1 npu_inst_pe_1_5_4_U133 ( .A(npu_inst_pe_1_5_4_int_data_0_), .B(
        npu_inst_int_data_res_5__4__0_), .Z(npu_inst_pe_1_5_4_N73) );
  AND2_X1 npu_inst_pe_1_5_4_U132 ( .A1(npu_inst_int_data_res_5__4__0_), .A2(
        npu_inst_pe_1_5_4_int_data_0_), .ZN(npu_inst_pe_1_5_4_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_4_U131 ( .A(npu_inst_int_data_res_5__4__0_), .B(
        npu_inst_pe_1_5_4_n12), .ZN(npu_inst_pe_1_5_4_N65) );
  OR2_X1 npu_inst_pe_1_5_4_U130 ( .A1(npu_inst_pe_1_5_4_n12), .A2(
        npu_inst_int_data_res_5__4__0_), .ZN(npu_inst_pe_1_5_4_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_4_U129 ( .A(npu_inst_int_data_res_5__4__2_), .B(
        npu_inst_pe_1_5_4_add_79_carry_2_), .Z(npu_inst_pe_1_5_4_N75) );
  AND2_X1 npu_inst_pe_1_5_4_U128 ( .A1(npu_inst_pe_1_5_4_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_5__4__2_), .ZN(
        npu_inst_pe_1_5_4_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_4_U127 ( .A(npu_inst_int_data_res_5__4__3_), .B(
        npu_inst_pe_1_5_4_add_79_carry_3_), .Z(npu_inst_pe_1_5_4_N76) );
  AND2_X1 npu_inst_pe_1_5_4_U126 ( .A1(npu_inst_pe_1_5_4_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_5__4__3_), .ZN(
        npu_inst_pe_1_5_4_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_4_U125 ( .A(npu_inst_int_data_res_5__4__4_), .B(
        npu_inst_pe_1_5_4_add_79_carry_4_), .Z(npu_inst_pe_1_5_4_N77) );
  AND2_X1 npu_inst_pe_1_5_4_U124 ( .A1(npu_inst_pe_1_5_4_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_5__4__4_), .ZN(
        npu_inst_pe_1_5_4_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_4_U123 ( .A(npu_inst_int_data_res_5__4__5_), .B(
        npu_inst_pe_1_5_4_add_79_carry_5_), .Z(npu_inst_pe_1_5_4_N78) );
  AND2_X1 npu_inst_pe_1_5_4_U122 ( .A1(npu_inst_pe_1_5_4_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_5__4__5_), .ZN(
        npu_inst_pe_1_5_4_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_4_U121 ( .A(npu_inst_int_data_res_5__4__6_), .B(
        npu_inst_pe_1_5_4_add_79_carry_6_), .Z(npu_inst_pe_1_5_4_N79) );
  AND2_X1 npu_inst_pe_1_5_4_U120 ( .A1(npu_inst_pe_1_5_4_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_5__4__6_), .ZN(
        npu_inst_pe_1_5_4_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_4_U119 ( .A(npu_inst_int_data_res_5__4__7_), .B(
        npu_inst_pe_1_5_4_add_79_carry_7_), .Z(npu_inst_pe_1_5_4_N80) );
  XNOR2_X1 npu_inst_pe_1_5_4_U118 ( .A(npu_inst_pe_1_5_4_sub_77_carry_2_), .B(
        npu_inst_int_data_res_5__4__2_), .ZN(npu_inst_pe_1_5_4_N67) );
  OR2_X1 npu_inst_pe_1_5_4_U117 ( .A1(npu_inst_int_data_res_5__4__2_), .A2(
        npu_inst_pe_1_5_4_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_5_4_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_4_U116 ( .A(npu_inst_pe_1_5_4_sub_77_carry_3_), .B(
        npu_inst_int_data_res_5__4__3_), .ZN(npu_inst_pe_1_5_4_N68) );
  OR2_X1 npu_inst_pe_1_5_4_U115 ( .A1(npu_inst_int_data_res_5__4__3_), .A2(
        npu_inst_pe_1_5_4_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_5_4_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_4_U114 ( .A(npu_inst_pe_1_5_4_sub_77_carry_4_), .B(
        npu_inst_int_data_res_5__4__4_), .ZN(npu_inst_pe_1_5_4_N69) );
  OR2_X1 npu_inst_pe_1_5_4_U113 ( .A1(npu_inst_int_data_res_5__4__4_), .A2(
        npu_inst_pe_1_5_4_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_5_4_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_4_U112 ( .A(npu_inst_pe_1_5_4_sub_77_carry_5_), .B(
        npu_inst_int_data_res_5__4__5_), .ZN(npu_inst_pe_1_5_4_N70) );
  OR2_X1 npu_inst_pe_1_5_4_U111 ( .A1(npu_inst_int_data_res_5__4__5_), .A2(
        npu_inst_pe_1_5_4_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_5_4_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_4_U110 ( .A(npu_inst_pe_1_5_4_sub_77_carry_6_), .B(
        npu_inst_int_data_res_5__4__6_), .ZN(npu_inst_pe_1_5_4_N71) );
  OR2_X1 npu_inst_pe_1_5_4_U109 ( .A1(npu_inst_int_data_res_5__4__6_), .A2(
        npu_inst_pe_1_5_4_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_5_4_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_4_U108 ( .A(npu_inst_int_data_res_5__4__7_), .B(
        npu_inst_pe_1_5_4_sub_77_carry_7_), .ZN(npu_inst_pe_1_5_4_N72) );
  INV_X1 npu_inst_pe_1_5_4_U107 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_5_4_n6)
         );
  INV_X1 npu_inst_pe_1_5_4_U106 ( .A(npu_inst_pe_1_5_4_n6), .ZN(
        npu_inst_pe_1_5_4_n5) );
  INV_X1 npu_inst_pe_1_5_4_U105 ( .A(npu_inst_n36), .ZN(npu_inst_pe_1_5_4_n2)
         );
  AOI22_X1 npu_inst_pe_1_5_4_U104 ( .A1(npu_inst_int_data_y_6__4__0_), .A2(
        npu_inst_pe_1_5_4_n58), .B1(npu_inst_pe_1_5_4_n118), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_4_n57) );
  INV_X1 npu_inst_pe_1_5_4_U103 ( .A(npu_inst_pe_1_5_4_n57), .ZN(
        npu_inst_pe_1_5_4_n107) );
  AOI22_X1 npu_inst_pe_1_5_4_U102 ( .A1(npu_inst_int_data_y_6__4__0_), .A2(
        npu_inst_pe_1_5_4_n54), .B1(npu_inst_pe_1_5_4_n117), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_4_n53) );
  INV_X1 npu_inst_pe_1_5_4_U99 ( .A(npu_inst_pe_1_5_4_n53), .ZN(
        npu_inst_pe_1_5_4_n108) );
  AOI22_X1 npu_inst_pe_1_5_4_U98 ( .A1(npu_inst_int_data_y_6__4__0_), .A2(
        npu_inst_pe_1_5_4_n50), .B1(npu_inst_pe_1_5_4_n116), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_4_n49) );
  INV_X1 npu_inst_pe_1_5_4_U97 ( .A(npu_inst_pe_1_5_4_n49), .ZN(
        npu_inst_pe_1_5_4_n109) );
  AOI22_X1 npu_inst_pe_1_5_4_U96 ( .A1(npu_inst_int_data_y_6__4__0_), .A2(
        npu_inst_pe_1_5_4_n46), .B1(npu_inst_pe_1_5_4_n115), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_4_n45) );
  INV_X1 npu_inst_pe_1_5_4_U95 ( .A(npu_inst_pe_1_5_4_n45), .ZN(
        npu_inst_pe_1_5_4_n110) );
  AOI22_X1 npu_inst_pe_1_5_4_U94 ( .A1(npu_inst_int_data_y_6__4__0_), .A2(
        npu_inst_pe_1_5_4_n42), .B1(npu_inst_pe_1_5_4_n114), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_4_n41) );
  INV_X1 npu_inst_pe_1_5_4_U93 ( .A(npu_inst_pe_1_5_4_n41), .ZN(
        npu_inst_pe_1_5_4_n111) );
  AOI22_X1 npu_inst_pe_1_5_4_U92 ( .A1(npu_inst_int_data_y_6__4__1_), .A2(
        npu_inst_pe_1_5_4_n58), .B1(npu_inst_pe_1_5_4_n118), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_4_n59) );
  INV_X1 npu_inst_pe_1_5_4_U91 ( .A(npu_inst_pe_1_5_4_n59), .ZN(
        npu_inst_pe_1_5_4_n101) );
  AOI22_X1 npu_inst_pe_1_5_4_U90 ( .A1(npu_inst_int_data_y_6__4__1_), .A2(
        npu_inst_pe_1_5_4_n54), .B1(npu_inst_pe_1_5_4_n117), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_4_n55) );
  INV_X1 npu_inst_pe_1_5_4_U89 ( .A(npu_inst_pe_1_5_4_n55), .ZN(
        npu_inst_pe_1_5_4_n102) );
  AOI22_X1 npu_inst_pe_1_5_4_U88 ( .A1(npu_inst_int_data_y_6__4__1_), .A2(
        npu_inst_pe_1_5_4_n50), .B1(npu_inst_pe_1_5_4_n116), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_4_n51) );
  INV_X1 npu_inst_pe_1_5_4_U87 ( .A(npu_inst_pe_1_5_4_n51), .ZN(
        npu_inst_pe_1_5_4_n103) );
  AOI22_X1 npu_inst_pe_1_5_4_U86 ( .A1(npu_inst_int_data_y_6__4__1_), .A2(
        npu_inst_pe_1_5_4_n46), .B1(npu_inst_pe_1_5_4_n115), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_4_n47) );
  INV_X1 npu_inst_pe_1_5_4_U85 ( .A(npu_inst_pe_1_5_4_n47), .ZN(
        npu_inst_pe_1_5_4_n104) );
  AOI22_X1 npu_inst_pe_1_5_4_U84 ( .A1(npu_inst_int_data_y_6__4__1_), .A2(
        npu_inst_pe_1_5_4_n42), .B1(npu_inst_pe_1_5_4_n114), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_4_n43) );
  INV_X1 npu_inst_pe_1_5_4_U83 ( .A(npu_inst_pe_1_5_4_n43), .ZN(
        npu_inst_pe_1_5_4_n105) );
  AOI22_X1 npu_inst_pe_1_5_4_U82 ( .A1(npu_inst_pe_1_5_4_n38), .A2(
        npu_inst_int_data_y_6__4__1_), .B1(npu_inst_pe_1_5_4_n113), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_4_n39) );
  INV_X1 npu_inst_pe_1_5_4_U81 ( .A(npu_inst_pe_1_5_4_n39), .ZN(
        npu_inst_pe_1_5_4_n106) );
  AND2_X1 npu_inst_pe_1_5_4_U80 ( .A1(npu_inst_pe_1_5_4_N93), .A2(npu_inst_n36), .ZN(npu_inst_int_data_y_5__4__0_) );
  NAND2_X1 npu_inst_pe_1_5_4_U79 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_4_n60), .ZN(npu_inst_pe_1_5_4_n74) );
  OAI21_X1 npu_inst_pe_1_5_4_U78 ( .B1(npu_inst_pe_1_5_4_n63), .B2(
        npu_inst_pe_1_5_4_n60), .A(npu_inst_pe_1_5_4_n74), .ZN(
        npu_inst_pe_1_5_4_n97) );
  NAND2_X1 npu_inst_pe_1_5_4_U77 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_4_n60), .ZN(npu_inst_pe_1_5_4_n73) );
  OAI21_X1 npu_inst_pe_1_5_4_U76 ( .B1(npu_inst_pe_1_5_4_n61), .B2(
        npu_inst_pe_1_5_4_n60), .A(npu_inst_pe_1_5_4_n73), .ZN(
        npu_inst_pe_1_5_4_n96) );
  NAND2_X1 npu_inst_pe_1_5_4_U75 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_4_n56), .ZN(npu_inst_pe_1_5_4_n72) );
  OAI21_X1 npu_inst_pe_1_5_4_U74 ( .B1(npu_inst_pe_1_5_4_n63), .B2(
        npu_inst_pe_1_5_4_n56), .A(npu_inst_pe_1_5_4_n72), .ZN(
        npu_inst_pe_1_5_4_n95) );
  NAND2_X1 npu_inst_pe_1_5_4_U73 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_4_n56), .ZN(npu_inst_pe_1_5_4_n71) );
  OAI21_X1 npu_inst_pe_1_5_4_U72 ( .B1(npu_inst_pe_1_5_4_n61), .B2(
        npu_inst_pe_1_5_4_n56), .A(npu_inst_pe_1_5_4_n71), .ZN(
        npu_inst_pe_1_5_4_n94) );
  NAND2_X1 npu_inst_pe_1_5_4_U71 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_4_n52), .ZN(npu_inst_pe_1_5_4_n70) );
  OAI21_X1 npu_inst_pe_1_5_4_U70 ( .B1(npu_inst_pe_1_5_4_n63), .B2(
        npu_inst_pe_1_5_4_n52), .A(npu_inst_pe_1_5_4_n70), .ZN(
        npu_inst_pe_1_5_4_n93) );
  NAND2_X1 npu_inst_pe_1_5_4_U69 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_4_n52), .ZN(npu_inst_pe_1_5_4_n69) );
  OAI21_X1 npu_inst_pe_1_5_4_U68 ( .B1(npu_inst_pe_1_5_4_n61), .B2(
        npu_inst_pe_1_5_4_n52), .A(npu_inst_pe_1_5_4_n69), .ZN(
        npu_inst_pe_1_5_4_n92) );
  NAND2_X1 npu_inst_pe_1_5_4_U67 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_4_n48), .ZN(npu_inst_pe_1_5_4_n68) );
  OAI21_X1 npu_inst_pe_1_5_4_U66 ( .B1(npu_inst_pe_1_5_4_n63), .B2(
        npu_inst_pe_1_5_4_n48), .A(npu_inst_pe_1_5_4_n68), .ZN(
        npu_inst_pe_1_5_4_n91) );
  NAND2_X1 npu_inst_pe_1_5_4_U65 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_4_n48), .ZN(npu_inst_pe_1_5_4_n67) );
  OAI21_X1 npu_inst_pe_1_5_4_U64 ( .B1(npu_inst_pe_1_5_4_n61), .B2(
        npu_inst_pe_1_5_4_n48), .A(npu_inst_pe_1_5_4_n67), .ZN(
        npu_inst_pe_1_5_4_n90) );
  NAND2_X1 npu_inst_pe_1_5_4_U63 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_4_n44), .ZN(npu_inst_pe_1_5_4_n66) );
  OAI21_X1 npu_inst_pe_1_5_4_U62 ( .B1(npu_inst_pe_1_5_4_n63), .B2(
        npu_inst_pe_1_5_4_n44), .A(npu_inst_pe_1_5_4_n66), .ZN(
        npu_inst_pe_1_5_4_n89) );
  NAND2_X1 npu_inst_pe_1_5_4_U61 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_4_n44), .ZN(npu_inst_pe_1_5_4_n65) );
  OAI21_X1 npu_inst_pe_1_5_4_U60 ( .B1(npu_inst_pe_1_5_4_n61), .B2(
        npu_inst_pe_1_5_4_n44), .A(npu_inst_pe_1_5_4_n65), .ZN(
        npu_inst_pe_1_5_4_n88) );
  NAND2_X1 npu_inst_pe_1_5_4_U59 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_4_n40), .ZN(npu_inst_pe_1_5_4_n64) );
  OAI21_X1 npu_inst_pe_1_5_4_U58 ( .B1(npu_inst_pe_1_5_4_n63), .B2(
        npu_inst_pe_1_5_4_n40), .A(npu_inst_pe_1_5_4_n64), .ZN(
        npu_inst_pe_1_5_4_n87) );
  NAND2_X1 npu_inst_pe_1_5_4_U57 ( .A1(npu_inst_pe_1_5_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_4_n40), .ZN(npu_inst_pe_1_5_4_n62) );
  OAI21_X1 npu_inst_pe_1_5_4_U56 ( .B1(npu_inst_pe_1_5_4_n61), .B2(
        npu_inst_pe_1_5_4_n40), .A(npu_inst_pe_1_5_4_n62), .ZN(
        npu_inst_pe_1_5_4_n86) );
  AOI22_X1 npu_inst_pe_1_5_4_U55 ( .A1(npu_inst_pe_1_5_4_n38), .A2(
        npu_inst_int_data_y_6__4__0_), .B1(npu_inst_pe_1_5_4_n113), .B2(
        npu_inst_pe_1_5_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_4_n37) );
  INV_X1 npu_inst_pe_1_5_4_U54 ( .A(npu_inst_pe_1_5_4_n37), .ZN(
        npu_inst_pe_1_5_4_n112) );
  AND2_X1 npu_inst_pe_1_5_4_U53 ( .A1(npu_inst_n36), .A2(npu_inst_pe_1_5_4_N94), .ZN(npu_inst_int_data_y_5__4__1_) );
  AOI222_X1 npu_inst_pe_1_5_4_U52 ( .A1(npu_inst_int_data_res_6__4__0_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N73), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N65), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n84) );
  INV_X1 npu_inst_pe_1_5_4_U51 ( .A(npu_inst_pe_1_5_4_n84), .ZN(
        npu_inst_pe_1_5_4_n100) );
  AOI222_X1 npu_inst_pe_1_5_4_U50 ( .A1(npu_inst_pe_1_5_4_n1), .A2(
        npu_inst_int_data_res_6__4__7_), .B1(npu_inst_pe_1_5_4_N80), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N72), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n75) );
  INV_X1 npu_inst_pe_1_5_4_U49 ( .A(npu_inst_pe_1_5_4_n75), .ZN(
        npu_inst_pe_1_5_4_n32) );
  AOI222_X1 npu_inst_pe_1_5_4_U48 ( .A1(npu_inst_int_data_res_6__4__1_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N74), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N66), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n83) );
  INV_X1 npu_inst_pe_1_5_4_U47 ( .A(npu_inst_pe_1_5_4_n83), .ZN(
        npu_inst_pe_1_5_4_n99) );
  AOI222_X1 npu_inst_pe_1_5_4_U46 ( .A1(npu_inst_int_data_res_6__4__3_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N76), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N68), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n81) );
  INV_X1 npu_inst_pe_1_5_4_U45 ( .A(npu_inst_pe_1_5_4_n81), .ZN(
        npu_inst_pe_1_5_4_n36) );
  AOI222_X1 npu_inst_pe_1_5_4_U44 ( .A1(npu_inst_int_data_res_6__4__4_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N77), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N69), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n80) );
  INV_X1 npu_inst_pe_1_5_4_U43 ( .A(npu_inst_pe_1_5_4_n80), .ZN(
        npu_inst_pe_1_5_4_n35) );
  AOI222_X1 npu_inst_pe_1_5_4_U42 ( .A1(npu_inst_int_data_res_6__4__5_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N78), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N70), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n79) );
  INV_X1 npu_inst_pe_1_5_4_U41 ( .A(npu_inst_pe_1_5_4_n79), .ZN(
        npu_inst_pe_1_5_4_n34) );
  AOI222_X1 npu_inst_pe_1_5_4_U40 ( .A1(npu_inst_int_data_res_6__4__6_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N79), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N71), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n78) );
  INV_X1 npu_inst_pe_1_5_4_U39 ( .A(npu_inst_pe_1_5_4_n78), .ZN(
        npu_inst_pe_1_5_4_n33) );
  NOR3_X1 npu_inst_pe_1_5_4_U38 ( .A1(npu_inst_pe_1_5_4_n26), .A2(npu_inst_n36), .A3(npu_inst_int_ckg[19]), .ZN(npu_inst_pe_1_5_4_n85) );
  OR2_X1 npu_inst_pe_1_5_4_U37 ( .A1(npu_inst_pe_1_5_4_n85), .A2(
        npu_inst_pe_1_5_4_n1), .ZN(npu_inst_pe_1_5_4_N84) );
  AND2_X1 npu_inst_pe_1_5_4_U36 ( .A1(npu_inst_int_data_x_5__4__1_), .A2(
        npu_inst_pe_1_5_4_int_q_weight_1_), .ZN(npu_inst_pe_1_5_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_4_U35 ( .A1(npu_inst_int_data_x_5__4__0_), .A2(
        npu_inst_pe_1_5_4_int_q_weight_1_), .ZN(npu_inst_pe_1_5_4_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_5_4_U34 ( .A(npu_inst_pe_1_5_4_int_data_1_), .ZN(
        npu_inst_pe_1_5_4_n13) );
  AOI222_X1 npu_inst_pe_1_5_4_U33 ( .A1(npu_inst_int_data_res_6__4__2_), .A2(
        npu_inst_pe_1_5_4_n1), .B1(npu_inst_pe_1_5_4_N75), .B2(
        npu_inst_pe_1_5_4_n76), .C1(npu_inst_pe_1_5_4_N67), .C2(
        npu_inst_pe_1_5_4_n77), .ZN(npu_inst_pe_1_5_4_n82) );
  INV_X1 npu_inst_pe_1_5_4_U32 ( .A(npu_inst_pe_1_5_4_n82), .ZN(
        npu_inst_pe_1_5_4_n98) );
  AOI22_X1 npu_inst_pe_1_5_4_U31 ( .A1(npu_inst_n36), .A2(
        npu_inst_int_data_y_6__4__1_), .B1(npu_inst_pe_1_5_4_n2), .B2(
        npu_inst_int_data_x_5__5__1_), .ZN(npu_inst_pe_1_5_4_n63) );
  AOI22_X1 npu_inst_pe_1_5_4_U30 ( .A1(npu_inst_n36), .A2(
        npu_inst_int_data_y_6__4__0_), .B1(npu_inst_pe_1_5_4_n2), .B2(
        npu_inst_int_data_x_5__5__0_), .ZN(npu_inst_pe_1_5_4_n61) );
  INV_X1 npu_inst_pe_1_5_4_U29 ( .A(npu_inst_pe_1_5_4_int_data_0_), .ZN(
        npu_inst_pe_1_5_4_n12) );
  INV_X1 npu_inst_pe_1_5_4_U28 ( .A(npu_inst_n50), .ZN(npu_inst_pe_1_5_4_n4)
         );
  OR3_X1 npu_inst_pe_1_5_4_U27 ( .A1(npu_inst_pe_1_5_4_n5), .A2(
        npu_inst_pe_1_5_4_n7), .A3(npu_inst_pe_1_5_4_n4), .ZN(
        npu_inst_pe_1_5_4_n56) );
  OR3_X1 npu_inst_pe_1_5_4_U26 ( .A1(npu_inst_pe_1_5_4_n4), .A2(
        npu_inst_pe_1_5_4_n7), .A3(npu_inst_pe_1_5_4_n6), .ZN(
        npu_inst_pe_1_5_4_n48) );
  INV_X1 npu_inst_pe_1_5_4_U25 ( .A(npu_inst_pe_1_5_4_n4), .ZN(
        npu_inst_pe_1_5_4_n3) );
  OR3_X1 npu_inst_pe_1_5_4_U24 ( .A1(npu_inst_pe_1_5_4_n3), .A2(
        npu_inst_pe_1_5_4_n7), .A3(npu_inst_pe_1_5_4_n6), .ZN(
        npu_inst_pe_1_5_4_n52) );
  OR3_X1 npu_inst_pe_1_5_4_U23 ( .A1(npu_inst_pe_1_5_4_n5), .A2(
        npu_inst_pe_1_5_4_n7), .A3(npu_inst_pe_1_5_4_n3), .ZN(
        npu_inst_pe_1_5_4_n60) );
  BUF_X1 npu_inst_pe_1_5_4_U22 ( .A(npu_inst_n17), .Z(npu_inst_pe_1_5_4_n1) );
  NOR2_X1 npu_inst_pe_1_5_4_U21 ( .A1(npu_inst_pe_1_5_4_n60), .A2(
        npu_inst_pe_1_5_4_n2), .ZN(npu_inst_pe_1_5_4_n58) );
  NOR2_X1 npu_inst_pe_1_5_4_U20 ( .A1(npu_inst_pe_1_5_4_n56), .A2(
        npu_inst_pe_1_5_4_n2), .ZN(npu_inst_pe_1_5_4_n54) );
  NOR2_X1 npu_inst_pe_1_5_4_U19 ( .A1(npu_inst_pe_1_5_4_n52), .A2(
        npu_inst_pe_1_5_4_n2), .ZN(npu_inst_pe_1_5_4_n50) );
  NOR2_X1 npu_inst_pe_1_5_4_U18 ( .A1(npu_inst_pe_1_5_4_n48), .A2(
        npu_inst_pe_1_5_4_n2), .ZN(npu_inst_pe_1_5_4_n46) );
  NOR2_X1 npu_inst_pe_1_5_4_U17 ( .A1(npu_inst_pe_1_5_4_n40), .A2(
        npu_inst_pe_1_5_4_n2), .ZN(npu_inst_pe_1_5_4_n38) );
  NOR2_X1 npu_inst_pe_1_5_4_U16 ( .A1(npu_inst_pe_1_5_4_n44), .A2(
        npu_inst_pe_1_5_4_n2), .ZN(npu_inst_pe_1_5_4_n42) );
  BUF_X1 npu_inst_pe_1_5_4_U15 ( .A(npu_inst_n78), .Z(npu_inst_pe_1_5_4_n7) );
  INV_X1 npu_inst_pe_1_5_4_U14 ( .A(npu_inst_n105), .ZN(npu_inst_pe_1_5_4_n11)
         );
  INV_X1 npu_inst_pe_1_5_4_U13 ( .A(npu_inst_pe_1_5_4_n38), .ZN(
        npu_inst_pe_1_5_4_n113) );
  INV_X1 npu_inst_pe_1_5_4_U12 ( .A(npu_inst_pe_1_5_4_n58), .ZN(
        npu_inst_pe_1_5_4_n118) );
  INV_X1 npu_inst_pe_1_5_4_U11 ( .A(npu_inst_pe_1_5_4_n54), .ZN(
        npu_inst_pe_1_5_4_n117) );
  INV_X1 npu_inst_pe_1_5_4_U10 ( .A(npu_inst_pe_1_5_4_n50), .ZN(
        npu_inst_pe_1_5_4_n116) );
  INV_X1 npu_inst_pe_1_5_4_U9 ( .A(npu_inst_pe_1_5_4_n46), .ZN(
        npu_inst_pe_1_5_4_n115) );
  INV_X1 npu_inst_pe_1_5_4_U8 ( .A(npu_inst_pe_1_5_4_n42), .ZN(
        npu_inst_pe_1_5_4_n114) );
  BUF_X1 npu_inst_pe_1_5_4_U7 ( .A(npu_inst_pe_1_5_4_n11), .Z(
        npu_inst_pe_1_5_4_n10) );
  BUF_X1 npu_inst_pe_1_5_4_U6 ( .A(npu_inst_pe_1_5_4_n11), .Z(
        npu_inst_pe_1_5_4_n9) );
  BUF_X1 npu_inst_pe_1_5_4_U5 ( .A(npu_inst_pe_1_5_4_n11), .Z(
        npu_inst_pe_1_5_4_n8) );
  NOR2_X1 npu_inst_pe_1_5_4_U4 ( .A1(npu_inst_pe_1_5_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_4_n1), .ZN(npu_inst_pe_1_5_4_n76) );
  NOR2_X1 npu_inst_pe_1_5_4_U3 ( .A1(npu_inst_pe_1_5_4_n27), .A2(
        npu_inst_pe_1_5_4_n1), .ZN(npu_inst_pe_1_5_4_n77) );
  FA_X1 npu_inst_pe_1_5_4_sub_77_U2_1 ( .A(npu_inst_int_data_res_5__4__1_), 
        .B(npu_inst_pe_1_5_4_n13), .CI(npu_inst_pe_1_5_4_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_5_4_sub_77_carry_2_), .S(npu_inst_pe_1_5_4_N66) );
  FA_X1 npu_inst_pe_1_5_4_add_79_U1_1 ( .A(npu_inst_int_data_res_5__4__1_), 
        .B(npu_inst_pe_1_5_4_int_data_1_), .CI(
        npu_inst_pe_1_5_4_add_79_carry_1_), .CO(
        npu_inst_pe_1_5_4_add_79_carry_2_), .S(npu_inst_pe_1_5_4_N74) );
  NAND3_X1 npu_inst_pe_1_5_4_U101 ( .A1(npu_inst_pe_1_5_4_n4), .A2(
        npu_inst_pe_1_5_4_n6), .A3(npu_inst_pe_1_5_4_n7), .ZN(
        npu_inst_pe_1_5_4_n44) );
  NAND3_X1 npu_inst_pe_1_5_4_U100 ( .A1(npu_inst_pe_1_5_4_n3), .A2(
        npu_inst_pe_1_5_4_n6), .A3(npu_inst_pe_1_5_4_n7), .ZN(
        npu_inst_pe_1_5_4_n40) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_4_n33), .CK(
        npu_inst_pe_1_5_4_net3466), .RN(npu_inst_pe_1_5_4_n8), .Q(
        npu_inst_int_data_res_5__4__6_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_4_n34), .CK(
        npu_inst_pe_1_5_4_net3466), .RN(npu_inst_pe_1_5_4_n8), .Q(
        npu_inst_int_data_res_5__4__5_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_4_n35), .CK(
        npu_inst_pe_1_5_4_net3466), .RN(npu_inst_pe_1_5_4_n8), .Q(
        npu_inst_int_data_res_5__4__4_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_4_n36), .CK(
        npu_inst_pe_1_5_4_net3466), .RN(npu_inst_pe_1_5_4_n8), .Q(
        npu_inst_int_data_res_5__4__3_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_4_n98), .CK(
        npu_inst_pe_1_5_4_net3466), .RN(npu_inst_pe_1_5_4_n8), .Q(
        npu_inst_int_data_res_5__4__2_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_4_n99), .CK(
        npu_inst_pe_1_5_4_net3466), .RN(npu_inst_pe_1_5_4_n8), .Q(
        npu_inst_int_data_res_5__4__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_4_n32), .CK(
        npu_inst_pe_1_5_4_net3466), .RN(npu_inst_pe_1_5_4_n8), .Q(
        npu_inst_int_data_res_5__4__7_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_4_n100), 
        .CK(npu_inst_pe_1_5_4_net3466), .RN(npu_inst_pe_1_5_4_n8), .Q(
        npu_inst_int_data_res_5__4__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_weight_reg_0_ ( .D(npu_inst_n91), .CK(
        npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n8), .Q(
        npu_inst_pe_1_5_4_int_q_weight_0_), .QN(npu_inst_pe_1_5_4_n27) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_weight_reg_1_ ( .D(npu_inst_n97), .CK(
        npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n8), .Q(
        npu_inst_pe_1_5_4_int_q_weight_1_), .QN(npu_inst_pe_1_5_4_n26) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_4_n112), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n8), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_4_n106), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n8), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_4_n111), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_4_n105), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_4_n110), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_4_n104), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_4_n109), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_4_n103), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_4_n108), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_4_n102), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_4_n107), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_4_n101), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_4_n86), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_4_n87), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n9), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_4_n88), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_4_n89), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_4_n90), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_4_n91), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_4_n92), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_4_n93), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_4_n94), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_4_n95), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_4_n96), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_4_n97), 
        .CK(npu_inst_pe_1_5_4_net3472), .RN(npu_inst_pe_1_5_4_n10), .Q(
        npu_inst_pe_1_5_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_4_net3466) );
  CLKGATETST_X1 npu_inst_pe_1_5_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n44), .SE(1'b0), .GCK(npu_inst_pe_1_5_4_net3472) );
  MUX2_X1 npu_inst_pe_1_5_5_U153 ( .A(npu_inst_pe_1_5_5_n31), .B(
        npu_inst_pe_1_5_5_n28), .S(npu_inst_pe_1_5_5_n7), .Z(
        npu_inst_pe_1_5_5_N93) );
  MUX2_X1 npu_inst_pe_1_5_5_U152 ( .A(npu_inst_pe_1_5_5_n30), .B(
        npu_inst_pe_1_5_5_n29), .S(npu_inst_pe_1_5_5_n5), .Z(
        npu_inst_pe_1_5_5_n31) );
  MUX2_X1 npu_inst_pe_1_5_5_U151 ( .A(npu_inst_pe_1_5_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_5_n3), .Z(
        npu_inst_pe_1_5_5_n30) );
  MUX2_X1 npu_inst_pe_1_5_5_U150 ( .A(npu_inst_pe_1_5_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_5_n3), .Z(
        npu_inst_pe_1_5_5_n29) );
  MUX2_X1 npu_inst_pe_1_5_5_U149 ( .A(npu_inst_pe_1_5_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_5_n3), .Z(
        npu_inst_pe_1_5_5_n28) );
  MUX2_X1 npu_inst_pe_1_5_5_U148 ( .A(npu_inst_pe_1_5_5_n25), .B(
        npu_inst_pe_1_5_5_n22), .S(npu_inst_pe_1_5_5_n7), .Z(
        npu_inst_pe_1_5_5_N94) );
  MUX2_X1 npu_inst_pe_1_5_5_U147 ( .A(npu_inst_pe_1_5_5_n24), .B(
        npu_inst_pe_1_5_5_n23), .S(npu_inst_pe_1_5_5_n5), .Z(
        npu_inst_pe_1_5_5_n25) );
  MUX2_X1 npu_inst_pe_1_5_5_U146 ( .A(npu_inst_pe_1_5_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_5_n3), .Z(
        npu_inst_pe_1_5_5_n24) );
  MUX2_X1 npu_inst_pe_1_5_5_U145 ( .A(npu_inst_pe_1_5_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_5_n3), .Z(
        npu_inst_pe_1_5_5_n23) );
  MUX2_X1 npu_inst_pe_1_5_5_U144 ( .A(npu_inst_pe_1_5_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_5_n3), .Z(
        npu_inst_pe_1_5_5_n22) );
  MUX2_X1 npu_inst_pe_1_5_5_U143 ( .A(npu_inst_pe_1_5_5_n21), .B(
        npu_inst_pe_1_5_5_n18), .S(npu_inst_pe_1_5_5_n7), .Z(
        npu_inst_int_data_x_5__5__1_) );
  MUX2_X1 npu_inst_pe_1_5_5_U142 ( .A(npu_inst_pe_1_5_5_n20), .B(
        npu_inst_pe_1_5_5_n19), .S(npu_inst_pe_1_5_5_n5), .Z(
        npu_inst_pe_1_5_5_n21) );
  MUX2_X1 npu_inst_pe_1_5_5_U141 ( .A(npu_inst_pe_1_5_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_5_n3), .Z(
        npu_inst_pe_1_5_5_n20) );
  MUX2_X1 npu_inst_pe_1_5_5_U140 ( .A(npu_inst_pe_1_5_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_5_n3), .Z(
        npu_inst_pe_1_5_5_n19) );
  MUX2_X1 npu_inst_pe_1_5_5_U139 ( .A(npu_inst_pe_1_5_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_5_n3), .Z(
        npu_inst_pe_1_5_5_n18) );
  MUX2_X1 npu_inst_pe_1_5_5_U138 ( .A(npu_inst_pe_1_5_5_n17), .B(
        npu_inst_pe_1_5_5_n14), .S(npu_inst_pe_1_5_5_n7), .Z(
        npu_inst_int_data_x_5__5__0_) );
  MUX2_X1 npu_inst_pe_1_5_5_U137 ( .A(npu_inst_pe_1_5_5_n16), .B(
        npu_inst_pe_1_5_5_n15), .S(npu_inst_pe_1_5_5_n5), .Z(
        npu_inst_pe_1_5_5_n17) );
  MUX2_X1 npu_inst_pe_1_5_5_U136 ( .A(npu_inst_pe_1_5_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_5_n3), .Z(
        npu_inst_pe_1_5_5_n16) );
  MUX2_X1 npu_inst_pe_1_5_5_U135 ( .A(npu_inst_pe_1_5_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_5_n3), .Z(
        npu_inst_pe_1_5_5_n15) );
  MUX2_X1 npu_inst_pe_1_5_5_U134 ( .A(npu_inst_pe_1_5_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_5_n3), .Z(
        npu_inst_pe_1_5_5_n14) );
  XOR2_X1 npu_inst_pe_1_5_5_U133 ( .A(npu_inst_pe_1_5_5_int_data_0_), .B(
        npu_inst_int_data_res_5__5__0_), .Z(npu_inst_pe_1_5_5_N73) );
  AND2_X1 npu_inst_pe_1_5_5_U132 ( .A1(npu_inst_int_data_res_5__5__0_), .A2(
        npu_inst_pe_1_5_5_int_data_0_), .ZN(npu_inst_pe_1_5_5_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_5_U131 ( .A(npu_inst_int_data_res_5__5__0_), .B(
        npu_inst_pe_1_5_5_n12), .ZN(npu_inst_pe_1_5_5_N65) );
  OR2_X1 npu_inst_pe_1_5_5_U130 ( .A1(npu_inst_pe_1_5_5_n12), .A2(
        npu_inst_int_data_res_5__5__0_), .ZN(npu_inst_pe_1_5_5_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_5_U129 ( .A(npu_inst_int_data_res_5__5__2_), .B(
        npu_inst_pe_1_5_5_add_79_carry_2_), .Z(npu_inst_pe_1_5_5_N75) );
  AND2_X1 npu_inst_pe_1_5_5_U128 ( .A1(npu_inst_pe_1_5_5_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_5__5__2_), .ZN(
        npu_inst_pe_1_5_5_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_5_U127 ( .A(npu_inst_int_data_res_5__5__3_), .B(
        npu_inst_pe_1_5_5_add_79_carry_3_), .Z(npu_inst_pe_1_5_5_N76) );
  AND2_X1 npu_inst_pe_1_5_5_U126 ( .A1(npu_inst_pe_1_5_5_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_5__5__3_), .ZN(
        npu_inst_pe_1_5_5_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_5_U125 ( .A(npu_inst_int_data_res_5__5__4_), .B(
        npu_inst_pe_1_5_5_add_79_carry_4_), .Z(npu_inst_pe_1_5_5_N77) );
  AND2_X1 npu_inst_pe_1_5_5_U124 ( .A1(npu_inst_pe_1_5_5_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_5__5__4_), .ZN(
        npu_inst_pe_1_5_5_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_5_U123 ( .A(npu_inst_int_data_res_5__5__5_), .B(
        npu_inst_pe_1_5_5_add_79_carry_5_), .Z(npu_inst_pe_1_5_5_N78) );
  AND2_X1 npu_inst_pe_1_5_5_U122 ( .A1(npu_inst_pe_1_5_5_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_5__5__5_), .ZN(
        npu_inst_pe_1_5_5_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_5_U121 ( .A(npu_inst_int_data_res_5__5__6_), .B(
        npu_inst_pe_1_5_5_add_79_carry_6_), .Z(npu_inst_pe_1_5_5_N79) );
  AND2_X1 npu_inst_pe_1_5_5_U120 ( .A1(npu_inst_pe_1_5_5_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_5__5__6_), .ZN(
        npu_inst_pe_1_5_5_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_5_U119 ( .A(npu_inst_int_data_res_5__5__7_), .B(
        npu_inst_pe_1_5_5_add_79_carry_7_), .Z(npu_inst_pe_1_5_5_N80) );
  XNOR2_X1 npu_inst_pe_1_5_5_U118 ( .A(npu_inst_pe_1_5_5_sub_77_carry_2_), .B(
        npu_inst_int_data_res_5__5__2_), .ZN(npu_inst_pe_1_5_5_N67) );
  OR2_X1 npu_inst_pe_1_5_5_U117 ( .A1(npu_inst_int_data_res_5__5__2_), .A2(
        npu_inst_pe_1_5_5_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_5_5_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_5_U116 ( .A(npu_inst_pe_1_5_5_sub_77_carry_3_), .B(
        npu_inst_int_data_res_5__5__3_), .ZN(npu_inst_pe_1_5_5_N68) );
  OR2_X1 npu_inst_pe_1_5_5_U115 ( .A1(npu_inst_int_data_res_5__5__3_), .A2(
        npu_inst_pe_1_5_5_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_5_5_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_5_U114 ( .A(npu_inst_pe_1_5_5_sub_77_carry_4_), .B(
        npu_inst_int_data_res_5__5__4_), .ZN(npu_inst_pe_1_5_5_N69) );
  OR2_X1 npu_inst_pe_1_5_5_U113 ( .A1(npu_inst_int_data_res_5__5__4_), .A2(
        npu_inst_pe_1_5_5_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_5_5_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_5_U112 ( .A(npu_inst_pe_1_5_5_sub_77_carry_5_), .B(
        npu_inst_int_data_res_5__5__5_), .ZN(npu_inst_pe_1_5_5_N70) );
  OR2_X1 npu_inst_pe_1_5_5_U111 ( .A1(npu_inst_int_data_res_5__5__5_), .A2(
        npu_inst_pe_1_5_5_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_5_5_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_5_U110 ( .A(npu_inst_pe_1_5_5_sub_77_carry_6_), .B(
        npu_inst_int_data_res_5__5__6_), .ZN(npu_inst_pe_1_5_5_N71) );
  OR2_X1 npu_inst_pe_1_5_5_U109 ( .A1(npu_inst_int_data_res_5__5__6_), .A2(
        npu_inst_pe_1_5_5_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_5_5_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_5_U108 ( .A(npu_inst_int_data_res_5__5__7_), .B(
        npu_inst_pe_1_5_5_sub_77_carry_7_), .ZN(npu_inst_pe_1_5_5_N72) );
  INV_X1 npu_inst_pe_1_5_5_U107 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_5_5_n6)
         );
  INV_X1 npu_inst_pe_1_5_5_U106 ( .A(npu_inst_pe_1_5_5_n6), .ZN(
        npu_inst_pe_1_5_5_n5) );
  INV_X1 npu_inst_pe_1_5_5_U105 ( .A(npu_inst_n36), .ZN(npu_inst_pe_1_5_5_n2)
         );
  AOI22_X1 npu_inst_pe_1_5_5_U104 ( .A1(npu_inst_int_data_y_6__5__0_), .A2(
        npu_inst_pe_1_5_5_n58), .B1(npu_inst_pe_1_5_5_n118), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_5_n57) );
  INV_X1 npu_inst_pe_1_5_5_U103 ( .A(npu_inst_pe_1_5_5_n57), .ZN(
        npu_inst_pe_1_5_5_n107) );
  AOI22_X1 npu_inst_pe_1_5_5_U102 ( .A1(npu_inst_int_data_y_6__5__0_), .A2(
        npu_inst_pe_1_5_5_n54), .B1(npu_inst_pe_1_5_5_n117), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_5_n53) );
  INV_X1 npu_inst_pe_1_5_5_U99 ( .A(npu_inst_pe_1_5_5_n53), .ZN(
        npu_inst_pe_1_5_5_n108) );
  AOI22_X1 npu_inst_pe_1_5_5_U98 ( .A1(npu_inst_int_data_y_6__5__0_), .A2(
        npu_inst_pe_1_5_5_n50), .B1(npu_inst_pe_1_5_5_n116), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_5_n49) );
  INV_X1 npu_inst_pe_1_5_5_U97 ( .A(npu_inst_pe_1_5_5_n49), .ZN(
        npu_inst_pe_1_5_5_n109) );
  AOI22_X1 npu_inst_pe_1_5_5_U96 ( .A1(npu_inst_int_data_y_6__5__0_), .A2(
        npu_inst_pe_1_5_5_n46), .B1(npu_inst_pe_1_5_5_n115), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_5_n45) );
  INV_X1 npu_inst_pe_1_5_5_U95 ( .A(npu_inst_pe_1_5_5_n45), .ZN(
        npu_inst_pe_1_5_5_n110) );
  AOI22_X1 npu_inst_pe_1_5_5_U94 ( .A1(npu_inst_int_data_y_6__5__0_), .A2(
        npu_inst_pe_1_5_5_n42), .B1(npu_inst_pe_1_5_5_n114), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_5_n41) );
  INV_X1 npu_inst_pe_1_5_5_U93 ( .A(npu_inst_pe_1_5_5_n41), .ZN(
        npu_inst_pe_1_5_5_n111) );
  AOI22_X1 npu_inst_pe_1_5_5_U92 ( .A1(npu_inst_int_data_y_6__5__1_), .A2(
        npu_inst_pe_1_5_5_n58), .B1(npu_inst_pe_1_5_5_n118), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_5_n59) );
  INV_X1 npu_inst_pe_1_5_5_U91 ( .A(npu_inst_pe_1_5_5_n59), .ZN(
        npu_inst_pe_1_5_5_n101) );
  AOI22_X1 npu_inst_pe_1_5_5_U90 ( .A1(npu_inst_int_data_y_6__5__1_), .A2(
        npu_inst_pe_1_5_5_n54), .B1(npu_inst_pe_1_5_5_n117), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_5_n55) );
  INV_X1 npu_inst_pe_1_5_5_U89 ( .A(npu_inst_pe_1_5_5_n55), .ZN(
        npu_inst_pe_1_5_5_n102) );
  AOI22_X1 npu_inst_pe_1_5_5_U88 ( .A1(npu_inst_int_data_y_6__5__1_), .A2(
        npu_inst_pe_1_5_5_n50), .B1(npu_inst_pe_1_5_5_n116), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_5_n51) );
  INV_X1 npu_inst_pe_1_5_5_U87 ( .A(npu_inst_pe_1_5_5_n51), .ZN(
        npu_inst_pe_1_5_5_n103) );
  AOI22_X1 npu_inst_pe_1_5_5_U86 ( .A1(npu_inst_int_data_y_6__5__1_), .A2(
        npu_inst_pe_1_5_5_n46), .B1(npu_inst_pe_1_5_5_n115), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_5_n47) );
  INV_X1 npu_inst_pe_1_5_5_U85 ( .A(npu_inst_pe_1_5_5_n47), .ZN(
        npu_inst_pe_1_5_5_n104) );
  AOI22_X1 npu_inst_pe_1_5_5_U84 ( .A1(npu_inst_int_data_y_6__5__1_), .A2(
        npu_inst_pe_1_5_5_n42), .B1(npu_inst_pe_1_5_5_n114), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_5_n43) );
  INV_X1 npu_inst_pe_1_5_5_U83 ( .A(npu_inst_pe_1_5_5_n43), .ZN(
        npu_inst_pe_1_5_5_n105) );
  AOI22_X1 npu_inst_pe_1_5_5_U82 ( .A1(npu_inst_pe_1_5_5_n38), .A2(
        npu_inst_int_data_y_6__5__1_), .B1(npu_inst_pe_1_5_5_n113), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_5_n39) );
  INV_X1 npu_inst_pe_1_5_5_U81 ( .A(npu_inst_pe_1_5_5_n39), .ZN(
        npu_inst_pe_1_5_5_n106) );
  AND2_X1 npu_inst_pe_1_5_5_U80 ( .A1(npu_inst_pe_1_5_5_N93), .A2(npu_inst_n36), .ZN(npu_inst_int_data_y_5__5__0_) );
  NAND2_X1 npu_inst_pe_1_5_5_U79 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_5_n60), .ZN(npu_inst_pe_1_5_5_n74) );
  OAI21_X1 npu_inst_pe_1_5_5_U78 ( .B1(npu_inst_pe_1_5_5_n63), .B2(
        npu_inst_pe_1_5_5_n60), .A(npu_inst_pe_1_5_5_n74), .ZN(
        npu_inst_pe_1_5_5_n97) );
  NAND2_X1 npu_inst_pe_1_5_5_U77 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_5_n60), .ZN(npu_inst_pe_1_5_5_n73) );
  OAI21_X1 npu_inst_pe_1_5_5_U76 ( .B1(npu_inst_pe_1_5_5_n61), .B2(
        npu_inst_pe_1_5_5_n60), .A(npu_inst_pe_1_5_5_n73), .ZN(
        npu_inst_pe_1_5_5_n96) );
  NAND2_X1 npu_inst_pe_1_5_5_U75 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_5_n56), .ZN(npu_inst_pe_1_5_5_n72) );
  OAI21_X1 npu_inst_pe_1_5_5_U74 ( .B1(npu_inst_pe_1_5_5_n63), .B2(
        npu_inst_pe_1_5_5_n56), .A(npu_inst_pe_1_5_5_n72), .ZN(
        npu_inst_pe_1_5_5_n95) );
  NAND2_X1 npu_inst_pe_1_5_5_U73 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_5_n56), .ZN(npu_inst_pe_1_5_5_n71) );
  OAI21_X1 npu_inst_pe_1_5_5_U72 ( .B1(npu_inst_pe_1_5_5_n61), .B2(
        npu_inst_pe_1_5_5_n56), .A(npu_inst_pe_1_5_5_n71), .ZN(
        npu_inst_pe_1_5_5_n94) );
  NAND2_X1 npu_inst_pe_1_5_5_U71 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_5_n52), .ZN(npu_inst_pe_1_5_5_n70) );
  OAI21_X1 npu_inst_pe_1_5_5_U70 ( .B1(npu_inst_pe_1_5_5_n63), .B2(
        npu_inst_pe_1_5_5_n52), .A(npu_inst_pe_1_5_5_n70), .ZN(
        npu_inst_pe_1_5_5_n93) );
  NAND2_X1 npu_inst_pe_1_5_5_U69 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_5_n52), .ZN(npu_inst_pe_1_5_5_n69) );
  OAI21_X1 npu_inst_pe_1_5_5_U68 ( .B1(npu_inst_pe_1_5_5_n61), .B2(
        npu_inst_pe_1_5_5_n52), .A(npu_inst_pe_1_5_5_n69), .ZN(
        npu_inst_pe_1_5_5_n92) );
  NAND2_X1 npu_inst_pe_1_5_5_U67 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_5_n48), .ZN(npu_inst_pe_1_5_5_n68) );
  OAI21_X1 npu_inst_pe_1_5_5_U66 ( .B1(npu_inst_pe_1_5_5_n63), .B2(
        npu_inst_pe_1_5_5_n48), .A(npu_inst_pe_1_5_5_n68), .ZN(
        npu_inst_pe_1_5_5_n91) );
  NAND2_X1 npu_inst_pe_1_5_5_U65 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_5_n48), .ZN(npu_inst_pe_1_5_5_n67) );
  OAI21_X1 npu_inst_pe_1_5_5_U64 ( .B1(npu_inst_pe_1_5_5_n61), .B2(
        npu_inst_pe_1_5_5_n48), .A(npu_inst_pe_1_5_5_n67), .ZN(
        npu_inst_pe_1_5_5_n90) );
  NAND2_X1 npu_inst_pe_1_5_5_U63 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_5_n44), .ZN(npu_inst_pe_1_5_5_n66) );
  OAI21_X1 npu_inst_pe_1_5_5_U62 ( .B1(npu_inst_pe_1_5_5_n63), .B2(
        npu_inst_pe_1_5_5_n44), .A(npu_inst_pe_1_5_5_n66), .ZN(
        npu_inst_pe_1_5_5_n89) );
  NAND2_X1 npu_inst_pe_1_5_5_U61 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_5_n44), .ZN(npu_inst_pe_1_5_5_n65) );
  OAI21_X1 npu_inst_pe_1_5_5_U60 ( .B1(npu_inst_pe_1_5_5_n61), .B2(
        npu_inst_pe_1_5_5_n44), .A(npu_inst_pe_1_5_5_n65), .ZN(
        npu_inst_pe_1_5_5_n88) );
  NAND2_X1 npu_inst_pe_1_5_5_U59 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_5_n40), .ZN(npu_inst_pe_1_5_5_n64) );
  OAI21_X1 npu_inst_pe_1_5_5_U58 ( .B1(npu_inst_pe_1_5_5_n63), .B2(
        npu_inst_pe_1_5_5_n40), .A(npu_inst_pe_1_5_5_n64), .ZN(
        npu_inst_pe_1_5_5_n87) );
  NAND2_X1 npu_inst_pe_1_5_5_U57 ( .A1(npu_inst_pe_1_5_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_5_n40), .ZN(npu_inst_pe_1_5_5_n62) );
  OAI21_X1 npu_inst_pe_1_5_5_U56 ( .B1(npu_inst_pe_1_5_5_n61), .B2(
        npu_inst_pe_1_5_5_n40), .A(npu_inst_pe_1_5_5_n62), .ZN(
        npu_inst_pe_1_5_5_n86) );
  AOI22_X1 npu_inst_pe_1_5_5_U55 ( .A1(npu_inst_pe_1_5_5_n38), .A2(
        npu_inst_int_data_y_6__5__0_), .B1(npu_inst_pe_1_5_5_n113), .B2(
        npu_inst_pe_1_5_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_5_n37) );
  INV_X1 npu_inst_pe_1_5_5_U54 ( .A(npu_inst_pe_1_5_5_n37), .ZN(
        npu_inst_pe_1_5_5_n112) );
  AND2_X1 npu_inst_pe_1_5_5_U53 ( .A1(npu_inst_n36), .A2(npu_inst_pe_1_5_5_N94), .ZN(npu_inst_int_data_y_5__5__1_) );
  AOI222_X1 npu_inst_pe_1_5_5_U52 ( .A1(npu_inst_int_data_res_6__5__0_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N73), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N65), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n84) );
  INV_X1 npu_inst_pe_1_5_5_U51 ( .A(npu_inst_pe_1_5_5_n84), .ZN(
        npu_inst_pe_1_5_5_n100) );
  AOI222_X1 npu_inst_pe_1_5_5_U50 ( .A1(npu_inst_pe_1_5_5_n1), .A2(
        npu_inst_int_data_res_6__5__7_), .B1(npu_inst_pe_1_5_5_N80), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N72), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n75) );
  INV_X1 npu_inst_pe_1_5_5_U49 ( .A(npu_inst_pe_1_5_5_n75), .ZN(
        npu_inst_pe_1_5_5_n32) );
  AOI222_X1 npu_inst_pe_1_5_5_U48 ( .A1(npu_inst_int_data_res_6__5__1_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N74), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N66), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n83) );
  INV_X1 npu_inst_pe_1_5_5_U47 ( .A(npu_inst_pe_1_5_5_n83), .ZN(
        npu_inst_pe_1_5_5_n99) );
  AOI222_X1 npu_inst_pe_1_5_5_U46 ( .A1(npu_inst_int_data_res_6__5__3_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N76), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N68), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n81) );
  INV_X1 npu_inst_pe_1_5_5_U45 ( .A(npu_inst_pe_1_5_5_n81), .ZN(
        npu_inst_pe_1_5_5_n36) );
  AOI222_X1 npu_inst_pe_1_5_5_U44 ( .A1(npu_inst_int_data_res_6__5__4_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N77), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N69), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n80) );
  INV_X1 npu_inst_pe_1_5_5_U43 ( .A(npu_inst_pe_1_5_5_n80), .ZN(
        npu_inst_pe_1_5_5_n35) );
  AOI222_X1 npu_inst_pe_1_5_5_U42 ( .A1(npu_inst_int_data_res_6__5__5_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N78), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N70), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n79) );
  INV_X1 npu_inst_pe_1_5_5_U41 ( .A(npu_inst_pe_1_5_5_n79), .ZN(
        npu_inst_pe_1_5_5_n34) );
  AOI222_X1 npu_inst_pe_1_5_5_U40 ( .A1(npu_inst_int_data_res_6__5__6_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N79), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N71), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n78) );
  INV_X1 npu_inst_pe_1_5_5_U39 ( .A(npu_inst_pe_1_5_5_n78), .ZN(
        npu_inst_pe_1_5_5_n33) );
  NOR3_X1 npu_inst_pe_1_5_5_U38 ( .A1(npu_inst_pe_1_5_5_n26), .A2(npu_inst_n36), .A3(npu_inst_int_ckg[18]), .ZN(npu_inst_pe_1_5_5_n85) );
  OR2_X1 npu_inst_pe_1_5_5_U37 ( .A1(npu_inst_pe_1_5_5_n85), .A2(
        npu_inst_pe_1_5_5_n1), .ZN(npu_inst_pe_1_5_5_N84) );
  AND2_X1 npu_inst_pe_1_5_5_U36 ( .A1(npu_inst_int_data_x_5__5__1_), .A2(
        npu_inst_pe_1_5_5_int_q_weight_1_), .ZN(npu_inst_pe_1_5_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_5_U35 ( .A1(npu_inst_int_data_x_5__5__0_), .A2(
        npu_inst_pe_1_5_5_int_q_weight_1_), .ZN(npu_inst_pe_1_5_5_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_5_5_U34 ( .A(npu_inst_pe_1_5_5_int_data_1_), .ZN(
        npu_inst_pe_1_5_5_n13) );
  AOI222_X1 npu_inst_pe_1_5_5_U33 ( .A1(npu_inst_int_data_res_6__5__2_), .A2(
        npu_inst_pe_1_5_5_n1), .B1(npu_inst_pe_1_5_5_N75), .B2(
        npu_inst_pe_1_5_5_n76), .C1(npu_inst_pe_1_5_5_N67), .C2(
        npu_inst_pe_1_5_5_n77), .ZN(npu_inst_pe_1_5_5_n82) );
  INV_X1 npu_inst_pe_1_5_5_U32 ( .A(npu_inst_pe_1_5_5_n82), .ZN(
        npu_inst_pe_1_5_5_n98) );
  AOI22_X1 npu_inst_pe_1_5_5_U31 ( .A1(npu_inst_n36), .A2(
        npu_inst_int_data_y_6__5__1_), .B1(npu_inst_pe_1_5_5_n2), .B2(
        npu_inst_int_data_x_5__6__1_), .ZN(npu_inst_pe_1_5_5_n63) );
  AOI22_X1 npu_inst_pe_1_5_5_U30 ( .A1(npu_inst_n36), .A2(
        npu_inst_int_data_y_6__5__0_), .B1(npu_inst_pe_1_5_5_n2), .B2(
        npu_inst_int_data_x_5__6__0_), .ZN(npu_inst_pe_1_5_5_n61) );
  INV_X1 npu_inst_pe_1_5_5_U29 ( .A(npu_inst_pe_1_5_5_int_data_0_), .ZN(
        npu_inst_pe_1_5_5_n12) );
  INV_X1 npu_inst_pe_1_5_5_U28 ( .A(npu_inst_n50), .ZN(npu_inst_pe_1_5_5_n4)
         );
  OR3_X1 npu_inst_pe_1_5_5_U27 ( .A1(npu_inst_pe_1_5_5_n5), .A2(
        npu_inst_pe_1_5_5_n7), .A3(npu_inst_pe_1_5_5_n4), .ZN(
        npu_inst_pe_1_5_5_n56) );
  OR3_X1 npu_inst_pe_1_5_5_U26 ( .A1(npu_inst_pe_1_5_5_n4), .A2(
        npu_inst_pe_1_5_5_n7), .A3(npu_inst_pe_1_5_5_n6), .ZN(
        npu_inst_pe_1_5_5_n48) );
  INV_X1 npu_inst_pe_1_5_5_U25 ( .A(npu_inst_pe_1_5_5_n4), .ZN(
        npu_inst_pe_1_5_5_n3) );
  OR3_X1 npu_inst_pe_1_5_5_U24 ( .A1(npu_inst_pe_1_5_5_n3), .A2(
        npu_inst_pe_1_5_5_n7), .A3(npu_inst_pe_1_5_5_n6), .ZN(
        npu_inst_pe_1_5_5_n52) );
  OR3_X1 npu_inst_pe_1_5_5_U23 ( .A1(npu_inst_pe_1_5_5_n5), .A2(
        npu_inst_pe_1_5_5_n7), .A3(npu_inst_pe_1_5_5_n3), .ZN(
        npu_inst_pe_1_5_5_n60) );
  BUF_X1 npu_inst_pe_1_5_5_U22 ( .A(npu_inst_n17), .Z(npu_inst_pe_1_5_5_n1) );
  NOR2_X1 npu_inst_pe_1_5_5_U21 ( .A1(npu_inst_pe_1_5_5_n60), .A2(
        npu_inst_pe_1_5_5_n2), .ZN(npu_inst_pe_1_5_5_n58) );
  NOR2_X1 npu_inst_pe_1_5_5_U20 ( .A1(npu_inst_pe_1_5_5_n56), .A2(
        npu_inst_pe_1_5_5_n2), .ZN(npu_inst_pe_1_5_5_n54) );
  NOR2_X1 npu_inst_pe_1_5_5_U19 ( .A1(npu_inst_pe_1_5_5_n52), .A2(
        npu_inst_pe_1_5_5_n2), .ZN(npu_inst_pe_1_5_5_n50) );
  NOR2_X1 npu_inst_pe_1_5_5_U18 ( .A1(npu_inst_pe_1_5_5_n48), .A2(
        npu_inst_pe_1_5_5_n2), .ZN(npu_inst_pe_1_5_5_n46) );
  NOR2_X1 npu_inst_pe_1_5_5_U17 ( .A1(npu_inst_pe_1_5_5_n40), .A2(
        npu_inst_pe_1_5_5_n2), .ZN(npu_inst_pe_1_5_5_n38) );
  NOR2_X1 npu_inst_pe_1_5_5_U16 ( .A1(npu_inst_pe_1_5_5_n44), .A2(
        npu_inst_pe_1_5_5_n2), .ZN(npu_inst_pe_1_5_5_n42) );
  BUF_X1 npu_inst_pe_1_5_5_U15 ( .A(npu_inst_n78), .Z(npu_inst_pe_1_5_5_n7) );
  INV_X1 npu_inst_pe_1_5_5_U14 ( .A(npu_inst_n105), .ZN(npu_inst_pe_1_5_5_n11)
         );
  INV_X1 npu_inst_pe_1_5_5_U13 ( .A(npu_inst_pe_1_5_5_n38), .ZN(
        npu_inst_pe_1_5_5_n113) );
  INV_X1 npu_inst_pe_1_5_5_U12 ( .A(npu_inst_pe_1_5_5_n58), .ZN(
        npu_inst_pe_1_5_5_n118) );
  INV_X1 npu_inst_pe_1_5_5_U11 ( .A(npu_inst_pe_1_5_5_n54), .ZN(
        npu_inst_pe_1_5_5_n117) );
  INV_X1 npu_inst_pe_1_5_5_U10 ( .A(npu_inst_pe_1_5_5_n50), .ZN(
        npu_inst_pe_1_5_5_n116) );
  INV_X1 npu_inst_pe_1_5_5_U9 ( .A(npu_inst_pe_1_5_5_n46), .ZN(
        npu_inst_pe_1_5_5_n115) );
  INV_X1 npu_inst_pe_1_5_5_U8 ( .A(npu_inst_pe_1_5_5_n42), .ZN(
        npu_inst_pe_1_5_5_n114) );
  BUF_X1 npu_inst_pe_1_5_5_U7 ( .A(npu_inst_pe_1_5_5_n11), .Z(
        npu_inst_pe_1_5_5_n10) );
  BUF_X1 npu_inst_pe_1_5_5_U6 ( .A(npu_inst_pe_1_5_5_n11), .Z(
        npu_inst_pe_1_5_5_n9) );
  BUF_X1 npu_inst_pe_1_5_5_U5 ( .A(npu_inst_pe_1_5_5_n11), .Z(
        npu_inst_pe_1_5_5_n8) );
  NOR2_X1 npu_inst_pe_1_5_5_U4 ( .A1(npu_inst_pe_1_5_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_5_n1), .ZN(npu_inst_pe_1_5_5_n76) );
  NOR2_X1 npu_inst_pe_1_5_5_U3 ( .A1(npu_inst_pe_1_5_5_n27), .A2(
        npu_inst_pe_1_5_5_n1), .ZN(npu_inst_pe_1_5_5_n77) );
  FA_X1 npu_inst_pe_1_5_5_sub_77_U2_1 ( .A(npu_inst_int_data_res_5__5__1_), 
        .B(npu_inst_pe_1_5_5_n13), .CI(npu_inst_pe_1_5_5_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_5_5_sub_77_carry_2_), .S(npu_inst_pe_1_5_5_N66) );
  FA_X1 npu_inst_pe_1_5_5_add_79_U1_1 ( .A(npu_inst_int_data_res_5__5__1_), 
        .B(npu_inst_pe_1_5_5_int_data_1_), .CI(
        npu_inst_pe_1_5_5_add_79_carry_1_), .CO(
        npu_inst_pe_1_5_5_add_79_carry_2_), .S(npu_inst_pe_1_5_5_N74) );
  NAND3_X1 npu_inst_pe_1_5_5_U101 ( .A1(npu_inst_pe_1_5_5_n4), .A2(
        npu_inst_pe_1_5_5_n6), .A3(npu_inst_pe_1_5_5_n7), .ZN(
        npu_inst_pe_1_5_5_n44) );
  NAND3_X1 npu_inst_pe_1_5_5_U100 ( .A1(npu_inst_pe_1_5_5_n3), .A2(
        npu_inst_pe_1_5_5_n6), .A3(npu_inst_pe_1_5_5_n7), .ZN(
        npu_inst_pe_1_5_5_n40) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_5_n33), .CK(
        npu_inst_pe_1_5_5_net3443), .RN(npu_inst_pe_1_5_5_n8), .Q(
        npu_inst_int_data_res_5__5__6_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_5_n34), .CK(
        npu_inst_pe_1_5_5_net3443), .RN(npu_inst_pe_1_5_5_n8), .Q(
        npu_inst_int_data_res_5__5__5_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_5_n35), .CK(
        npu_inst_pe_1_5_5_net3443), .RN(npu_inst_pe_1_5_5_n8), .Q(
        npu_inst_int_data_res_5__5__4_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_5_n36), .CK(
        npu_inst_pe_1_5_5_net3443), .RN(npu_inst_pe_1_5_5_n8), .Q(
        npu_inst_int_data_res_5__5__3_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_5_n98), .CK(
        npu_inst_pe_1_5_5_net3443), .RN(npu_inst_pe_1_5_5_n8), .Q(
        npu_inst_int_data_res_5__5__2_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_5_n99), .CK(
        npu_inst_pe_1_5_5_net3443), .RN(npu_inst_pe_1_5_5_n8), .Q(
        npu_inst_int_data_res_5__5__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_5_n32), .CK(
        npu_inst_pe_1_5_5_net3443), .RN(npu_inst_pe_1_5_5_n8), .Q(
        npu_inst_int_data_res_5__5__7_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_5_n100), 
        .CK(npu_inst_pe_1_5_5_net3443), .RN(npu_inst_pe_1_5_5_n8), .Q(
        npu_inst_int_data_res_5__5__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_weight_reg_0_ ( .D(npu_inst_n91), .CK(
        npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n8), .Q(
        npu_inst_pe_1_5_5_int_q_weight_0_), .QN(npu_inst_pe_1_5_5_n27) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_weight_reg_1_ ( .D(npu_inst_n97), .CK(
        npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n8), .Q(
        npu_inst_pe_1_5_5_int_q_weight_1_), .QN(npu_inst_pe_1_5_5_n26) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_5_n112), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n8), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_5_n106), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n8), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_5_n111), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_5_n105), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_5_n110), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_5_n104), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_5_n109), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_5_n103), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_5_n108), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_5_n102), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_5_n107), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_5_n101), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_5_n86), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_5_n87), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n9), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_5_n88), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_5_n89), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_5_n90), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_5_n91), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_5_n92), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_5_n93), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_5_n94), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_5_n95), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_5_n96), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_5_n97), 
        .CK(npu_inst_pe_1_5_5_net3449), .RN(npu_inst_pe_1_5_5_n10), .Q(
        npu_inst_pe_1_5_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_5_net3443) );
  CLKGATETST_X1 npu_inst_pe_1_5_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n44), .SE(1'b0), .GCK(npu_inst_pe_1_5_5_net3449) );
  MUX2_X1 npu_inst_pe_1_5_6_U153 ( .A(npu_inst_pe_1_5_6_n31), .B(
        npu_inst_pe_1_5_6_n28), .S(npu_inst_pe_1_5_6_n7), .Z(
        npu_inst_pe_1_5_6_N93) );
  MUX2_X1 npu_inst_pe_1_5_6_U152 ( .A(npu_inst_pe_1_5_6_n30), .B(
        npu_inst_pe_1_5_6_n29), .S(npu_inst_pe_1_5_6_n5), .Z(
        npu_inst_pe_1_5_6_n31) );
  MUX2_X1 npu_inst_pe_1_5_6_U151 ( .A(npu_inst_pe_1_5_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_6_n3), .Z(
        npu_inst_pe_1_5_6_n30) );
  MUX2_X1 npu_inst_pe_1_5_6_U150 ( .A(npu_inst_pe_1_5_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_6_n3), .Z(
        npu_inst_pe_1_5_6_n29) );
  MUX2_X1 npu_inst_pe_1_5_6_U149 ( .A(npu_inst_pe_1_5_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_6_n3), .Z(
        npu_inst_pe_1_5_6_n28) );
  MUX2_X1 npu_inst_pe_1_5_6_U148 ( .A(npu_inst_pe_1_5_6_n25), .B(
        npu_inst_pe_1_5_6_n22), .S(npu_inst_pe_1_5_6_n7), .Z(
        npu_inst_pe_1_5_6_N94) );
  MUX2_X1 npu_inst_pe_1_5_6_U147 ( .A(npu_inst_pe_1_5_6_n24), .B(
        npu_inst_pe_1_5_6_n23), .S(npu_inst_pe_1_5_6_n5), .Z(
        npu_inst_pe_1_5_6_n25) );
  MUX2_X1 npu_inst_pe_1_5_6_U146 ( .A(npu_inst_pe_1_5_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_6_n3), .Z(
        npu_inst_pe_1_5_6_n24) );
  MUX2_X1 npu_inst_pe_1_5_6_U145 ( .A(npu_inst_pe_1_5_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_6_n3), .Z(
        npu_inst_pe_1_5_6_n23) );
  MUX2_X1 npu_inst_pe_1_5_6_U144 ( .A(npu_inst_pe_1_5_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_6_n3), .Z(
        npu_inst_pe_1_5_6_n22) );
  MUX2_X1 npu_inst_pe_1_5_6_U143 ( .A(npu_inst_pe_1_5_6_n21), .B(
        npu_inst_pe_1_5_6_n18), .S(npu_inst_pe_1_5_6_n7), .Z(
        npu_inst_int_data_x_5__6__1_) );
  MUX2_X1 npu_inst_pe_1_5_6_U142 ( .A(npu_inst_pe_1_5_6_n20), .B(
        npu_inst_pe_1_5_6_n19), .S(npu_inst_pe_1_5_6_n5), .Z(
        npu_inst_pe_1_5_6_n21) );
  MUX2_X1 npu_inst_pe_1_5_6_U141 ( .A(npu_inst_pe_1_5_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_6_n3), .Z(
        npu_inst_pe_1_5_6_n20) );
  MUX2_X1 npu_inst_pe_1_5_6_U140 ( .A(npu_inst_pe_1_5_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_6_n3), .Z(
        npu_inst_pe_1_5_6_n19) );
  MUX2_X1 npu_inst_pe_1_5_6_U139 ( .A(npu_inst_pe_1_5_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_6_n3), .Z(
        npu_inst_pe_1_5_6_n18) );
  MUX2_X1 npu_inst_pe_1_5_6_U138 ( .A(npu_inst_pe_1_5_6_n17), .B(
        npu_inst_pe_1_5_6_n14), .S(npu_inst_pe_1_5_6_n7), .Z(
        npu_inst_int_data_x_5__6__0_) );
  MUX2_X1 npu_inst_pe_1_5_6_U137 ( .A(npu_inst_pe_1_5_6_n16), .B(
        npu_inst_pe_1_5_6_n15), .S(npu_inst_pe_1_5_6_n5), .Z(
        npu_inst_pe_1_5_6_n17) );
  MUX2_X1 npu_inst_pe_1_5_6_U136 ( .A(npu_inst_pe_1_5_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_6_n3), .Z(
        npu_inst_pe_1_5_6_n16) );
  MUX2_X1 npu_inst_pe_1_5_6_U135 ( .A(npu_inst_pe_1_5_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_6_n3), .Z(
        npu_inst_pe_1_5_6_n15) );
  MUX2_X1 npu_inst_pe_1_5_6_U134 ( .A(npu_inst_pe_1_5_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_6_n3), .Z(
        npu_inst_pe_1_5_6_n14) );
  XOR2_X1 npu_inst_pe_1_5_6_U133 ( .A(npu_inst_pe_1_5_6_int_data_0_), .B(
        npu_inst_int_data_res_5__6__0_), .Z(npu_inst_pe_1_5_6_N73) );
  AND2_X1 npu_inst_pe_1_5_6_U132 ( .A1(npu_inst_int_data_res_5__6__0_), .A2(
        npu_inst_pe_1_5_6_int_data_0_), .ZN(npu_inst_pe_1_5_6_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_6_U131 ( .A(npu_inst_int_data_res_5__6__0_), .B(
        npu_inst_pe_1_5_6_n12), .ZN(npu_inst_pe_1_5_6_N65) );
  OR2_X1 npu_inst_pe_1_5_6_U130 ( .A1(npu_inst_pe_1_5_6_n12), .A2(
        npu_inst_int_data_res_5__6__0_), .ZN(npu_inst_pe_1_5_6_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_6_U129 ( .A(npu_inst_int_data_res_5__6__2_), .B(
        npu_inst_pe_1_5_6_add_79_carry_2_), .Z(npu_inst_pe_1_5_6_N75) );
  AND2_X1 npu_inst_pe_1_5_6_U128 ( .A1(npu_inst_pe_1_5_6_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_5__6__2_), .ZN(
        npu_inst_pe_1_5_6_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_6_U127 ( .A(npu_inst_int_data_res_5__6__3_), .B(
        npu_inst_pe_1_5_6_add_79_carry_3_), .Z(npu_inst_pe_1_5_6_N76) );
  AND2_X1 npu_inst_pe_1_5_6_U126 ( .A1(npu_inst_pe_1_5_6_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_5__6__3_), .ZN(
        npu_inst_pe_1_5_6_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_6_U125 ( .A(npu_inst_int_data_res_5__6__4_), .B(
        npu_inst_pe_1_5_6_add_79_carry_4_), .Z(npu_inst_pe_1_5_6_N77) );
  AND2_X1 npu_inst_pe_1_5_6_U124 ( .A1(npu_inst_pe_1_5_6_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_5__6__4_), .ZN(
        npu_inst_pe_1_5_6_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_6_U123 ( .A(npu_inst_int_data_res_5__6__5_), .B(
        npu_inst_pe_1_5_6_add_79_carry_5_), .Z(npu_inst_pe_1_5_6_N78) );
  AND2_X1 npu_inst_pe_1_5_6_U122 ( .A1(npu_inst_pe_1_5_6_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_5__6__5_), .ZN(
        npu_inst_pe_1_5_6_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_6_U121 ( .A(npu_inst_int_data_res_5__6__6_), .B(
        npu_inst_pe_1_5_6_add_79_carry_6_), .Z(npu_inst_pe_1_5_6_N79) );
  AND2_X1 npu_inst_pe_1_5_6_U120 ( .A1(npu_inst_pe_1_5_6_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_5__6__6_), .ZN(
        npu_inst_pe_1_5_6_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_6_U119 ( .A(npu_inst_int_data_res_5__6__7_), .B(
        npu_inst_pe_1_5_6_add_79_carry_7_), .Z(npu_inst_pe_1_5_6_N80) );
  XNOR2_X1 npu_inst_pe_1_5_6_U118 ( .A(npu_inst_pe_1_5_6_sub_77_carry_2_), .B(
        npu_inst_int_data_res_5__6__2_), .ZN(npu_inst_pe_1_5_6_N67) );
  OR2_X1 npu_inst_pe_1_5_6_U117 ( .A1(npu_inst_int_data_res_5__6__2_), .A2(
        npu_inst_pe_1_5_6_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_5_6_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_6_U116 ( .A(npu_inst_pe_1_5_6_sub_77_carry_3_), .B(
        npu_inst_int_data_res_5__6__3_), .ZN(npu_inst_pe_1_5_6_N68) );
  OR2_X1 npu_inst_pe_1_5_6_U115 ( .A1(npu_inst_int_data_res_5__6__3_), .A2(
        npu_inst_pe_1_5_6_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_5_6_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_6_U114 ( .A(npu_inst_pe_1_5_6_sub_77_carry_4_), .B(
        npu_inst_int_data_res_5__6__4_), .ZN(npu_inst_pe_1_5_6_N69) );
  OR2_X1 npu_inst_pe_1_5_6_U113 ( .A1(npu_inst_int_data_res_5__6__4_), .A2(
        npu_inst_pe_1_5_6_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_5_6_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_6_U112 ( .A(npu_inst_pe_1_5_6_sub_77_carry_5_), .B(
        npu_inst_int_data_res_5__6__5_), .ZN(npu_inst_pe_1_5_6_N70) );
  OR2_X1 npu_inst_pe_1_5_6_U111 ( .A1(npu_inst_int_data_res_5__6__5_), .A2(
        npu_inst_pe_1_5_6_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_5_6_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_6_U110 ( .A(npu_inst_pe_1_5_6_sub_77_carry_6_), .B(
        npu_inst_int_data_res_5__6__6_), .ZN(npu_inst_pe_1_5_6_N71) );
  OR2_X1 npu_inst_pe_1_5_6_U109 ( .A1(npu_inst_int_data_res_5__6__6_), .A2(
        npu_inst_pe_1_5_6_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_5_6_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_6_U108 ( .A(npu_inst_int_data_res_5__6__7_), .B(
        npu_inst_pe_1_5_6_sub_77_carry_7_), .ZN(npu_inst_pe_1_5_6_N72) );
  INV_X1 npu_inst_pe_1_5_6_U107 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_5_6_n6)
         );
  INV_X1 npu_inst_pe_1_5_6_U106 ( .A(npu_inst_pe_1_5_6_n6), .ZN(
        npu_inst_pe_1_5_6_n5) );
  INV_X1 npu_inst_pe_1_5_6_U105 ( .A(npu_inst_n36), .ZN(npu_inst_pe_1_5_6_n2)
         );
  AOI22_X1 npu_inst_pe_1_5_6_U104 ( .A1(npu_inst_int_data_y_6__6__0_), .A2(
        npu_inst_pe_1_5_6_n58), .B1(npu_inst_pe_1_5_6_n118), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_6_n57) );
  INV_X1 npu_inst_pe_1_5_6_U103 ( .A(npu_inst_pe_1_5_6_n57), .ZN(
        npu_inst_pe_1_5_6_n107) );
  AOI22_X1 npu_inst_pe_1_5_6_U102 ( .A1(npu_inst_int_data_y_6__6__0_), .A2(
        npu_inst_pe_1_5_6_n54), .B1(npu_inst_pe_1_5_6_n117), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_6_n53) );
  INV_X1 npu_inst_pe_1_5_6_U99 ( .A(npu_inst_pe_1_5_6_n53), .ZN(
        npu_inst_pe_1_5_6_n108) );
  AOI22_X1 npu_inst_pe_1_5_6_U98 ( .A1(npu_inst_int_data_y_6__6__0_), .A2(
        npu_inst_pe_1_5_6_n50), .B1(npu_inst_pe_1_5_6_n116), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_6_n49) );
  INV_X1 npu_inst_pe_1_5_6_U97 ( .A(npu_inst_pe_1_5_6_n49), .ZN(
        npu_inst_pe_1_5_6_n109) );
  AOI22_X1 npu_inst_pe_1_5_6_U96 ( .A1(npu_inst_int_data_y_6__6__0_), .A2(
        npu_inst_pe_1_5_6_n46), .B1(npu_inst_pe_1_5_6_n115), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_6_n45) );
  INV_X1 npu_inst_pe_1_5_6_U95 ( .A(npu_inst_pe_1_5_6_n45), .ZN(
        npu_inst_pe_1_5_6_n110) );
  AOI22_X1 npu_inst_pe_1_5_6_U94 ( .A1(npu_inst_int_data_y_6__6__0_), .A2(
        npu_inst_pe_1_5_6_n42), .B1(npu_inst_pe_1_5_6_n114), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_6_n41) );
  INV_X1 npu_inst_pe_1_5_6_U93 ( .A(npu_inst_pe_1_5_6_n41), .ZN(
        npu_inst_pe_1_5_6_n111) );
  AOI22_X1 npu_inst_pe_1_5_6_U92 ( .A1(npu_inst_int_data_y_6__6__1_), .A2(
        npu_inst_pe_1_5_6_n58), .B1(npu_inst_pe_1_5_6_n118), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_6_n59) );
  INV_X1 npu_inst_pe_1_5_6_U91 ( .A(npu_inst_pe_1_5_6_n59), .ZN(
        npu_inst_pe_1_5_6_n101) );
  AOI22_X1 npu_inst_pe_1_5_6_U90 ( .A1(npu_inst_int_data_y_6__6__1_), .A2(
        npu_inst_pe_1_5_6_n54), .B1(npu_inst_pe_1_5_6_n117), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_6_n55) );
  INV_X1 npu_inst_pe_1_5_6_U89 ( .A(npu_inst_pe_1_5_6_n55), .ZN(
        npu_inst_pe_1_5_6_n102) );
  AOI22_X1 npu_inst_pe_1_5_6_U88 ( .A1(npu_inst_int_data_y_6__6__1_), .A2(
        npu_inst_pe_1_5_6_n50), .B1(npu_inst_pe_1_5_6_n116), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_6_n51) );
  INV_X1 npu_inst_pe_1_5_6_U87 ( .A(npu_inst_pe_1_5_6_n51), .ZN(
        npu_inst_pe_1_5_6_n103) );
  AOI22_X1 npu_inst_pe_1_5_6_U86 ( .A1(npu_inst_int_data_y_6__6__1_), .A2(
        npu_inst_pe_1_5_6_n46), .B1(npu_inst_pe_1_5_6_n115), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_6_n47) );
  INV_X1 npu_inst_pe_1_5_6_U85 ( .A(npu_inst_pe_1_5_6_n47), .ZN(
        npu_inst_pe_1_5_6_n104) );
  AOI22_X1 npu_inst_pe_1_5_6_U84 ( .A1(npu_inst_int_data_y_6__6__1_), .A2(
        npu_inst_pe_1_5_6_n42), .B1(npu_inst_pe_1_5_6_n114), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_6_n43) );
  INV_X1 npu_inst_pe_1_5_6_U83 ( .A(npu_inst_pe_1_5_6_n43), .ZN(
        npu_inst_pe_1_5_6_n105) );
  AOI22_X1 npu_inst_pe_1_5_6_U82 ( .A1(npu_inst_pe_1_5_6_n38), .A2(
        npu_inst_int_data_y_6__6__1_), .B1(npu_inst_pe_1_5_6_n113), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_6_n39) );
  INV_X1 npu_inst_pe_1_5_6_U81 ( .A(npu_inst_pe_1_5_6_n39), .ZN(
        npu_inst_pe_1_5_6_n106) );
  AND2_X1 npu_inst_pe_1_5_6_U80 ( .A1(npu_inst_pe_1_5_6_N93), .A2(npu_inst_n36), .ZN(npu_inst_int_data_y_5__6__0_) );
  NAND2_X1 npu_inst_pe_1_5_6_U79 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_6_n60), .ZN(npu_inst_pe_1_5_6_n74) );
  OAI21_X1 npu_inst_pe_1_5_6_U78 ( .B1(npu_inst_pe_1_5_6_n63), .B2(
        npu_inst_pe_1_5_6_n60), .A(npu_inst_pe_1_5_6_n74), .ZN(
        npu_inst_pe_1_5_6_n97) );
  NAND2_X1 npu_inst_pe_1_5_6_U77 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_6_n60), .ZN(npu_inst_pe_1_5_6_n73) );
  OAI21_X1 npu_inst_pe_1_5_6_U76 ( .B1(npu_inst_pe_1_5_6_n61), .B2(
        npu_inst_pe_1_5_6_n60), .A(npu_inst_pe_1_5_6_n73), .ZN(
        npu_inst_pe_1_5_6_n96) );
  NAND2_X1 npu_inst_pe_1_5_6_U75 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_6_n56), .ZN(npu_inst_pe_1_5_6_n72) );
  OAI21_X1 npu_inst_pe_1_5_6_U74 ( .B1(npu_inst_pe_1_5_6_n63), .B2(
        npu_inst_pe_1_5_6_n56), .A(npu_inst_pe_1_5_6_n72), .ZN(
        npu_inst_pe_1_5_6_n95) );
  NAND2_X1 npu_inst_pe_1_5_6_U73 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_6_n56), .ZN(npu_inst_pe_1_5_6_n71) );
  OAI21_X1 npu_inst_pe_1_5_6_U72 ( .B1(npu_inst_pe_1_5_6_n61), .B2(
        npu_inst_pe_1_5_6_n56), .A(npu_inst_pe_1_5_6_n71), .ZN(
        npu_inst_pe_1_5_6_n94) );
  NAND2_X1 npu_inst_pe_1_5_6_U71 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_6_n52), .ZN(npu_inst_pe_1_5_6_n70) );
  OAI21_X1 npu_inst_pe_1_5_6_U70 ( .B1(npu_inst_pe_1_5_6_n63), .B2(
        npu_inst_pe_1_5_6_n52), .A(npu_inst_pe_1_5_6_n70), .ZN(
        npu_inst_pe_1_5_6_n93) );
  NAND2_X1 npu_inst_pe_1_5_6_U69 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_6_n52), .ZN(npu_inst_pe_1_5_6_n69) );
  OAI21_X1 npu_inst_pe_1_5_6_U68 ( .B1(npu_inst_pe_1_5_6_n61), .B2(
        npu_inst_pe_1_5_6_n52), .A(npu_inst_pe_1_5_6_n69), .ZN(
        npu_inst_pe_1_5_6_n92) );
  NAND2_X1 npu_inst_pe_1_5_6_U67 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_6_n48), .ZN(npu_inst_pe_1_5_6_n68) );
  OAI21_X1 npu_inst_pe_1_5_6_U66 ( .B1(npu_inst_pe_1_5_6_n63), .B2(
        npu_inst_pe_1_5_6_n48), .A(npu_inst_pe_1_5_6_n68), .ZN(
        npu_inst_pe_1_5_6_n91) );
  NAND2_X1 npu_inst_pe_1_5_6_U65 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_6_n48), .ZN(npu_inst_pe_1_5_6_n67) );
  OAI21_X1 npu_inst_pe_1_5_6_U64 ( .B1(npu_inst_pe_1_5_6_n61), .B2(
        npu_inst_pe_1_5_6_n48), .A(npu_inst_pe_1_5_6_n67), .ZN(
        npu_inst_pe_1_5_6_n90) );
  NAND2_X1 npu_inst_pe_1_5_6_U63 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_6_n44), .ZN(npu_inst_pe_1_5_6_n66) );
  OAI21_X1 npu_inst_pe_1_5_6_U62 ( .B1(npu_inst_pe_1_5_6_n63), .B2(
        npu_inst_pe_1_5_6_n44), .A(npu_inst_pe_1_5_6_n66), .ZN(
        npu_inst_pe_1_5_6_n89) );
  NAND2_X1 npu_inst_pe_1_5_6_U61 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_6_n44), .ZN(npu_inst_pe_1_5_6_n65) );
  OAI21_X1 npu_inst_pe_1_5_6_U60 ( .B1(npu_inst_pe_1_5_6_n61), .B2(
        npu_inst_pe_1_5_6_n44), .A(npu_inst_pe_1_5_6_n65), .ZN(
        npu_inst_pe_1_5_6_n88) );
  NAND2_X1 npu_inst_pe_1_5_6_U59 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_6_n40), .ZN(npu_inst_pe_1_5_6_n64) );
  OAI21_X1 npu_inst_pe_1_5_6_U58 ( .B1(npu_inst_pe_1_5_6_n63), .B2(
        npu_inst_pe_1_5_6_n40), .A(npu_inst_pe_1_5_6_n64), .ZN(
        npu_inst_pe_1_5_6_n87) );
  NAND2_X1 npu_inst_pe_1_5_6_U57 ( .A1(npu_inst_pe_1_5_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_6_n40), .ZN(npu_inst_pe_1_5_6_n62) );
  OAI21_X1 npu_inst_pe_1_5_6_U56 ( .B1(npu_inst_pe_1_5_6_n61), .B2(
        npu_inst_pe_1_5_6_n40), .A(npu_inst_pe_1_5_6_n62), .ZN(
        npu_inst_pe_1_5_6_n86) );
  AOI22_X1 npu_inst_pe_1_5_6_U55 ( .A1(npu_inst_pe_1_5_6_n38), .A2(
        npu_inst_int_data_y_6__6__0_), .B1(npu_inst_pe_1_5_6_n113), .B2(
        npu_inst_pe_1_5_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_6_n37) );
  INV_X1 npu_inst_pe_1_5_6_U54 ( .A(npu_inst_pe_1_5_6_n37), .ZN(
        npu_inst_pe_1_5_6_n112) );
  AND2_X1 npu_inst_pe_1_5_6_U53 ( .A1(npu_inst_n36), .A2(npu_inst_pe_1_5_6_N94), .ZN(npu_inst_int_data_y_5__6__1_) );
  AOI222_X1 npu_inst_pe_1_5_6_U52 ( .A1(npu_inst_int_data_res_6__6__0_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N73), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N65), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n84) );
  INV_X1 npu_inst_pe_1_5_6_U51 ( .A(npu_inst_pe_1_5_6_n84), .ZN(
        npu_inst_pe_1_5_6_n100) );
  AOI222_X1 npu_inst_pe_1_5_6_U50 ( .A1(npu_inst_pe_1_5_6_n1), .A2(
        npu_inst_int_data_res_6__6__7_), .B1(npu_inst_pe_1_5_6_N80), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N72), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n75) );
  INV_X1 npu_inst_pe_1_5_6_U49 ( .A(npu_inst_pe_1_5_6_n75), .ZN(
        npu_inst_pe_1_5_6_n32) );
  AOI222_X1 npu_inst_pe_1_5_6_U48 ( .A1(npu_inst_int_data_res_6__6__1_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N74), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N66), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n83) );
  INV_X1 npu_inst_pe_1_5_6_U47 ( .A(npu_inst_pe_1_5_6_n83), .ZN(
        npu_inst_pe_1_5_6_n99) );
  AOI222_X1 npu_inst_pe_1_5_6_U46 ( .A1(npu_inst_int_data_res_6__6__3_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N76), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N68), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n81) );
  INV_X1 npu_inst_pe_1_5_6_U45 ( .A(npu_inst_pe_1_5_6_n81), .ZN(
        npu_inst_pe_1_5_6_n36) );
  AOI222_X1 npu_inst_pe_1_5_6_U44 ( .A1(npu_inst_int_data_res_6__6__4_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N77), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N69), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n80) );
  INV_X1 npu_inst_pe_1_5_6_U43 ( .A(npu_inst_pe_1_5_6_n80), .ZN(
        npu_inst_pe_1_5_6_n35) );
  AOI222_X1 npu_inst_pe_1_5_6_U42 ( .A1(npu_inst_int_data_res_6__6__5_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N78), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N70), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n79) );
  INV_X1 npu_inst_pe_1_5_6_U41 ( .A(npu_inst_pe_1_5_6_n79), .ZN(
        npu_inst_pe_1_5_6_n34) );
  AOI222_X1 npu_inst_pe_1_5_6_U40 ( .A1(npu_inst_int_data_res_6__6__6_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N79), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N71), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n78) );
  INV_X1 npu_inst_pe_1_5_6_U39 ( .A(npu_inst_pe_1_5_6_n78), .ZN(
        npu_inst_pe_1_5_6_n33) );
  NOR3_X1 npu_inst_pe_1_5_6_U38 ( .A1(npu_inst_pe_1_5_6_n26), .A2(npu_inst_n36), .A3(npu_inst_int_ckg[17]), .ZN(npu_inst_pe_1_5_6_n85) );
  OR2_X1 npu_inst_pe_1_5_6_U37 ( .A1(npu_inst_pe_1_5_6_n85), .A2(
        npu_inst_pe_1_5_6_n1), .ZN(npu_inst_pe_1_5_6_N84) );
  AND2_X1 npu_inst_pe_1_5_6_U36 ( .A1(npu_inst_int_data_x_5__6__1_), .A2(
        npu_inst_pe_1_5_6_int_q_weight_1_), .ZN(npu_inst_pe_1_5_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_6_U35 ( .A1(npu_inst_int_data_x_5__6__0_), .A2(
        npu_inst_pe_1_5_6_int_q_weight_1_), .ZN(npu_inst_pe_1_5_6_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_5_6_U34 ( .A(npu_inst_pe_1_5_6_int_data_1_), .ZN(
        npu_inst_pe_1_5_6_n13) );
  AOI222_X1 npu_inst_pe_1_5_6_U33 ( .A1(npu_inst_int_data_res_6__6__2_), .A2(
        npu_inst_pe_1_5_6_n1), .B1(npu_inst_pe_1_5_6_N75), .B2(
        npu_inst_pe_1_5_6_n76), .C1(npu_inst_pe_1_5_6_N67), .C2(
        npu_inst_pe_1_5_6_n77), .ZN(npu_inst_pe_1_5_6_n82) );
  INV_X1 npu_inst_pe_1_5_6_U32 ( .A(npu_inst_pe_1_5_6_n82), .ZN(
        npu_inst_pe_1_5_6_n98) );
  AOI22_X1 npu_inst_pe_1_5_6_U31 ( .A1(npu_inst_n36), .A2(
        npu_inst_int_data_y_6__6__1_), .B1(npu_inst_pe_1_5_6_n2), .B2(
        npu_inst_int_data_x_5__7__1_), .ZN(npu_inst_pe_1_5_6_n63) );
  AOI22_X1 npu_inst_pe_1_5_6_U30 ( .A1(npu_inst_n36), .A2(
        npu_inst_int_data_y_6__6__0_), .B1(npu_inst_pe_1_5_6_n2), .B2(
        npu_inst_int_data_x_5__7__0_), .ZN(npu_inst_pe_1_5_6_n61) );
  INV_X1 npu_inst_pe_1_5_6_U29 ( .A(npu_inst_pe_1_5_6_int_data_0_), .ZN(
        npu_inst_pe_1_5_6_n12) );
  INV_X1 npu_inst_pe_1_5_6_U28 ( .A(npu_inst_n50), .ZN(npu_inst_pe_1_5_6_n4)
         );
  OR3_X1 npu_inst_pe_1_5_6_U27 ( .A1(npu_inst_pe_1_5_6_n5), .A2(
        npu_inst_pe_1_5_6_n7), .A3(npu_inst_pe_1_5_6_n4), .ZN(
        npu_inst_pe_1_5_6_n56) );
  OR3_X1 npu_inst_pe_1_5_6_U26 ( .A1(npu_inst_pe_1_5_6_n4), .A2(
        npu_inst_pe_1_5_6_n7), .A3(npu_inst_pe_1_5_6_n6), .ZN(
        npu_inst_pe_1_5_6_n48) );
  INV_X1 npu_inst_pe_1_5_6_U25 ( .A(npu_inst_pe_1_5_6_n4), .ZN(
        npu_inst_pe_1_5_6_n3) );
  OR3_X1 npu_inst_pe_1_5_6_U24 ( .A1(npu_inst_pe_1_5_6_n3), .A2(
        npu_inst_pe_1_5_6_n7), .A3(npu_inst_pe_1_5_6_n6), .ZN(
        npu_inst_pe_1_5_6_n52) );
  OR3_X1 npu_inst_pe_1_5_6_U23 ( .A1(npu_inst_pe_1_5_6_n5), .A2(
        npu_inst_pe_1_5_6_n7), .A3(npu_inst_pe_1_5_6_n3), .ZN(
        npu_inst_pe_1_5_6_n60) );
  BUF_X1 npu_inst_pe_1_5_6_U22 ( .A(npu_inst_n16), .Z(npu_inst_pe_1_5_6_n1) );
  NOR2_X1 npu_inst_pe_1_5_6_U21 ( .A1(npu_inst_pe_1_5_6_n60), .A2(
        npu_inst_pe_1_5_6_n2), .ZN(npu_inst_pe_1_5_6_n58) );
  NOR2_X1 npu_inst_pe_1_5_6_U20 ( .A1(npu_inst_pe_1_5_6_n56), .A2(
        npu_inst_pe_1_5_6_n2), .ZN(npu_inst_pe_1_5_6_n54) );
  NOR2_X1 npu_inst_pe_1_5_6_U19 ( .A1(npu_inst_pe_1_5_6_n52), .A2(
        npu_inst_pe_1_5_6_n2), .ZN(npu_inst_pe_1_5_6_n50) );
  NOR2_X1 npu_inst_pe_1_5_6_U18 ( .A1(npu_inst_pe_1_5_6_n48), .A2(
        npu_inst_pe_1_5_6_n2), .ZN(npu_inst_pe_1_5_6_n46) );
  NOR2_X1 npu_inst_pe_1_5_6_U17 ( .A1(npu_inst_pe_1_5_6_n40), .A2(
        npu_inst_pe_1_5_6_n2), .ZN(npu_inst_pe_1_5_6_n38) );
  NOR2_X1 npu_inst_pe_1_5_6_U16 ( .A1(npu_inst_pe_1_5_6_n44), .A2(
        npu_inst_pe_1_5_6_n2), .ZN(npu_inst_pe_1_5_6_n42) );
  BUF_X1 npu_inst_pe_1_5_6_U15 ( .A(npu_inst_n78), .Z(npu_inst_pe_1_5_6_n7) );
  INV_X1 npu_inst_pe_1_5_6_U14 ( .A(npu_inst_n105), .ZN(npu_inst_pe_1_5_6_n11)
         );
  INV_X1 npu_inst_pe_1_5_6_U13 ( .A(npu_inst_pe_1_5_6_n38), .ZN(
        npu_inst_pe_1_5_6_n113) );
  INV_X1 npu_inst_pe_1_5_6_U12 ( .A(npu_inst_pe_1_5_6_n58), .ZN(
        npu_inst_pe_1_5_6_n118) );
  INV_X1 npu_inst_pe_1_5_6_U11 ( .A(npu_inst_pe_1_5_6_n54), .ZN(
        npu_inst_pe_1_5_6_n117) );
  INV_X1 npu_inst_pe_1_5_6_U10 ( .A(npu_inst_pe_1_5_6_n50), .ZN(
        npu_inst_pe_1_5_6_n116) );
  INV_X1 npu_inst_pe_1_5_6_U9 ( .A(npu_inst_pe_1_5_6_n46), .ZN(
        npu_inst_pe_1_5_6_n115) );
  INV_X1 npu_inst_pe_1_5_6_U8 ( .A(npu_inst_pe_1_5_6_n42), .ZN(
        npu_inst_pe_1_5_6_n114) );
  BUF_X1 npu_inst_pe_1_5_6_U7 ( .A(npu_inst_pe_1_5_6_n11), .Z(
        npu_inst_pe_1_5_6_n10) );
  BUF_X1 npu_inst_pe_1_5_6_U6 ( .A(npu_inst_pe_1_5_6_n11), .Z(
        npu_inst_pe_1_5_6_n9) );
  BUF_X1 npu_inst_pe_1_5_6_U5 ( .A(npu_inst_pe_1_5_6_n11), .Z(
        npu_inst_pe_1_5_6_n8) );
  NOR2_X1 npu_inst_pe_1_5_6_U4 ( .A1(npu_inst_pe_1_5_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_6_n1), .ZN(npu_inst_pe_1_5_6_n76) );
  NOR2_X1 npu_inst_pe_1_5_6_U3 ( .A1(npu_inst_pe_1_5_6_n27), .A2(
        npu_inst_pe_1_5_6_n1), .ZN(npu_inst_pe_1_5_6_n77) );
  FA_X1 npu_inst_pe_1_5_6_sub_77_U2_1 ( .A(npu_inst_int_data_res_5__6__1_), 
        .B(npu_inst_pe_1_5_6_n13), .CI(npu_inst_pe_1_5_6_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_5_6_sub_77_carry_2_), .S(npu_inst_pe_1_5_6_N66) );
  FA_X1 npu_inst_pe_1_5_6_add_79_U1_1 ( .A(npu_inst_int_data_res_5__6__1_), 
        .B(npu_inst_pe_1_5_6_int_data_1_), .CI(
        npu_inst_pe_1_5_6_add_79_carry_1_), .CO(
        npu_inst_pe_1_5_6_add_79_carry_2_), .S(npu_inst_pe_1_5_6_N74) );
  NAND3_X1 npu_inst_pe_1_5_6_U101 ( .A1(npu_inst_pe_1_5_6_n4), .A2(
        npu_inst_pe_1_5_6_n6), .A3(npu_inst_pe_1_5_6_n7), .ZN(
        npu_inst_pe_1_5_6_n44) );
  NAND3_X1 npu_inst_pe_1_5_6_U100 ( .A1(npu_inst_pe_1_5_6_n3), .A2(
        npu_inst_pe_1_5_6_n6), .A3(npu_inst_pe_1_5_6_n7), .ZN(
        npu_inst_pe_1_5_6_n40) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_6_n33), .CK(
        npu_inst_pe_1_5_6_net3420), .RN(npu_inst_pe_1_5_6_n8), .Q(
        npu_inst_int_data_res_5__6__6_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_6_n34), .CK(
        npu_inst_pe_1_5_6_net3420), .RN(npu_inst_pe_1_5_6_n8), .Q(
        npu_inst_int_data_res_5__6__5_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_6_n35), .CK(
        npu_inst_pe_1_5_6_net3420), .RN(npu_inst_pe_1_5_6_n8), .Q(
        npu_inst_int_data_res_5__6__4_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_6_n36), .CK(
        npu_inst_pe_1_5_6_net3420), .RN(npu_inst_pe_1_5_6_n8), .Q(
        npu_inst_int_data_res_5__6__3_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_6_n98), .CK(
        npu_inst_pe_1_5_6_net3420), .RN(npu_inst_pe_1_5_6_n8), .Q(
        npu_inst_int_data_res_5__6__2_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_6_n99), .CK(
        npu_inst_pe_1_5_6_net3420), .RN(npu_inst_pe_1_5_6_n8), .Q(
        npu_inst_int_data_res_5__6__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_6_n32), .CK(
        npu_inst_pe_1_5_6_net3420), .RN(npu_inst_pe_1_5_6_n8), .Q(
        npu_inst_int_data_res_5__6__7_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_6_n100), 
        .CK(npu_inst_pe_1_5_6_net3420), .RN(npu_inst_pe_1_5_6_n8), .Q(
        npu_inst_int_data_res_5__6__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_weight_reg_0_ ( .D(npu_inst_n91), .CK(
        npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n8), .Q(
        npu_inst_pe_1_5_6_int_q_weight_0_), .QN(npu_inst_pe_1_5_6_n27) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_weight_reg_1_ ( .D(npu_inst_n97), .CK(
        npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n8), .Q(
        npu_inst_pe_1_5_6_int_q_weight_1_), .QN(npu_inst_pe_1_5_6_n26) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_6_n112), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n8), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_6_n106), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n8), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_6_n111), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_6_n105), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_6_n110), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_6_n104), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_6_n109), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_6_n103), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_6_n108), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_6_n102), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_6_n107), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_6_n101), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_6_n86), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_6_n87), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n9), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_6_n88), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_6_n89), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_6_n90), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_6_n91), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_6_n92), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_6_n93), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_6_n94), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_6_n95), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_6_n96), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_6_n97), 
        .CK(npu_inst_pe_1_5_6_net3426), .RN(npu_inst_pe_1_5_6_n10), .Q(
        npu_inst_pe_1_5_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_6_net3420) );
  CLKGATETST_X1 npu_inst_pe_1_5_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n44), .SE(1'b0), .GCK(npu_inst_pe_1_5_6_net3426) );
  MUX2_X1 npu_inst_pe_1_5_7_U153 ( .A(npu_inst_pe_1_5_7_n31), .B(
        npu_inst_pe_1_5_7_n28), .S(npu_inst_pe_1_5_7_n7), .Z(
        npu_inst_pe_1_5_7_N93) );
  MUX2_X1 npu_inst_pe_1_5_7_U152 ( .A(npu_inst_pe_1_5_7_n30), .B(
        npu_inst_pe_1_5_7_n29), .S(npu_inst_pe_1_5_7_n5), .Z(
        npu_inst_pe_1_5_7_n31) );
  MUX2_X1 npu_inst_pe_1_5_7_U151 ( .A(npu_inst_pe_1_5_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_5_7_n3), .Z(
        npu_inst_pe_1_5_7_n30) );
  MUX2_X1 npu_inst_pe_1_5_7_U150 ( .A(npu_inst_pe_1_5_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_5_7_n3), .Z(
        npu_inst_pe_1_5_7_n29) );
  MUX2_X1 npu_inst_pe_1_5_7_U149 ( .A(npu_inst_pe_1_5_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_5_7_n3), .Z(
        npu_inst_pe_1_5_7_n28) );
  MUX2_X1 npu_inst_pe_1_5_7_U148 ( .A(npu_inst_pe_1_5_7_n25), .B(
        npu_inst_pe_1_5_7_n22), .S(npu_inst_pe_1_5_7_n7), .Z(
        npu_inst_pe_1_5_7_N94) );
  MUX2_X1 npu_inst_pe_1_5_7_U147 ( .A(npu_inst_pe_1_5_7_n24), .B(
        npu_inst_pe_1_5_7_n23), .S(npu_inst_pe_1_5_7_n5), .Z(
        npu_inst_pe_1_5_7_n25) );
  MUX2_X1 npu_inst_pe_1_5_7_U146 ( .A(npu_inst_pe_1_5_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_5_7_n3), .Z(
        npu_inst_pe_1_5_7_n24) );
  MUX2_X1 npu_inst_pe_1_5_7_U145 ( .A(npu_inst_pe_1_5_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_5_7_n3), .Z(
        npu_inst_pe_1_5_7_n23) );
  MUX2_X1 npu_inst_pe_1_5_7_U144 ( .A(npu_inst_pe_1_5_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_5_7_n3), .Z(
        npu_inst_pe_1_5_7_n22) );
  MUX2_X1 npu_inst_pe_1_5_7_U143 ( .A(npu_inst_pe_1_5_7_n21), .B(
        npu_inst_pe_1_5_7_n18), .S(npu_inst_pe_1_5_7_n7), .Z(
        npu_inst_int_data_x_5__7__1_) );
  MUX2_X1 npu_inst_pe_1_5_7_U142 ( .A(npu_inst_pe_1_5_7_n20), .B(
        npu_inst_pe_1_5_7_n19), .S(npu_inst_pe_1_5_7_n5), .Z(
        npu_inst_pe_1_5_7_n21) );
  MUX2_X1 npu_inst_pe_1_5_7_U141 ( .A(npu_inst_pe_1_5_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_5_7_n3), .Z(
        npu_inst_pe_1_5_7_n20) );
  MUX2_X1 npu_inst_pe_1_5_7_U140 ( .A(npu_inst_pe_1_5_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_5_7_n3), .Z(
        npu_inst_pe_1_5_7_n19) );
  MUX2_X1 npu_inst_pe_1_5_7_U139 ( .A(npu_inst_pe_1_5_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_5_7_n3), .Z(
        npu_inst_pe_1_5_7_n18) );
  MUX2_X1 npu_inst_pe_1_5_7_U138 ( .A(npu_inst_pe_1_5_7_n17), .B(
        npu_inst_pe_1_5_7_n14), .S(npu_inst_pe_1_5_7_n7), .Z(
        npu_inst_int_data_x_5__7__0_) );
  MUX2_X1 npu_inst_pe_1_5_7_U137 ( .A(npu_inst_pe_1_5_7_n16), .B(
        npu_inst_pe_1_5_7_n15), .S(npu_inst_pe_1_5_7_n5), .Z(
        npu_inst_pe_1_5_7_n17) );
  MUX2_X1 npu_inst_pe_1_5_7_U136 ( .A(npu_inst_pe_1_5_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_5_7_n3), .Z(
        npu_inst_pe_1_5_7_n16) );
  MUX2_X1 npu_inst_pe_1_5_7_U135 ( .A(npu_inst_pe_1_5_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_5_7_n3), .Z(
        npu_inst_pe_1_5_7_n15) );
  MUX2_X1 npu_inst_pe_1_5_7_U134 ( .A(npu_inst_pe_1_5_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_5_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_5_7_n3), .Z(
        npu_inst_pe_1_5_7_n14) );
  XOR2_X1 npu_inst_pe_1_5_7_U133 ( .A(npu_inst_pe_1_5_7_int_data_0_), .B(
        npu_inst_int_data_res_5__7__0_), .Z(npu_inst_pe_1_5_7_N73) );
  AND2_X1 npu_inst_pe_1_5_7_U132 ( .A1(npu_inst_int_data_res_5__7__0_), .A2(
        npu_inst_pe_1_5_7_int_data_0_), .ZN(npu_inst_pe_1_5_7_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_5_7_U131 ( .A(npu_inst_int_data_res_5__7__0_), .B(
        npu_inst_pe_1_5_7_n12), .ZN(npu_inst_pe_1_5_7_N65) );
  OR2_X1 npu_inst_pe_1_5_7_U130 ( .A1(npu_inst_pe_1_5_7_n12), .A2(
        npu_inst_int_data_res_5__7__0_), .ZN(npu_inst_pe_1_5_7_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_5_7_U129 ( .A(npu_inst_int_data_res_5__7__2_), .B(
        npu_inst_pe_1_5_7_add_79_carry_2_), .Z(npu_inst_pe_1_5_7_N75) );
  AND2_X1 npu_inst_pe_1_5_7_U128 ( .A1(npu_inst_pe_1_5_7_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_5__7__2_), .ZN(
        npu_inst_pe_1_5_7_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_5_7_U127 ( .A(npu_inst_int_data_res_5__7__3_), .B(
        npu_inst_pe_1_5_7_add_79_carry_3_), .Z(npu_inst_pe_1_5_7_N76) );
  AND2_X1 npu_inst_pe_1_5_7_U126 ( .A1(npu_inst_pe_1_5_7_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_5__7__3_), .ZN(
        npu_inst_pe_1_5_7_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_5_7_U125 ( .A(npu_inst_int_data_res_5__7__4_), .B(
        npu_inst_pe_1_5_7_add_79_carry_4_), .Z(npu_inst_pe_1_5_7_N77) );
  AND2_X1 npu_inst_pe_1_5_7_U124 ( .A1(npu_inst_pe_1_5_7_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_5__7__4_), .ZN(
        npu_inst_pe_1_5_7_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_5_7_U123 ( .A(npu_inst_int_data_res_5__7__5_), .B(
        npu_inst_pe_1_5_7_add_79_carry_5_), .Z(npu_inst_pe_1_5_7_N78) );
  AND2_X1 npu_inst_pe_1_5_7_U122 ( .A1(npu_inst_pe_1_5_7_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_5__7__5_), .ZN(
        npu_inst_pe_1_5_7_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_5_7_U121 ( .A(npu_inst_int_data_res_5__7__6_), .B(
        npu_inst_pe_1_5_7_add_79_carry_6_), .Z(npu_inst_pe_1_5_7_N79) );
  AND2_X1 npu_inst_pe_1_5_7_U120 ( .A1(npu_inst_pe_1_5_7_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_5__7__6_), .ZN(
        npu_inst_pe_1_5_7_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_5_7_U119 ( .A(npu_inst_int_data_res_5__7__7_), .B(
        npu_inst_pe_1_5_7_add_79_carry_7_), .Z(npu_inst_pe_1_5_7_N80) );
  XNOR2_X1 npu_inst_pe_1_5_7_U118 ( .A(npu_inst_pe_1_5_7_sub_77_carry_2_), .B(
        npu_inst_int_data_res_5__7__2_), .ZN(npu_inst_pe_1_5_7_N67) );
  OR2_X1 npu_inst_pe_1_5_7_U117 ( .A1(npu_inst_int_data_res_5__7__2_), .A2(
        npu_inst_pe_1_5_7_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_5_7_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_5_7_U116 ( .A(npu_inst_pe_1_5_7_sub_77_carry_3_), .B(
        npu_inst_int_data_res_5__7__3_), .ZN(npu_inst_pe_1_5_7_N68) );
  OR2_X1 npu_inst_pe_1_5_7_U115 ( .A1(npu_inst_int_data_res_5__7__3_), .A2(
        npu_inst_pe_1_5_7_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_5_7_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_5_7_U114 ( .A(npu_inst_pe_1_5_7_sub_77_carry_4_), .B(
        npu_inst_int_data_res_5__7__4_), .ZN(npu_inst_pe_1_5_7_N69) );
  OR2_X1 npu_inst_pe_1_5_7_U113 ( .A1(npu_inst_int_data_res_5__7__4_), .A2(
        npu_inst_pe_1_5_7_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_5_7_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_5_7_U112 ( .A(npu_inst_pe_1_5_7_sub_77_carry_5_), .B(
        npu_inst_int_data_res_5__7__5_), .ZN(npu_inst_pe_1_5_7_N70) );
  OR2_X1 npu_inst_pe_1_5_7_U111 ( .A1(npu_inst_int_data_res_5__7__5_), .A2(
        npu_inst_pe_1_5_7_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_5_7_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_5_7_U110 ( .A(npu_inst_pe_1_5_7_sub_77_carry_6_), .B(
        npu_inst_int_data_res_5__7__6_), .ZN(npu_inst_pe_1_5_7_N71) );
  OR2_X1 npu_inst_pe_1_5_7_U109 ( .A1(npu_inst_int_data_res_5__7__6_), .A2(
        npu_inst_pe_1_5_7_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_5_7_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_5_7_U108 ( .A(npu_inst_int_data_res_5__7__7_), .B(
        npu_inst_pe_1_5_7_sub_77_carry_7_), .ZN(npu_inst_pe_1_5_7_N72) );
  INV_X1 npu_inst_pe_1_5_7_U107 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_5_7_n6)
         );
  INV_X1 npu_inst_pe_1_5_7_U106 ( .A(npu_inst_pe_1_5_7_n6), .ZN(
        npu_inst_pe_1_5_7_n5) );
  INV_X1 npu_inst_pe_1_5_7_U105 ( .A(npu_inst_n36), .ZN(npu_inst_pe_1_5_7_n2)
         );
  AOI22_X1 npu_inst_pe_1_5_7_U104 ( .A1(npu_inst_int_data_y_6__7__0_), .A2(
        npu_inst_pe_1_5_7_n58), .B1(npu_inst_pe_1_5_7_n118), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_5_7_n57) );
  INV_X1 npu_inst_pe_1_5_7_U103 ( .A(npu_inst_pe_1_5_7_n57), .ZN(
        npu_inst_pe_1_5_7_n107) );
  AOI22_X1 npu_inst_pe_1_5_7_U102 ( .A1(npu_inst_int_data_y_6__7__0_), .A2(
        npu_inst_pe_1_5_7_n54), .B1(npu_inst_pe_1_5_7_n117), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_5_7_n53) );
  INV_X1 npu_inst_pe_1_5_7_U99 ( .A(npu_inst_pe_1_5_7_n53), .ZN(
        npu_inst_pe_1_5_7_n108) );
  AOI22_X1 npu_inst_pe_1_5_7_U98 ( .A1(npu_inst_int_data_y_6__7__0_), .A2(
        npu_inst_pe_1_5_7_n50), .B1(npu_inst_pe_1_5_7_n116), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_5_7_n49) );
  INV_X1 npu_inst_pe_1_5_7_U97 ( .A(npu_inst_pe_1_5_7_n49), .ZN(
        npu_inst_pe_1_5_7_n109) );
  AOI22_X1 npu_inst_pe_1_5_7_U96 ( .A1(npu_inst_int_data_y_6__7__0_), .A2(
        npu_inst_pe_1_5_7_n46), .B1(npu_inst_pe_1_5_7_n115), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_5_7_n45) );
  INV_X1 npu_inst_pe_1_5_7_U95 ( .A(npu_inst_pe_1_5_7_n45), .ZN(
        npu_inst_pe_1_5_7_n110) );
  AOI22_X1 npu_inst_pe_1_5_7_U94 ( .A1(npu_inst_int_data_y_6__7__0_), .A2(
        npu_inst_pe_1_5_7_n42), .B1(npu_inst_pe_1_5_7_n114), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_5_7_n41) );
  INV_X1 npu_inst_pe_1_5_7_U93 ( .A(npu_inst_pe_1_5_7_n41), .ZN(
        npu_inst_pe_1_5_7_n111) );
  AOI22_X1 npu_inst_pe_1_5_7_U92 ( .A1(npu_inst_int_data_y_6__7__1_), .A2(
        npu_inst_pe_1_5_7_n58), .B1(npu_inst_pe_1_5_7_n118), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_5_7_n59) );
  INV_X1 npu_inst_pe_1_5_7_U91 ( .A(npu_inst_pe_1_5_7_n59), .ZN(
        npu_inst_pe_1_5_7_n101) );
  AOI22_X1 npu_inst_pe_1_5_7_U90 ( .A1(npu_inst_int_data_y_6__7__1_), .A2(
        npu_inst_pe_1_5_7_n54), .B1(npu_inst_pe_1_5_7_n117), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_5_7_n55) );
  INV_X1 npu_inst_pe_1_5_7_U89 ( .A(npu_inst_pe_1_5_7_n55), .ZN(
        npu_inst_pe_1_5_7_n102) );
  AOI22_X1 npu_inst_pe_1_5_7_U88 ( .A1(npu_inst_int_data_y_6__7__1_), .A2(
        npu_inst_pe_1_5_7_n50), .B1(npu_inst_pe_1_5_7_n116), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_5_7_n51) );
  INV_X1 npu_inst_pe_1_5_7_U87 ( .A(npu_inst_pe_1_5_7_n51), .ZN(
        npu_inst_pe_1_5_7_n103) );
  AOI22_X1 npu_inst_pe_1_5_7_U86 ( .A1(npu_inst_int_data_y_6__7__1_), .A2(
        npu_inst_pe_1_5_7_n46), .B1(npu_inst_pe_1_5_7_n115), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_5_7_n47) );
  INV_X1 npu_inst_pe_1_5_7_U85 ( .A(npu_inst_pe_1_5_7_n47), .ZN(
        npu_inst_pe_1_5_7_n104) );
  AOI22_X1 npu_inst_pe_1_5_7_U84 ( .A1(npu_inst_int_data_y_6__7__1_), .A2(
        npu_inst_pe_1_5_7_n42), .B1(npu_inst_pe_1_5_7_n114), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_5_7_n43) );
  INV_X1 npu_inst_pe_1_5_7_U83 ( .A(npu_inst_pe_1_5_7_n43), .ZN(
        npu_inst_pe_1_5_7_n105) );
  AOI22_X1 npu_inst_pe_1_5_7_U82 ( .A1(npu_inst_pe_1_5_7_n38), .A2(
        npu_inst_int_data_y_6__7__1_), .B1(npu_inst_pe_1_5_7_n113), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_5_7_n39) );
  INV_X1 npu_inst_pe_1_5_7_U81 ( .A(npu_inst_pe_1_5_7_n39), .ZN(
        npu_inst_pe_1_5_7_n106) );
  AND2_X1 npu_inst_pe_1_5_7_U80 ( .A1(npu_inst_pe_1_5_7_N93), .A2(npu_inst_n36), .ZN(npu_inst_int_data_y_5__7__0_) );
  AOI22_X1 npu_inst_pe_1_5_7_U79 ( .A1(npu_inst_pe_1_5_7_n38), .A2(
        npu_inst_int_data_y_6__7__0_), .B1(npu_inst_pe_1_5_7_n113), .B2(
        npu_inst_pe_1_5_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_5_7_n37) );
  INV_X1 npu_inst_pe_1_5_7_U78 ( .A(npu_inst_pe_1_5_7_n37), .ZN(
        npu_inst_pe_1_5_7_n112) );
  AND2_X1 npu_inst_pe_1_5_7_U77 ( .A1(npu_inst_n36), .A2(npu_inst_pe_1_5_7_N94), .ZN(npu_inst_int_data_y_5__7__1_) );
  AOI222_X1 npu_inst_pe_1_5_7_U76 ( .A1(npu_inst_int_data_res_6__7__0_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N73), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N65), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n84) );
  INV_X1 npu_inst_pe_1_5_7_U75 ( .A(npu_inst_pe_1_5_7_n84), .ZN(
        npu_inst_pe_1_5_7_n100) );
  AOI222_X1 npu_inst_pe_1_5_7_U74 ( .A1(npu_inst_pe_1_5_7_n1), .A2(
        npu_inst_int_data_res_6__7__7_), .B1(npu_inst_pe_1_5_7_N80), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N72), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n75) );
  INV_X1 npu_inst_pe_1_5_7_U73 ( .A(npu_inst_pe_1_5_7_n75), .ZN(
        npu_inst_pe_1_5_7_n32) );
  AOI222_X1 npu_inst_pe_1_5_7_U72 ( .A1(npu_inst_int_data_res_6__7__1_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N74), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N66), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n83) );
  INV_X1 npu_inst_pe_1_5_7_U71 ( .A(npu_inst_pe_1_5_7_n83), .ZN(
        npu_inst_pe_1_5_7_n99) );
  AOI222_X1 npu_inst_pe_1_5_7_U70 ( .A1(npu_inst_int_data_res_6__7__3_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N76), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N68), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n81) );
  INV_X1 npu_inst_pe_1_5_7_U69 ( .A(npu_inst_pe_1_5_7_n81), .ZN(
        npu_inst_pe_1_5_7_n36) );
  AOI222_X1 npu_inst_pe_1_5_7_U68 ( .A1(npu_inst_int_data_res_6__7__4_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N77), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N69), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n80) );
  INV_X1 npu_inst_pe_1_5_7_U67 ( .A(npu_inst_pe_1_5_7_n80), .ZN(
        npu_inst_pe_1_5_7_n35) );
  AOI222_X1 npu_inst_pe_1_5_7_U66 ( .A1(npu_inst_int_data_res_6__7__5_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N78), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N70), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n79) );
  INV_X1 npu_inst_pe_1_5_7_U65 ( .A(npu_inst_pe_1_5_7_n79), .ZN(
        npu_inst_pe_1_5_7_n34) );
  AOI222_X1 npu_inst_pe_1_5_7_U64 ( .A1(npu_inst_int_data_res_6__7__6_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N79), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N71), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n78) );
  INV_X1 npu_inst_pe_1_5_7_U63 ( .A(npu_inst_pe_1_5_7_n78), .ZN(
        npu_inst_pe_1_5_7_n33) );
  NOR3_X1 npu_inst_pe_1_5_7_U62 ( .A1(npu_inst_pe_1_5_7_n26), .A2(npu_inst_n36), .A3(npu_inst_int_ckg[16]), .ZN(npu_inst_pe_1_5_7_n85) );
  OR2_X1 npu_inst_pe_1_5_7_U61 ( .A1(npu_inst_pe_1_5_7_n85), .A2(
        npu_inst_pe_1_5_7_n1), .ZN(npu_inst_pe_1_5_7_N84) );
  AND2_X1 npu_inst_pe_1_5_7_U60 ( .A1(npu_inst_int_data_x_5__7__1_), .A2(
        npu_inst_pe_1_5_7_int_q_weight_1_), .ZN(npu_inst_pe_1_5_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_5_7_U59 ( .A1(npu_inst_int_data_x_5__7__0_), .A2(
        npu_inst_pe_1_5_7_int_q_weight_1_), .ZN(npu_inst_pe_1_5_7_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_5_7_U58 ( .A(npu_inst_pe_1_5_7_int_data_1_), .ZN(
        npu_inst_pe_1_5_7_n13) );
  NAND2_X1 npu_inst_pe_1_5_7_U57 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_5_7_n60), .ZN(npu_inst_pe_1_5_7_n74) );
  OAI21_X1 npu_inst_pe_1_5_7_U56 ( .B1(npu_inst_pe_1_5_7_n63), .B2(
        npu_inst_pe_1_5_7_n60), .A(npu_inst_pe_1_5_7_n74), .ZN(
        npu_inst_pe_1_5_7_n97) );
  NAND2_X1 npu_inst_pe_1_5_7_U55 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_5_7_n60), .ZN(npu_inst_pe_1_5_7_n73) );
  OAI21_X1 npu_inst_pe_1_5_7_U54 ( .B1(npu_inst_pe_1_5_7_n61), .B2(
        npu_inst_pe_1_5_7_n60), .A(npu_inst_pe_1_5_7_n73), .ZN(
        npu_inst_pe_1_5_7_n96) );
  NAND2_X1 npu_inst_pe_1_5_7_U53 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_5_7_n56), .ZN(npu_inst_pe_1_5_7_n72) );
  OAI21_X1 npu_inst_pe_1_5_7_U52 ( .B1(npu_inst_pe_1_5_7_n63), .B2(
        npu_inst_pe_1_5_7_n56), .A(npu_inst_pe_1_5_7_n72), .ZN(
        npu_inst_pe_1_5_7_n95) );
  NAND2_X1 npu_inst_pe_1_5_7_U51 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_5_7_n56), .ZN(npu_inst_pe_1_5_7_n71) );
  OAI21_X1 npu_inst_pe_1_5_7_U50 ( .B1(npu_inst_pe_1_5_7_n61), .B2(
        npu_inst_pe_1_5_7_n56), .A(npu_inst_pe_1_5_7_n71), .ZN(
        npu_inst_pe_1_5_7_n94) );
  NAND2_X1 npu_inst_pe_1_5_7_U49 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_5_7_n52), .ZN(npu_inst_pe_1_5_7_n70) );
  OAI21_X1 npu_inst_pe_1_5_7_U48 ( .B1(npu_inst_pe_1_5_7_n63), .B2(
        npu_inst_pe_1_5_7_n52), .A(npu_inst_pe_1_5_7_n70), .ZN(
        npu_inst_pe_1_5_7_n93) );
  NAND2_X1 npu_inst_pe_1_5_7_U47 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_5_7_n52), .ZN(npu_inst_pe_1_5_7_n69) );
  OAI21_X1 npu_inst_pe_1_5_7_U46 ( .B1(npu_inst_pe_1_5_7_n61), .B2(
        npu_inst_pe_1_5_7_n52), .A(npu_inst_pe_1_5_7_n69), .ZN(
        npu_inst_pe_1_5_7_n92) );
  NAND2_X1 npu_inst_pe_1_5_7_U45 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_5_7_n48), .ZN(npu_inst_pe_1_5_7_n68) );
  OAI21_X1 npu_inst_pe_1_5_7_U44 ( .B1(npu_inst_pe_1_5_7_n63), .B2(
        npu_inst_pe_1_5_7_n48), .A(npu_inst_pe_1_5_7_n68), .ZN(
        npu_inst_pe_1_5_7_n91) );
  NAND2_X1 npu_inst_pe_1_5_7_U43 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_5_7_n48), .ZN(npu_inst_pe_1_5_7_n67) );
  OAI21_X1 npu_inst_pe_1_5_7_U42 ( .B1(npu_inst_pe_1_5_7_n61), .B2(
        npu_inst_pe_1_5_7_n48), .A(npu_inst_pe_1_5_7_n67), .ZN(
        npu_inst_pe_1_5_7_n90) );
  NAND2_X1 npu_inst_pe_1_5_7_U41 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_5_7_n44), .ZN(npu_inst_pe_1_5_7_n66) );
  OAI21_X1 npu_inst_pe_1_5_7_U40 ( .B1(npu_inst_pe_1_5_7_n63), .B2(
        npu_inst_pe_1_5_7_n44), .A(npu_inst_pe_1_5_7_n66), .ZN(
        npu_inst_pe_1_5_7_n89) );
  NAND2_X1 npu_inst_pe_1_5_7_U39 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_5_7_n44), .ZN(npu_inst_pe_1_5_7_n65) );
  OAI21_X1 npu_inst_pe_1_5_7_U38 ( .B1(npu_inst_pe_1_5_7_n61), .B2(
        npu_inst_pe_1_5_7_n44), .A(npu_inst_pe_1_5_7_n65), .ZN(
        npu_inst_pe_1_5_7_n88) );
  NAND2_X1 npu_inst_pe_1_5_7_U37 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_5_7_n40), .ZN(npu_inst_pe_1_5_7_n64) );
  OAI21_X1 npu_inst_pe_1_5_7_U36 ( .B1(npu_inst_pe_1_5_7_n63), .B2(
        npu_inst_pe_1_5_7_n40), .A(npu_inst_pe_1_5_7_n64), .ZN(
        npu_inst_pe_1_5_7_n87) );
  NAND2_X1 npu_inst_pe_1_5_7_U35 ( .A1(npu_inst_pe_1_5_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_5_7_n40), .ZN(npu_inst_pe_1_5_7_n62) );
  OAI21_X1 npu_inst_pe_1_5_7_U34 ( .B1(npu_inst_pe_1_5_7_n61), .B2(
        npu_inst_pe_1_5_7_n40), .A(npu_inst_pe_1_5_7_n62), .ZN(
        npu_inst_pe_1_5_7_n86) );
  AOI222_X1 npu_inst_pe_1_5_7_U33 ( .A1(npu_inst_int_data_res_6__7__2_), .A2(
        npu_inst_pe_1_5_7_n1), .B1(npu_inst_pe_1_5_7_N75), .B2(
        npu_inst_pe_1_5_7_n76), .C1(npu_inst_pe_1_5_7_N67), .C2(
        npu_inst_pe_1_5_7_n77), .ZN(npu_inst_pe_1_5_7_n82) );
  INV_X1 npu_inst_pe_1_5_7_U32 ( .A(npu_inst_pe_1_5_7_n82), .ZN(
        npu_inst_pe_1_5_7_n98) );
  INV_X1 npu_inst_pe_1_5_7_U31 ( .A(npu_inst_pe_1_5_7_int_data_0_), .ZN(
        npu_inst_pe_1_5_7_n12) );
  INV_X1 npu_inst_pe_1_5_7_U30 ( .A(npu_inst_n50), .ZN(npu_inst_pe_1_5_7_n4)
         );
  AOI22_X1 npu_inst_pe_1_5_7_U29 ( .A1(npu_inst_n36), .A2(
        npu_inst_int_data_y_6__7__1_), .B1(npu_inst_pe_1_5_7_n2), .B2(
        int_i_data_h_npu[5]), .ZN(npu_inst_pe_1_5_7_n63) );
  AOI22_X1 npu_inst_pe_1_5_7_U28 ( .A1(npu_inst_n36), .A2(
        npu_inst_int_data_y_6__7__0_), .B1(npu_inst_pe_1_5_7_n2), .B2(
        int_i_data_h_npu[4]), .ZN(npu_inst_pe_1_5_7_n61) );
  OR3_X1 npu_inst_pe_1_5_7_U27 ( .A1(npu_inst_pe_1_5_7_n5), .A2(
        npu_inst_pe_1_5_7_n7), .A3(npu_inst_pe_1_5_7_n4), .ZN(
        npu_inst_pe_1_5_7_n56) );
  OR3_X1 npu_inst_pe_1_5_7_U26 ( .A1(npu_inst_pe_1_5_7_n4), .A2(
        npu_inst_pe_1_5_7_n7), .A3(npu_inst_pe_1_5_7_n6), .ZN(
        npu_inst_pe_1_5_7_n48) );
  INV_X1 npu_inst_pe_1_5_7_U25 ( .A(npu_inst_pe_1_5_7_n4), .ZN(
        npu_inst_pe_1_5_7_n3) );
  OR3_X1 npu_inst_pe_1_5_7_U24 ( .A1(npu_inst_pe_1_5_7_n3), .A2(
        npu_inst_pe_1_5_7_n7), .A3(npu_inst_pe_1_5_7_n6), .ZN(
        npu_inst_pe_1_5_7_n52) );
  OR3_X1 npu_inst_pe_1_5_7_U23 ( .A1(npu_inst_pe_1_5_7_n5), .A2(
        npu_inst_pe_1_5_7_n7), .A3(npu_inst_pe_1_5_7_n3), .ZN(
        npu_inst_pe_1_5_7_n60) );
  BUF_X1 npu_inst_pe_1_5_7_U22 ( .A(npu_inst_n16), .Z(npu_inst_pe_1_5_7_n1) );
  NOR2_X1 npu_inst_pe_1_5_7_U21 ( .A1(npu_inst_pe_1_5_7_n60), .A2(
        npu_inst_pe_1_5_7_n2), .ZN(npu_inst_pe_1_5_7_n58) );
  NOR2_X1 npu_inst_pe_1_5_7_U20 ( .A1(npu_inst_pe_1_5_7_n56), .A2(
        npu_inst_pe_1_5_7_n2), .ZN(npu_inst_pe_1_5_7_n54) );
  NOR2_X1 npu_inst_pe_1_5_7_U19 ( .A1(npu_inst_pe_1_5_7_n52), .A2(
        npu_inst_pe_1_5_7_n2), .ZN(npu_inst_pe_1_5_7_n50) );
  NOR2_X1 npu_inst_pe_1_5_7_U18 ( .A1(npu_inst_pe_1_5_7_n48), .A2(
        npu_inst_pe_1_5_7_n2), .ZN(npu_inst_pe_1_5_7_n46) );
  NOR2_X1 npu_inst_pe_1_5_7_U17 ( .A1(npu_inst_pe_1_5_7_n40), .A2(
        npu_inst_pe_1_5_7_n2), .ZN(npu_inst_pe_1_5_7_n38) );
  NOR2_X1 npu_inst_pe_1_5_7_U16 ( .A1(npu_inst_pe_1_5_7_n44), .A2(
        npu_inst_pe_1_5_7_n2), .ZN(npu_inst_pe_1_5_7_n42) );
  BUF_X1 npu_inst_pe_1_5_7_U15 ( .A(npu_inst_n78), .Z(npu_inst_pe_1_5_7_n7) );
  INV_X1 npu_inst_pe_1_5_7_U14 ( .A(npu_inst_n105), .ZN(npu_inst_pe_1_5_7_n11)
         );
  INV_X1 npu_inst_pe_1_5_7_U13 ( .A(npu_inst_pe_1_5_7_n38), .ZN(
        npu_inst_pe_1_5_7_n113) );
  INV_X1 npu_inst_pe_1_5_7_U12 ( .A(npu_inst_pe_1_5_7_n58), .ZN(
        npu_inst_pe_1_5_7_n118) );
  INV_X1 npu_inst_pe_1_5_7_U11 ( .A(npu_inst_pe_1_5_7_n54), .ZN(
        npu_inst_pe_1_5_7_n117) );
  INV_X1 npu_inst_pe_1_5_7_U10 ( .A(npu_inst_pe_1_5_7_n50), .ZN(
        npu_inst_pe_1_5_7_n116) );
  INV_X1 npu_inst_pe_1_5_7_U9 ( .A(npu_inst_pe_1_5_7_n46), .ZN(
        npu_inst_pe_1_5_7_n115) );
  INV_X1 npu_inst_pe_1_5_7_U8 ( .A(npu_inst_pe_1_5_7_n42), .ZN(
        npu_inst_pe_1_5_7_n114) );
  BUF_X1 npu_inst_pe_1_5_7_U7 ( .A(npu_inst_pe_1_5_7_n11), .Z(
        npu_inst_pe_1_5_7_n10) );
  BUF_X1 npu_inst_pe_1_5_7_U6 ( .A(npu_inst_pe_1_5_7_n11), .Z(
        npu_inst_pe_1_5_7_n9) );
  BUF_X1 npu_inst_pe_1_5_7_U5 ( .A(npu_inst_pe_1_5_7_n11), .Z(
        npu_inst_pe_1_5_7_n8) );
  NOR2_X1 npu_inst_pe_1_5_7_U4 ( .A1(npu_inst_pe_1_5_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_5_7_n1), .ZN(npu_inst_pe_1_5_7_n76) );
  NOR2_X1 npu_inst_pe_1_5_7_U3 ( .A1(npu_inst_pe_1_5_7_n27), .A2(
        npu_inst_pe_1_5_7_n1), .ZN(npu_inst_pe_1_5_7_n77) );
  FA_X1 npu_inst_pe_1_5_7_sub_77_U2_1 ( .A(npu_inst_int_data_res_5__7__1_), 
        .B(npu_inst_pe_1_5_7_n13), .CI(npu_inst_pe_1_5_7_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_5_7_sub_77_carry_2_), .S(npu_inst_pe_1_5_7_N66) );
  FA_X1 npu_inst_pe_1_5_7_add_79_U1_1 ( .A(npu_inst_int_data_res_5__7__1_), 
        .B(npu_inst_pe_1_5_7_int_data_1_), .CI(
        npu_inst_pe_1_5_7_add_79_carry_1_), .CO(
        npu_inst_pe_1_5_7_add_79_carry_2_), .S(npu_inst_pe_1_5_7_N74) );
  NAND3_X1 npu_inst_pe_1_5_7_U101 ( .A1(npu_inst_pe_1_5_7_n4), .A2(
        npu_inst_pe_1_5_7_n6), .A3(npu_inst_pe_1_5_7_n7), .ZN(
        npu_inst_pe_1_5_7_n44) );
  NAND3_X1 npu_inst_pe_1_5_7_U100 ( .A1(npu_inst_pe_1_5_7_n3), .A2(
        npu_inst_pe_1_5_7_n6), .A3(npu_inst_pe_1_5_7_n7), .ZN(
        npu_inst_pe_1_5_7_n40) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_5_7_n33), .CK(
        npu_inst_pe_1_5_7_net3397), .RN(npu_inst_pe_1_5_7_n8), .Q(
        npu_inst_int_data_res_5__7__6_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_5_7_n34), .CK(
        npu_inst_pe_1_5_7_net3397), .RN(npu_inst_pe_1_5_7_n8), .Q(
        npu_inst_int_data_res_5__7__5_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_5_7_n35), .CK(
        npu_inst_pe_1_5_7_net3397), .RN(npu_inst_pe_1_5_7_n8), .Q(
        npu_inst_int_data_res_5__7__4_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_5_7_n36), .CK(
        npu_inst_pe_1_5_7_net3397), .RN(npu_inst_pe_1_5_7_n8), .Q(
        npu_inst_int_data_res_5__7__3_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_5_7_n98), .CK(
        npu_inst_pe_1_5_7_net3397), .RN(npu_inst_pe_1_5_7_n8), .Q(
        npu_inst_int_data_res_5__7__2_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_5_7_n99), .CK(
        npu_inst_pe_1_5_7_net3397), .RN(npu_inst_pe_1_5_7_n8), .Q(
        npu_inst_int_data_res_5__7__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_5_7_n32), .CK(
        npu_inst_pe_1_5_7_net3397), .RN(npu_inst_pe_1_5_7_n8), .Q(
        npu_inst_int_data_res_5__7__7_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_5_7_n100), 
        .CK(npu_inst_pe_1_5_7_net3397), .RN(npu_inst_pe_1_5_7_n8), .Q(
        npu_inst_int_data_res_5__7__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_weight_reg_0_ ( .D(npu_inst_n91), .CK(
        npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n8), .Q(
        npu_inst_pe_1_5_7_int_q_weight_0_), .QN(npu_inst_pe_1_5_7_n27) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_weight_reg_1_ ( .D(npu_inst_n97), .CK(
        npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n8), .Q(
        npu_inst_pe_1_5_7_int_q_weight_1_), .QN(npu_inst_pe_1_5_7_n26) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_5_7_n112), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n8), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_5_7_n106), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n8), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_5_7_n111), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_5_7_n105), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_5_7_n110), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_5_7_n104), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_5_7_n109), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_5_7_n103), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_5_7_n108), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_5_7_n102), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_5_7_n107), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_5_7_n101), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_5_7_n86), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_5_7_n87), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n9), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_5_7_n88), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_5_7_n89), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_5_7_n90), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_5_7_n91), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_5_7_n92), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_5_7_n93), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_5_7_n94), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_5_7_n95), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_5_7_n96), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_5_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_5_7_n97), 
        .CK(npu_inst_pe_1_5_7_net3403), .RN(npu_inst_pe_1_5_7_n10), .Q(
        npu_inst_pe_1_5_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_5_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_5_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_5_7_net3397) );
  CLKGATETST_X1 npu_inst_pe_1_5_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n44), .SE(1'b0), .GCK(npu_inst_pe_1_5_7_net3403) );
  MUX2_X1 npu_inst_pe_1_6_0_U153 ( .A(npu_inst_pe_1_6_0_n31), .B(
        npu_inst_pe_1_6_0_n28), .S(npu_inst_pe_1_6_0_n7), .Z(
        npu_inst_pe_1_6_0_N93) );
  MUX2_X1 npu_inst_pe_1_6_0_U152 ( .A(npu_inst_pe_1_6_0_n30), .B(
        npu_inst_pe_1_6_0_n29), .S(npu_inst_pe_1_6_0_n5), .Z(
        npu_inst_pe_1_6_0_n31) );
  MUX2_X1 npu_inst_pe_1_6_0_U151 ( .A(npu_inst_pe_1_6_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_0_n3), .Z(
        npu_inst_pe_1_6_0_n30) );
  MUX2_X1 npu_inst_pe_1_6_0_U150 ( .A(npu_inst_pe_1_6_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_0_n3), .Z(
        npu_inst_pe_1_6_0_n29) );
  MUX2_X1 npu_inst_pe_1_6_0_U149 ( .A(npu_inst_pe_1_6_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_0_n3), .Z(
        npu_inst_pe_1_6_0_n28) );
  MUX2_X1 npu_inst_pe_1_6_0_U148 ( .A(npu_inst_pe_1_6_0_n25), .B(
        npu_inst_pe_1_6_0_n22), .S(npu_inst_pe_1_6_0_n7), .Z(
        npu_inst_pe_1_6_0_N94) );
  MUX2_X1 npu_inst_pe_1_6_0_U147 ( .A(npu_inst_pe_1_6_0_n24), .B(
        npu_inst_pe_1_6_0_n23), .S(npu_inst_pe_1_6_0_n5), .Z(
        npu_inst_pe_1_6_0_n25) );
  MUX2_X1 npu_inst_pe_1_6_0_U146 ( .A(npu_inst_pe_1_6_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_0_n3), .Z(
        npu_inst_pe_1_6_0_n24) );
  MUX2_X1 npu_inst_pe_1_6_0_U145 ( .A(npu_inst_pe_1_6_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_0_n3), .Z(
        npu_inst_pe_1_6_0_n23) );
  MUX2_X1 npu_inst_pe_1_6_0_U144 ( .A(npu_inst_pe_1_6_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_0_n3), .Z(
        npu_inst_pe_1_6_0_n22) );
  MUX2_X1 npu_inst_pe_1_6_0_U143 ( .A(npu_inst_pe_1_6_0_n21), .B(
        npu_inst_pe_1_6_0_n18), .S(npu_inst_pe_1_6_0_n7), .Z(
        npu_inst_pe_1_6_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_6_0_U142 ( .A(npu_inst_pe_1_6_0_n20), .B(
        npu_inst_pe_1_6_0_n19), .S(npu_inst_pe_1_6_0_n5), .Z(
        npu_inst_pe_1_6_0_n21) );
  MUX2_X1 npu_inst_pe_1_6_0_U141 ( .A(npu_inst_pe_1_6_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_0_n3), .Z(
        npu_inst_pe_1_6_0_n20) );
  MUX2_X1 npu_inst_pe_1_6_0_U140 ( .A(npu_inst_pe_1_6_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_0_n3), .Z(
        npu_inst_pe_1_6_0_n19) );
  MUX2_X1 npu_inst_pe_1_6_0_U139 ( .A(npu_inst_pe_1_6_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_0_n3), .Z(
        npu_inst_pe_1_6_0_n18) );
  MUX2_X1 npu_inst_pe_1_6_0_U138 ( .A(npu_inst_pe_1_6_0_n17), .B(
        npu_inst_pe_1_6_0_n14), .S(npu_inst_pe_1_6_0_n7), .Z(
        npu_inst_pe_1_6_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_6_0_U137 ( .A(npu_inst_pe_1_6_0_n16), .B(
        npu_inst_pe_1_6_0_n15), .S(npu_inst_pe_1_6_0_n5), .Z(
        npu_inst_pe_1_6_0_n17) );
  MUX2_X1 npu_inst_pe_1_6_0_U136 ( .A(npu_inst_pe_1_6_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_0_n3), .Z(
        npu_inst_pe_1_6_0_n16) );
  MUX2_X1 npu_inst_pe_1_6_0_U135 ( .A(npu_inst_pe_1_6_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_0_n3), .Z(
        npu_inst_pe_1_6_0_n15) );
  MUX2_X1 npu_inst_pe_1_6_0_U134 ( .A(npu_inst_pe_1_6_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_0_n3), .Z(
        npu_inst_pe_1_6_0_n14) );
  XOR2_X1 npu_inst_pe_1_6_0_U133 ( .A(npu_inst_pe_1_6_0_int_data_0_), .B(
        npu_inst_int_data_res_6__0__0_), .Z(npu_inst_pe_1_6_0_N73) );
  AND2_X1 npu_inst_pe_1_6_0_U132 ( .A1(npu_inst_int_data_res_6__0__0_), .A2(
        npu_inst_pe_1_6_0_int_data_0_), .ZN(npu_inst_pe_1_6_0_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_0_U131 ( .A(npu_inst_int_data_res_6__0__0_), .B(
        npu_inst_pe_1_6_0_n12), .ZN(npu_inst_pe_1_6_0_N65) );
  OR2_X1 npu_inst_pe_1_6_0_U130 ( .A1(npu_inst_pe_1_6_0_n12), .A2(
        npu_inst_int_data_res_6__0__0_), .ZN(npu_inst_pe_1_6_0_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_0_U129 ( .A(npu_inst_int_data_res_6__0__2_), .B(
        npu_inst_pe_1_6_0_add_79_carry_2_), .Z(npu_inst_pe_1_6_0_N75) );
  AND2_X1 npu_inst_pe_1_6_0_U128 ( .A1(npu_inst_pe_1_6_0_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_6__0__2_), .ZN(
        npu_inst_pe_1_6_0_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_0_U127 ( .A(npu_inst_int_data_res_6__0__3_), .B(
        npu_inst_pe_1_6_0_add_79_carry_3_), .Z(npu_inst_pe_1_6_0_N76) );
  AND2_X1 npu_inst_pe_1_6_0_U126 ( .A1(npu_inst_pe_1_6_0_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_6__0__3_), .ZN(
        npu_inst_pe_1_6_0_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_0_U125 ( .A(npu_inst_int_data_res_6__0__4_), .B(
        npu_inst_pe_1_6_0_add_79_carry_4_), .Z(npu_inst_pe_1_6_0_N77) );
  AND2_X1 npu_inst_pe_1_6_0_U124 ( .A1(npu_inst_pe_1_6_0_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_6__0__4_), .ZN(
        npu_inst_pe_1_6_0_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_0_U123 ( .A(npu_inst_int_data_res_6__0__5_), .B(
        npu_inst_pe_1_6_0_add_79_carry_5_), .Z(npu_inst_pe_1_6_0_N78) );
  AND2_X1 npu_inst_pe_1_6_0_U122 ( .A1(npu_inst_pe_1_6_0_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_6__0__5_), .ZN(
        npu_inst_pe_1_6_0_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_0_U121 ( .A(npu_inst_int_data_res_6__0__6_), .B(
        npu_inst_pe_1_6_0_add_79_carry_6_), .Z(npu_inst_pe_1_6_0_N79) );
  AND2_X1 npu_inst_pe_1_6_0_U120 ( .A1(npu_inst_pe_1_6_0_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_6__0__6_), .ZN(
        npu_inst_pe_1_6_0_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_0_U119 ( .A(npu_inst_int_data_res_6__0__7_), .B(
        npu_inst_pe_1_6_0_add_79_carry_7_), .Z(npu_inst_pe_1_6_0_N80) );
  XNOR2_X1 npu_inst_pe_1_6_0_U118 ( .A(npu_inst_pe_1_6_0_sub_77_carry_2_), .B(
        npu_inst_int_data_res_6__0__2_), .ZN(npu_inst_pe_1_6_0_N67) );
  OR2_X1 npu_inst_pe_1_6_0_U117 ( .A1(npu_inst_int_data_res_6__0__2_), .A2(
        npu_inst_pe_1_6_0_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_6_0_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_0_U116 ( .A(npu_inst_pe_1_6_0_sub_77_carry_3_), .B(
        npu_inst_int_data_res_6__0__3_), .ZN(npu_inst_pe_1_6_0_N68) );
  OR2_X1 npu_inst_pe_1_6_0_U115 ( .A1(npu_inst_int_data_res_6__0__3_), .A2(
        npu_inst_pe_1_6_0_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_6_0_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_0_U114 ( .A(npu_inst_pe_1_6_0_sub_77_carry_4_), .B(
        npu_inst_int_data_res_6__0__4_), .ZN(npu_inst_pe_1_6_0_N69) );
  OR2_X1 npu_inst_pe_1_6_0_U113 ( .A1(npu_inst_int_data_res_6__0__4_), .A2(
        npu_inst_pe_1_6_0_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_6_0_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_0_U112 ( .A(npu_inst_pe_1_6_0_sub_77_carry_5_), .B(
        npu_inst_int_data_res_6__0__5_), .ZN(npu_inst_pe_1_6_0_N70) );
  OR2_X1 npu_inst_pe_1_6_0_U111 ( .A1(npu_inst_int_data_res_6__0__5_), .A2(
        npu_inst_pe_1_6_0_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_6_0_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_0_U110 ( .A(npu_inst_pe_1_6_0_sub_77_carry_6_), .B(
        npu_inst_int_data_res_6__0__6_), .ZN(npu_inst_pe_1_6_0_N71) );
  OR2_X1 npu_inst_pe_1_6_0_U109 ( .A1(npu_inst_int_data_res_6__0__6_), .A2(
        npu_inst_pe_1_6_0_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_6_0_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_0_U108 ( .A(npu_inst_int_data_res_6__0__7_), .B(
        npu_inst_pe_1_6_0_sub_77_carry_7_), .ZN(npu_inst_pe_1_6_0_N72) );
  INV_X1 npu_inst_pe_1_6_0_U107 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_6_0_n6)
         );
  INV_X1 npu_inst_pe_1_6_0_U106 ( .A(npu_inst_pe_1_6_0_n6), .ZN(
        npu_inst_pe_1_6_0_n5) );
  INV_X1 npu_inst_pe_1_6_0_U105 ( .A(npu_inst_n36), .ZN(npu_inst_pe_1_6_0_n2)
         );
  AOI22_X1 npu_inst_pe_1_6_0_U104 ( .A1(npu_inst_int_data_y_7__0__0_), .A2(
        npu_inst_pe_1_6_0_n58), .B1(npu_inst_pe_1_6_0_n118), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_0_n57) );
  INV_X1 npu_inst_pe_1_6_0_U103 ( .A(npu_inst_pe_1_6_0_n57), .ZN(
        npu_inst_pe_1_6_0_n107) );
  AOI22_X1 npu_inst_pe_1_6_0_U102 ( .A1(npu_inst_int_data_y_7__0__0_), .A2(
        npu_inst_pe_1_6_0_n54), .B1(npu_inst_pe_1_6_0_n117), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_0_n53) );
  INV_X1 npu_inst_pe_1_6_0_U99 ( .A(npu_inst_pe_1_6_0_n53), .ZN(
        npu_inst_pe_1_6_0_n108) );
  AOI22_X1 npu_inst_pe_1_6_0_U98 ( .A1(npu_inst_int_data_y_7__0__0_), .A2(
        npu_inst_pe_1_6_0_n50), .B1(npu_inst_pe_1_6_0_n116), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_0_n49) );
  INV_X1 npu_inst_pe_1_6_0_U97 ( .A(npu_inst_pe_1_6_0_n49), .ZN(
        npu_inst_pe_1_6_0_n109) );
  AOI22_X1 npu_inst_pe_1_6_0_U96 ( .A1(npu_inst_int_data_y_7__0__0_), .A2(
        npu_inst_pe_1_6_0_n46), .B1(npu_inst_pe_1_6_0_n115), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_0_n45) );
  INV_X1 npu_inst_pe_1_6_0_U95 ( .A(npu_inst_pe_1_6_0_n45), .ZN(
        npu_inst_pe_1_6_0_n110) );
  AOI22_X1 npu_inst_pe_1_6_0_U94 ( .A1(npu_inst_int_data_y_7__0__0_), .A2(
        npu_inst_pe_1_6_0_n42), .B1(npu_inst_pe_1_6_0_n114), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_0_n41) );
  INV_X1 npu_inst_pe_1_6_0_U93 ( .A(npu_inst_pe_1_6_0_n41), .ZN(
        npu_inst_pe_1_6_0_n111) );
  AOI22_X1 npu_inst_pe_1_6_0_U92 ( .A1(npu_inst_int_data_y_7__0__1_), .A2(
        npu_inst_pe_1_6_0_n58), .B1(npu_inst_pe_1_6_0_n118), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_0_n59) );
  INV_X1 npu_inst_pe_1_6_0_U91 ( .A(npu_inst_pe_1_6_0_n59), .ZN(
        npu_inst_pe_1_6_0_n101) );
  AOI22_X1 npu_inst_pe_1_6_0_U90 ( .A1(npu_inst_int_data_y_7__0__1_), .A2(
        npu_inst_pe_1_6_0_n54), .B1(npu_inst_pe_1_6_0_n117), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_0_n55) );
  INV_X1 npu_inst_pe_1_6_0_U89 ( .A(npu_inst_pe_1_6_0_n55), .ZN(
        npu_inst_pe_1_6_0_n102) );
  AOI22_X1 npu_inst_pe_1_6_0_U88 ( .A1(npu_inst_int_data_y_7__0__1_), .A2(
        npu_inst_pe_1_6_0_n50), .B1(npu_inst_pe_1_6_0_n116), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_0_n51) );
  INV_X1 npu_inst_pe_1_6_0_U87 ( .A(npu_inst_pe_1_6_0_n51), .ZN(
        npu_inst_pe_1_6_0_n103) );
  AOI22_X1 npu_inst_pe_1_6_0_U86 ( .A1(npu_inst_int_data_y_7__0__1_), .A2(
        npu_inst_pe_1_6_0_n46), .B1(npu_inst_pe_1_6_0_n115), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_0_n47) );
  INV_X1 npu_inst_pe_1_6_0_U85 ( .A(npu_inst_pe_1_6_0_n47), .ZN(
        npu_inst_pe_1_6_0_n104) );
  AOI22_X1 npu_inst_pe_1_6_0_U84 ( .A1(npu_inst_int_data_y_7__0__1_), .A2(
        npu_inst_pe_1_6_0_n42), .B1(npu_inst_pe_1_6_0_n114), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_0_n43) );
  INV_X1 npu_inst_pe_1_6_0_U83 ( .A(npu_inst_pe_1_6_0_n43), .ZN(
        npu_inst_pe_1_6_0_n105) );
  AOI22_X1 npu_inst_pe_1_6_0_U82 ( .A1(npu_inst_pe_1_6_0_n38), .A2(
        npu_inst_int_data_y_7__0__1_), .B1(npu_inst_pe_1_6_0_n113), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_0_n39) );
  INV_X1 npu_inst_pe_1_6_0_U81 ( .A(npu_inst_pe_1_6_0_n39), .ZN(
        npu_inst_pe_1_6_0_n106) );
  AND2_X1 npu_inst_pe_1_6_0_U80 ( .A1(npu_inst_pe_1_6_0_N93), .A2(npu_inst_n36), .ZN(npu_inst_int_data_y_6__0__0_) );
  NAND2_X1 npu_inst_pe_1_6_0_U79 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_0_n60), .ZN(npu_inst_pe_1_6_0_n74) );
  OAI21_X1 npu_inst_pe_1_6_0_U78 ( .B1(npu_inst_pe_1_6_0_n63), .B2(
        npu_inst_pe_1_6_0_n60), .A(npu_inst_pe_1_6_0_n74), .ZN(
        npu_inst_pe_1_6_0_n97) );
  NAND2_X1 npu_inst_pe_1_6_0_U77 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_0_n60), .ZN(npu_inst_pe_1_6_0_n73) );
  OAI21_X1 npu_inst_pe_1_6_0_U76 ( .B1(npu_inst_pe_1_6_0_n61), .B2(
        npu_inst_pe_1_6_0_n60), .A(npu_inst_pe_1_6_0_n73), .ZN(
        npu_inst_pe_1_6_0_n96) );
  NAND2_X1 npu_inst_pe_1_6_0_U75 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_0_n56), .ZN(npu_inst_pe_1_6_0_n72) );
  OAI21_X1 npu_inst_pe_1_6_0_U74 ( .B1(npu_inst_pe_1_6_0_n63), .B2(
        npu_inst_pe_1_6_0_n56), .A(npu_inst_pe_1_6_0_n72), .ZN(
        npu_inst_pe_1_6_0_n95) );
  NAND2_X1 npu_inst_pe_1_6_0_U73 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_0_n56), .ZN(npu_inst_pe_1_6_0_n71) );
  OAI21_X1 npu_inst_pe_1_6_0_U72 ( .B1(npu_inst_pe_1_6_0_n61), .B2(
        npu_inst_pe_1_6_0_n56), .A(npu_inst_pe_1_6_0_n71), .ZN(
        npu_inst_pe_1_6_0_n94) );
  NAND2_X1 npu_inst_pe_1_6_0_U71 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_0_n52), .ZN(npu_inst_pe_1_6_0_n70) );
  OAI21_X1 npu_inst_pe_1_6_0_U70 ( .B1(npu_inst_pe_1_6_0_n63), .B2(
        npu_inst_pe_1_6_0_n52), .A(npu_inst_pe_1_6_0_n70), .ZN(
        npu_inst_pe_1_6_0_n93) );
  NAND2_X1 npu_inst_pe_1_6_0_U69 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_0_n52), .ZN(npu_inst_pe_1_6_0_n69) );
  OAI21_X1 npu_inst_pe_1_6_0_U68 ( .B1(npu_inst_pe_1_6_0_n61), .B2(
        npu_inst_pe_1_6_0_n52), .A(npu_inst_pe_1_6_0_n69), .ZN(
        npu_inst_pe_1_6_0_n92) );
  NAND2_X1 npu_inst_pe_1_6_0_U67 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_0_n48), .ZN(npu_inst_pe_1_6_0_n68) );
  OAI21_X1 npu_inst_pe_1_6_0_U66 ( .B1(npu_inst_pe_1_6_0_n63), .B2(
        npu_inst_pe_1_6_0_n48), .A(npu_inst_pe_1_6_0_n68), .ZN(
        npu_inst_pe_1_6_0_n91) );
  NAND2_X1 npu_inst_pe_1_6_0_U65 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_0_n48), .ZN(npu_inst_pe_1_6_0_n67) );
  OAI21_X1 npu_inst_pe_1_6_0_U64 ( .B1(npu_inst_pe_1_6_0_n61), .B2(
        npu_inst_pe_1_6_0_n48), .A(npu_inst_pe_1_6_0_n67), .ZN(
        npu_inst_pe_1_6_0_n90) );
  NAND2_X1 npu_inst_pe_1_6_0_U63 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_0_n44), .ZN(npu_inst_pe_1_6_0_n66) );
  OAI21_X1 npu_inst_pe_1_6_0_U62 ( .B1(npu_inst_pe_1_6_0_n63), .B2(
        npu_inst_pe_1_6_0_n44), .A(npu_inst_pe_1_6_0_n66), .ZN(
        npu_inst_pe_1_6_0_n89) );
  NAND2_X1 npu_inst_pe_1_6_0_U61 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_0_n44), .ZN(npu_inst_pe_1_6_0_n65) );
  OAI21_X1 npu_inst_pe_1_6_0_U60 ( .B1(npu_inst_pe_1_6_0_n61), .B2(
        npu_inst_pe_1_6_0_n44), .A(npu_inst_pe_1_6_0_n65), .ZN(
        npu_inst_pe_1_6_0_n88) );
  NAND2_X1 npu_inst_pe_1_6_0_U59 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_0_n40), .ZN(npu_inst_pe_1_6_0_n64) );
  OAI21_X1 npu_inst_pe_1_6_0_U58 ( .B1(npu_inst_pe_1_6_0_n63), .B2(
        npu_inst_pe_1_6_0_n40), .A(npu_inst_pe_1_6_0_n64), .ZN(
        npu_inst_pe_1_6_0_n87) );
  NAND2_X1 npu_inst_pe_1_6_0_U57 ( .A1(npu_inst_pe_1_6_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_0_n40), .ZN(npu_inst_pe_1_6_0_n62) );
  OAI21_X1 npu_inst_pe_1_6_0_U56 ( .B1(npu_inst_pe_1_6_0_n61), .B2(
        npu_inst_pe_1_6_0_n40), .A(npu_inst_pe_1_6_0_n62), .ZN(
        npu_inst_pe_1_6_0_n86) );
  AOI22_X1 npu_inst_pe_1_6_0_U55 ( .A1(npu_inst_pe_1_6_0_n38), .A2(
        npu_inst_int_data_y_7__0__0_), .B1(npu_inst_pe_1_6_0_n113), .B2(
        npu_inst_pe_1_6_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_0_n37) );
  INV_X1 npu_inst_pe_1_6_0_U54 ( .A(npu_inst_pe_1_6_0_n37), .ZN(
        npu_inst_pe_1_6_0_n112) );
  AND2_X1 npu_inst_pe_1_6_0_U53 ( .A1(npu_inst_n36), .A2(npu_inst_pe_1_6_0_N94), .ZN(npu_inst_int_data_y_6__0__1_) );
  AOI222_X1 npu_inst_pe_1_6_0_U52 ( .A1(npu_inst_int_data_res_7__0__0_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N73), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N65), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n84) );
  INV_X1 npu_inst_pe_1_6_0_U51 ( .A(npu_inst_pe_1_6_0_n84), .ZN(
        npu_inst_pe_1_6_0_n100) );
  AOI222_X1 npu_inst_pe_1_6_0_U50 ( .A1(npu_inst_pe_1_6_0_n1), .A2(
        npu_inst_int_data_res_7__0__7_), .B1(npu_inst_pe_1_6_0_N80), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N72), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n75) );
  INV_X1 npu_inst_pe_1_6_0_U49 ( .A(npu_inst_pe_1_6_0_n75), .ZN(
        npu_inst_pe_1_6_0_n32) );
  AOI222_X1 npu_inst_pe_1_6_0_U48 ( .A1(npu_inst_int_data_res_7__0__1_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N74), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N66), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n83) );
  INV_X1 npu_inst_pe_1_6_0_U47 ( .A(npu_inst_pe_1_6_0_n83), .ZN(
        npu_inst_pe_1_6_0_n99) );
  AOI222_X1 npu_inst_pe_1_6_0_U46 ( .A1(npu_inst_int_data_res_7__0__3_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N76), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N68), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n81) );
  INV_X1 npu_inst_pe_1_6_0_U45 ( .A(npu_inst_pe_1_6_0_n81), .ZN(
        npu_inst_pe_1_6_0_n36) );
  AOI222_X1 npu_inst_pe_1_6_0_U44 ( .A1(npu_inst_int_data_res_7__0__4_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N77), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N69), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n80) );
  INV_X1 npu_inst_pe_1_6_0_U43 ( .A(npu_inst_pe_1_6_0_n80), .ZN(
        npu_inst_pe_1_6_0_n35) );
  AOI222_X1 npu_inst_pe_1_6_0_U42 ( .A1(npu_inst_int_data_res_7__0__5_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N78), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N70), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n79) );
  INV_X1 npu_inst_pe_1_6_0_U41 ( .A(npu_inst_pe_1_6_0_n79), .ZN(
        npu_inst_pe_1_6_0_n34) );
  AOI222_X1 npu_inst_pe_1_6_0_U40 ( .A1(npu_inst_int_data_res_7__0__6_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N79), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N71), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n78) );
  INV_X1 npu_inst_pe_1_6_0_U39 ( .A(npu_inst_pe_1_6_0_n78), .ZN(
        npu_inst_pe_1_6_0_n33) );
  AND2_X1 npu_inst_pe_1_6_0_U38 ( .A1(npu_inst_pe_1_6_0_o_data_h_1_), .A2(
        npu_inst_pe_1_6_0_int_q_weight_1_), .ZN(npu_inst_pe_1_6_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_0_U37 ( .A1(npu_inst_pe_1_6_0_o_data_h_0_), .A2(
        npu_inst_pe_1_6_0_int_q_weight_1_), .ZN(npu_inst_pe_1_6_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_6_0_U36 ( .A(npu_inst_pe_1_6_0_int_data_1_), .ZN(
        npu_inst_pe_1_6_0_n13) );
  NOR3_X1 npu_inst_pe_1_6_0_U35 ( .A1(npu_inst_pe_1_6_0_n26), .A2(npu_inst_n36), .A3(npu_inst_int_ckg[15]), .ZN(npu_inst_pe_1_6_0_n85) );
  OR2_X1 npu_inst_pe_1_6_0_U34 ( .A1(npu_inst_pe_1_6_0_n85), .A2(
        npu_inst_pe_1_6_0_n1), .ZN(npu_inst_pe_1_6_0_N84) );
  AOI222_X1 npu_inst_pe_1_6_0_U33 ( .A1(npu_inst_int_data_res_7__0__2_), .A2(
        npu_inst_pe_1_6_0_n1), .B1(npu_inst_pe_1_6_0_N75), .B2(
        npu_inst_pe_1_6_0_n76), .C1(npu_inst_pe_1_6_0_N67), .C2(
        npu_inst_pe_1_6_0_n77), .ZN(npu_inst_pe_1_6_0_n82) );
  INV_X1 npu_inst_pe_1_6_0_U32 ( .A(npu_inst_pe_1_6_0_n82), .ZN(
        npu_inst_pe_1_6_0_n98) );
  AOI22_X1 npu_inst_pe_1_6_0_U31 ( .A1(npu_inst_n36), .A2(
        npu_inst_int_data_y_7__0__1_), .B1(npu_inst_pe_1_6_0_n2), .B2(
        npu_inst_int_data_x_6__1__1_), .ZN(npu_inst_pe_1_6_0_n63) );
  AOI22_X1 npu_inst_pe_1_6_0_U30 ( .A1(npu_inst_n36), .A2(
        npu_inst_int_data_y_7__0__0_), .B1(npu_inst_pe_1_6_0_n2), .B2(
        npu_inst_int_data_x_6__1__0_), .ZN(npu_inst_pe_1_6_0_n61) );
  INV_X1 npu_inst_pe_1_6_0_U29 ( .A(npu_inst_pe_1_6_0_int_data_0_), .ZN(
        npu_inst_pe_1_6_0_n12) );
  INV_X1 npu_inst_pe_1_6_0_U28 ( .A(npu_inst_n50), .ZN(npu_inst_pe_1_6_0_n4)
         );
  OR3_X1 npu_inst_pe_1_6_0_U27 ( .A1(npu_inst_pe_1_6_0_n5), .A2(
        npu_inst_pe_1_6_0_n7), .A3(npu_inst_pe_1_6_0_n4), .ZN(
        npu_inst_pe_1_6_0_n56) );
  OR3_X1 npu_inst_pe_1_6_0_U26 ( .A1(npu_inst_pe_1_6_0_n4), .A2(
        npu_inst_pe_1_6_0_n7), .A3(npu_inst_pe_1_6_0_n6), .ZN(
        npu_inst_pe_1_6_0_n48) );
  INV_X1 npu_inst_pe_1_6_0_U25 ( .A(npu_inst_pe_1_6_0_n4), .ZN(
        npu_inst_pe_1_6_0_n3) );
  OR3_X1 npu_inst_pe_1_6_0_U24 ( .A1(npu_inst_pe_1_6_0_n3), .A2(
        npu_inst_pe_1_6_0_n7), .A3(npu_inst_pe_1_6_0_n6), .ZN(
        npu_inst_pe_1_6_0_n52) );
  OR3_X1 npu_inst_pe_1_6_0_U23 ( .A1(npu_inst_pe_1_6_0_n5), .A2(
        npu_inst_pe_1_6_0_n7), .A3(npu_inst_pe_1_6_0_n3), .ZN(
        npu_inst_pe_1_6_0_n60) );
  BUF_X1 npu_inst_pe_1_6_0_U22 ( .A(npu_inst_n16), .Z(npu_inst_pe_1_6_0_n1) );
  NOR2_X1 npu_inst_pe_1_6_0_U21 ( .A1(npu_inst_pe_1_6_0_n60), .A2(
        npu_inst_pe_1_6_0_n2), .ZN(npu_inst_pe_1_6_0_n58) );
  NOR2_X1 npu_inst_pe_1_6_0_U20 ( .A1(npu_inst_pe_1_6_0_n56), .A2(
        npu_inst_pe_1_6_0_n2), .ZN(npu_inst_pe_1_6_0_n54) );
  NOR2_X1 npu_inst_pe_1_6_0_U19 ( .A1(npu_inst_pe_1_6_0_n52), .A2(
        npu_inst_pe_1_6_0_n2), .ZN(npu_inst_pe_1_6_0_n50) );
  NOR2_X1 npu_inst_pe_1_6_0_U18 ( .A1(npu_inst_pe_1_6_0_n48), .A2(
        npu_inst_pe_1_6_0_n2), .ZN(npu_inst_pe_1_6_0_n46) );
  NOR2_X1 npu_inst_pe_1_6_0_U17 ( .A1(npu_inst_pe_1_6_0_n40), .A2(
        npu_inst_pe_1_6_0_n2), .ZN(npu_inst_pe_1_6_0_n38) );
  NOR2_X1 npu_inst_pe_1_6_0_U16 ( .A1(npu_inst_pe_1_6_0_n44), .A2(
        npu_inst_pe_1_6_0_n2), .ZN(npu_inst_pe_1_6_0_n42) );
  BUF_X1 npu_inst_pe_1_6_0_U15 ( .A(npu_inst_n77), .Z(npu_inst_pe_1_6_0_n7) );
  INV_X1 npu_inst_pe_1_6_0_U14 ( .A(npu_inst_n105), .ZN(npu_inst_pe_1_6_0_n11)
         );
  INV_X1 npu_inst_pe_1_6_0_U13 ( .A(npu_inst_pe_1_6_0_n38), .ZN(
        npu_inst_pe_1_6_0_n113) );
  INV_X1 npu_inst_pe_1_6_0_U12 ( .A(npu_inst_pe_1_6_0_n58), .ZN(
        npu_inst_pe_1_6_0_n118) );
  INV_X1 npu_inst_pe_1_6_0_U11 ( .A(npu_inst_pe_1_6_0_n54), .ZN(
        npu_inst_pe_1_6_0_n117) );
  INV_X1 npu_inst_pe_1_6_0_U10 ( .A(npu_inst_pe_1_6_0_n50), .ZN(
        npu_inst_pe_1_6_0_n116) );
  INV_X1 npu_inst_pe_1_6_0_U9 ( .A(npu_inst_pe_1_6_0_n46), .ZN(
        npu_inst_pe_1_6_0_n115) );
  INV_X1 npu_inst_pe_1_6_0_U8 ( .A(npu_inst_pe_1_6_0_n42), .ZN(
        npu_inst_pe_1_6_0_n114) );
  BUF_X1 npu_inst_pe_1_6_0_U7 ( .A(npu_inst_pe_1_6_0_n11), .Z(
        npu_inst_pe_1_6_0_n10) );
  BUF_X1 npu_inst_pe_1_6_0_U6 ( .A(npu_inst_pe_1_6_0_n11), .Z(
        npu_inst_pe_1_6_0_n9) );
  BUF_X1 npu_inst_pe_1_6_0_U5 ( .A(npu_inst_pe_1_6_0_n11), .Z(
        npu_inst_pe_1_6_0_n8) );
  NOR2_X1 npu_inst_pe_1_6_0_U4 ( .A1(npu_inst_pe_1_6_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_0_n1), .ZN(npu_inst_pe_1_6_0_n76) );
  NOR2_X1 npu_inst_pe_1_6_0_U3 ( .A1(npu_inst_pe_1_6_0_n27), .A2(
        npu_inst_pe_1_6_0_n1), .ZN(npu_inst_pe_1_6_0_n77) );
  FA_X1 npu_inst_pe_1_6_0_sub_77_U2_1 ( .A(npu_inst_int_data_res_6__0__1_), 
        .B(npu_inst_pe_1_6_0_n13), .CI(npu_inst_pe_1_6_0_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_6_0_sub_77_carry_2_), .S(npu_inst_pe_1_6_0_N66) );
  FA_X1 npu_inst_pe_1_6_0_add_79_U1_1 ( .A(npu_inst_int_data_res_6__0__1_), 
        .B(npu_inst_pe_1_6_0_int_data_1_), .CI(
        npu_inst_pe_1_6_0_add_79_carry_1_), .CO(
        npu_inst_pe_1_6_0_add_79_carry_2_), .S(npu_inst_pe_1_6_0_N74) );
  NAND3_X1 npu_inst_pe_1_6_0_U101 ( .A1(npu_inst_pe_1_6_0_n4), .A2(
        npu_inst_pe_1_6_0_n6), .A3(npu_inst_pe_1_6_0_n7), .ZN(
        npu_inst_pe_1_6_0_n44) );
  NAND3_X1 npu_inst_pe_1_6_0_U100 ( .A1(npu_inst_pe_1_6_0_n3), .A2(
        npu_inst_pe_1_6_0_n6), .A3(npu_inst_pe_1_6_0_n7), .ZN(
        npu_inst_pe_1_6_0_n40) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_0_n33), .CK(
        npu_inst_pe_1_6_0_net3374), .RN(npu_inst_pe_1_6_0_n8), .Q(
        npu_inst_int_data_res_6__0__6_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_0_n34), .CK(
        npu_inst_pe_1_6_0_net3374), .RN(npu_inst_pe_1_6_0_n8), .Q(
        npu_inst_int_data_res_6__0__5_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_0_n35), .CK(
        npu_inst_pe_1_6_0_net3374), .RN(npu_inst_pe_1_6_0_n8), .Q(
        npu_inst_int_data_res_6__0__4_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_0_n36), .CK(
        npu_inst_pe_1_6_0_net3374), .RN(npu_inst_pe_1_6_0_n8), .Q(
        npu_inst_int_data_res_6__0__3_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_0_n98), .CK(
        npu_inst_pe_1_6_0_net3374), .RN(npu_inst_pe_1_6_0_n8), .Q(
        npu_inst_int_data_res_6__0__2_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_0_n99), .CK(
        npu_inst_pe_1_6_0_net3374), .RN(npu_inst_pe_1_6_0_n8), .Q(
        npu_inst_int_data_res_6__0__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_0_n32), .CK(
        npu_inst_pe_1_6_0_net3374), .RN(npu_inst_pe_1_6_0_n8), .Q(
        npu_inst_int_data_res_6__0__7_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_0_n100), 
        .CK(npu_inst_pe_1_6_0_net3374), .RN(npu_inst_pe_1_6_0_n8), .Q(
        npu_inst_int_data_res_6__0__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_weight_reg_0_ ( .D(npu_inst_n91), .CK(
        npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n8), .Q(
        npu_inst_pe_1_6_0_int_q_weight_0_), .QN(npu_inst_pe_1_6_0_n27) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_weight_reg_1_ ( .D(npu_inst_n97), .CK(
        npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n8), .Q(
        npu_inst_pe_1_6_0_int_q_weight_1_), .QN(npu_inst_pe_1_6_0_n26) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_0_n112), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n8), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_0_n106), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n8), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_0_n111), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_0_n105), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_0_n110), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_0_n104), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_0_n109), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_0_n103), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_0_n108), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_0_n102), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_0_n107), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_0_n101), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_0_n86), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_0_n87), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n9), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_0_n88), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_0_n89), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_0_n90), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_0_n91), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_0_n92), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_0_n93), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_0_n94), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_0_n95), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_0_n96), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_0_n97), 
        .CK(npu_inst_pe_1_6_0_net3380), .RN(npu_inst_pe_1_6_0_n10), .Q(
        npu_inst_pe_1_6_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_0_net3374) );
  CLKGATETST_X1 npu_inst_pe_1_6_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n44), .SE(1'b0), .GCK(npu_inst_pe_1_6_0_net3380) );
  MUX2_X1 npu_inst_pe_1_6_1_U153 ( .A(npu_inst_pe_1_6_1_n31), .B(
        npu_inst_pe_1_6_1_n28), .S(npu_inst_pe_1_6_1_n7), .Z(
        npu_inst_pe_1_6_1_N93) );
  MUX2_X1 npu_inst_pe_1_6_1_U152 ( .A(npu_inst_pe_1_6_1_n30), .B(
        npu_inst_pe_1_6_1_n29), .S(npu_inst_pe_1_6_1_n5), .Z(
        npu_inst_pe_1_6_1_n31) );
  MUX2_X1 npu_inst_pe_1_6_1_U151 ( .A(npu_inst_pe_1_6_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_1_n3), .Z(
        npu_inst_pe_1_6_1_n30) );
  MUX2_X1 npu_inst_pe_1_6_1_U150 ( .A(npu_inst_pe_1_6_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_1_n3), .Z(
        npu_inst_pe_1_6_1_n29) );
  MUX2_X1 npu_inst_pe_1_6_1_U149 ( .A(npu_inst_pe_1_6_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_1_n3), .Z(
        npu_inst_pe_1_6_1_n28) );
  MUX2_X1 npu_inst_pe_1_6_1_U148 ( .A(npu_inst_pe_1_6_1_n25), .B(
        npu_inst_pe_1_6_1_n22), .S(npu_inst_pe_1_6_1_n7), .Z(
        npu_inst_pe_1_6_1_N94) );
  MUX2_X1 npu_inst_pe_1_6_1_U147 ( .A(npu_inst_pe_1_6_1_n24), .B(
        npu_inst_pe_1_6_1_n23), .S(npu_inst_pe_1_6_1_n5), .Z(
        npu_inst_pe_1_6_1_n25) );
  MUX2_X1 npu_inst_pe_1_6_1_U146 ( .A(npu_inst_pe_1_6_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_1_n3), .Z(
        npu_inst_pe_1_6_1_n24) );
  MUX2_X1 npu_inst_pe_1_6_1_U145 ( .A(npu_inst_pe_1_6_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_1_n3), .Z(
        npu_inst_pe_1_6_1_n23) );
  MUX2_X1 npu_inst_pe_1_6_1_U144 ( .A(npu_inst_pe_1_6_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_1_n3), .Z(
        npu_inst_pe_1_6_1_n22) );
  MUX2_X1 npu_inst_pe_1_6_1_U143 ( .A(npu_inst_pe_1_6_1_n21), .B(
        npu_inst_pe_1_6_1_n18), .S(npu_inst_pe_1_6_1_n7), .Z(
        npu_inst_int_data_x_6__1__1_) );
  MUX2_X1 npu_inst_pe_1_6_1_U142 ( .A(npu_inst_pe_1_6_1_n20), .B(
        npu_inst_pe_1_6_1_n19), .S(npu_inst_pe_1_6_1_n5), .Z(
        npu_inst_pe_1_6_1_n21) );
  MUX2_X1 npu_inst_pe_1_6_1_U141 ( .A(npu_inst_pe_1_6_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_1_n3), .Z(
        npu_inst_pe_1_6_1_n20) );
  MUX2_X1 npu_inst_pe_1_6_1_U140 ( .A(npu_inst_pe_1_6_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_1_n3), .Z(
        npu_inst_pe_1_6_1_n19) );
  MUX2_X1 npu_inst_pe_1_6_1_U139 ( .A(npu_inst_pe_1_6_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_1_n3), .Z(
        npu_inst_pe_1_6_1_n18) );
  MUX2_X1 npu_inst_pe_1_6_1_U138 ( .A(npu_inst_pe_1_6_1_n17), .B(
        npu_inst_pe_1_6_1_n14), .S(npu_inst_pe_1_6_1_n7), .Z(
        npu_inst_int_data_x_6__1__0_) );
  MUX2_X1 npu_inst_pe_1_6_1_U137 ( .A(npu_inst_pe_1_6_1_n16), .B(
        npu_inst_pe_1_6_1_n15), .S(npu_inst_pe_1_6_1_n5), .Z(
        npu_inst_pe_1_6_1_n17) );
  MUX2_X1 npu_inst_pe_1_6_1_U136 ( .A(npu_inst_pe_1_6_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_1_n3), .Z(
        npu_inst_pe_1_6_1_n16) );
  MUX2_X1 npu_inst_pe_1_6_1_U135 ( .A(npu_inst_pe_1_6_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_1_n3), .Z(
        npu_inst_pe_1_6_1_n15) );
  MUX2_X1 npu_inst_pe_1_6_1_U134 ( .A(npu_inst_pe_1_6_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_1_n3), .Z(
        npu_inst_pe_1_6_1_n14) );
  XOR2_X1 npu_inst_pe_1_6_1_U133 ( .A(npu_inst_pe_1_6_1_int_data_0_), .B(
        npu_inst_int_data_res_6__1__0_), .Z(npu_inst_pe_1_6_1_N73) );
  AND2_X1 npu_inst_pe_1_6_1_U132 ( .A1(npu_inst_int_data_res_6__1__0_), .A2(
        npu_inst_pe_1_6_1_int_data_0_), .ZN(npu_inst_pe_1_6_1_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_1_U131 ( .A(npu_inst_int_data_res_6__1__0_), .B(
        npu_inst_pe_1_6_1_n12), .ZN(npu_inst_pe_1_6_1_N65) );
  OR2_X1 npu_inst_pe_1_6_1_U130 ( .A1(npu_inst_pe_1_6_1_n12), .A2(
        npu_inst_int_data_res_6__1__0_), .ZN(npu_inst_pe_1_6_1_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_1_U129 ( .A(npu_inst_int_data_res_6__1__2_), .B(
        npu_inst_pe_1_6_1_add_79_carry_2_), .Z(npu_inst_pe_1_6_1_N75) );
  AND2_X1 npu_inst_pe_1_6_1_U128 ( .A1(npu_inst_pe_1_6_1_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_6__1__2_), .ZN(
        npu_inst_pe_1_6_1_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_1_U127 ( .A(npu_inst_int_data_res_6__1__3_), .B(
        npu_inst_pe_1_6_1_add_79_carry_3_), .Z(npu_inst_pe_1_6_1_N76) );
  AND2_X1 npu_inst_pe_1_6_1_U126 ( .A1(npu_inst_pe_1_6_1_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_6__1__3_), .ZN(
        npu_inst_pe_1_6_1_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_1_U125 ( .A(npu_inst_int_data_res_6__1__4_), .B(
        npu_inst_pe_1_6_1_add_79_carry_4_), .Z(npu_inst_pe_1_6_1_N77) );
  AND2_X1 npu_inst_pe_1_6_1_U124 ( .A1(npu_inst_pe_1_6_1_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_6__1__4_), .ZN(
        npu_inst_pe_1_6_1_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_1_U123 ( .A(npu_inst_int_data_res_6__1__5_), .B(
        npu_inst_pe_1_6_1_add_79_carry_5_), .Z(npu_inst_pe_1_6_1_N78) );
  AND2_X1 npu_inst_pe_1_6_1_U122 ( .A1(npu_inst_pe_1_6_1_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_6__1__5_), .ZN(
        npu_inst_pe_1_6_1_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_1_U121 ( .A(npu_inst_int_data_res_6__1__6_), .B(
        npu_inst_pe_1_6_1_add_79_carry_6_), .Z(npu_inst_pe_1_6_1_N79) );
  AND2_X1 npu_inst_pe_1_6_1_U120 ( .A1(npu_inst_pe_1_6_1_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_6__1__6_), .ZN(
        npu_inst_pe_1_6_1_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_1_U119 ( .A(npu_inst_int_data_res_6__1__7_), .B(
        npu_inst_pe_1_6_1_add_79_carry_7_), .Z(npu_inst_pe_1_6_1_N80) );
  XNOR2_X1 npu_inst_pe_1_6_1_U118 ( .A(npu_inst_pe_1_6_1_sub_77_carry_2_), .B(
        npu_inst_int_data_res_6__1__2_), .ZN(npu_inst_pe_1_6_1_N67) );
  OR2_X1 npu_inst_pe_1_6_1_U117 ( .A1(npu_inst_int_data_res_6__1__2_), .A2(
        npu_inst_pe_1_6_1_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_6_1_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_1_U116 ( .A(npu_inst_pe_1_6_1_sub_77_carry_3_), .B(
        npu_inst_int_data_res_6__1__3_), .ZN(npu_inst_pe_1_6_1_N68) );
  OR2_X1 npu_inst_pe_1_6_1_U115 ( .A1(npu_inst_int_data_res_6__1__3_), .A2(
        npu_inst_pe_1_6_1_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_6_1_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_1_U114 ( .A(npu_inst_pe_1_6_1_sub_77_carry_4_), .B(
        npu_inst_int_data_res_6__1__4_), .ZN(npu_inst_pe_1_6_1_N69) );
  OR2_X1 npu_inst_pe_1_6_1_U113 ( .A1(npu_inst_int_data_res_6__1__4_), .A2(
        npu_inst_pe_1_6_1_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_6_1_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_1_U112 ( .A(npu_inst_pe_1_6_1_sub_77_carry_5_), .B(
        npu_inst_int_data_res_6__1__5_), .ZN(npu_inst_pe_1_6_1_N70) );
  OR2_X1 npu_inst_pe_1_6_1_U111 ( .A1(npu_inst_int_data_res_6__1__5_), .A2(
        npu_inst_pe_1_6_1_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_6_1_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_1_U110 ( .A(npu_inst_pe_1_6_1_sub_77_carry_6_), .B(
        npu_inst_int_data_res_6__1__6_), .ZN(npu_inst_pe_1_6_1_N71) );
  OR2_X1 npu_inst_pe_1_6_1_U109 ( .A1(npu_inst_int_data_res_6__1__6_), .A2(
        npu_inst_pe_1_6_1_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_6_1_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_1_U108 ( .A(npu_inst_int_data_res_6__1__7_), .B(
        npu_inst_pe_1_6_1_sub_77_carry_7_), .ZN(npu_inst_pe_1_6_1_N72) );
  INV_X1 npu_inst_pe_1_6_1_U107 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_6_1_n6)
         );
  INV_X1 npu_inst_pe_1_6_1_U106 ( .A(npu_inst_pe_1_6_1_n6), .ZN(
        npu_inst_pe_1_6_1_n5) );
  INV_X1 npu_inst_pe_1_6_1_U105 ( .A(npu_inst_n36), .ZN(npu_inst_pe_1_6_1_n2)
         );
  AOI22_X1 npu_inst_pe_1_6_1_U104 ( .A1(npu_inst_int_data_y_7__1__0_), .A2(
        npu_inst_pe_1_6_1_n58), .B1(npu_inst_pe_1_6_1_n118), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_1_n57) );
  INV_X1 npu_inst_pe_1_6_1_U103 ( .A(npu_inst_pe_1_6_1_n57), .ZN(
        npu_inst_pe_1_6_1_n107) );
  AOI22_X1 npu_inst_pe_1_6_1_U102 ( .A1(npu_inst_int_data_y_7__1__0_), .A2(
        npu_inst_pe_1_6_1_n54), .B1(npu_inst_pe_1_6_1_n117), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_1_n53) );
  INV_X1 npu_inst_pe_1_6_1_U99 ( .A(npu_inst_pe_1_6_1_n53), .ZN(
        npu_inst_pe_1_6_1_n108) );
  AOI22_X1 npu_inst_pe_1_6_1_U98 ( .A1(npu_inst_int_data_y_7__1__0_), .A2(
        npu_inst_pe_1_6_1_n50), .B1(npu_inst_pe_1_6_1_n116), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_1_n49) );
  INV_X1 npu_inst_pe_1_6_1_U97 ( .A(npu_inst_pe_1_6_1_n49), .ZN(
        npu_inst_pe_1_6_1_n109) );
  AOI22_X1 npu_inst_pe_1_6_1_U96 ( .A1(npu_inst_int_data_y_7__1__0_), .A2(
        npu_inst_pe_1_6_1_n46), .B1(npu_inst_pe_1_6_1_n115), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_1_n45) );
  INV_X1 npu_inst_pe_1_6_1_U95 ( .A(npu_inst_pe_1_6_1_n45), .ZN(
        npu_inst_pe_1_6_1_n110) );
  AOI22_X1 npu_inst_pe_1_6_1_U94 ( .A1(npu_inst_int_data_y_7__1__0_), .A2(
        npu_inst_pe_1_6_1_n42), .B1(npu_inst_pe_1_6_1_n114), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_1_n41) );
  INV_X1 npu_inst_pe_1_6_1_U93 ( .A(npu_inst_pe_1_6_1_n41), .ZN(
        npu_inst_pe_1_6_1_n111) );
  AOI22_X1 npu_inst_pe_1_6_1_U92 ( .A1(npu_inst_int_data_y_7__1__1_), .A2(
        npu_inst_pe_1_6_1_n58), .B1(npu_inst_pe_1_6_1_n118), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_1_n59) );
  INV_X1 npu_inst_pe_1_6_1_U91 ( .A(npu_inst_pe_1_6_1_n59), .ZN(
        npu_inst_pe_1_6_1_n101) );
  AOI22_X1 npu_inst_pe_1_6_1_U90 ( .A1(npu_inst_int_data_y_7__1__1_), .A2(
        npu_inst_pe_1_6_1_n54), .B1(npu_inst_pe_1_6_1_n117), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_1_n55) );
  INV_X1 npu_inst_pe_1_6_1_U89 ( .A(npu_inst_pe_1_6_1_n55), .ZN(
        npu_inst_pe_1_6_1_n102) );
  AOI22_X1 npu_inst_pe_1_6_1_U88 ( .A1(npu_inst_int_data_y_7__1__1_), .A2(
        npu_inst_pe_1_6_1_n50), .B1(npu_inst_pe_1_6_1_n116), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_1_n51) );
  INV_X1 npu_inst_pe_1_6_1_U87 ( .A(npu_inst_pe_1_6_1_n51), .ZN(
        npu_inst_pe_1_6_1_n103) );
  AOI22_X1 npu_inst_pe_1_6_1_U86 ( .A1(npu_inst_int_data_y_7__1__1_), .A2(
        npu_inst_pe_1_6_1_n46), .B1(npu_inst_pe_1_6_1_n115), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_1_n47) );
  INV_X1 npu_inst_pe_1_6_1_U85 ( .A(npu_inst_pe_1_6_1_n47), .ZN(
        npu_inst_pe_1_6_1_n104) );
  AOI22_X1 npu_inst_pe_1_6_1_U84 ( .A1(npu_inst_int_data_y_7__1__1_), .A2(
        npu_inst_pe_1_6_1_n42), .B1(npu_inst_pe_1_6_1_n114), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_1_n43) );
  INV_X1 npu_inst_pe_1_6_1_U83 ( .A(npu_inst_pe_1_6_1_n43), .ZN(
        npu_inst_pe_1_6_1_n105) );
  AOI22_X1 npu_inst_pe_1_6_1_U82 ( .A1(npu_inst_pe_1_6_1_n38), .A2(
        npu_inst_int_data_y_7__1__1_), .B1(npu_inst_pe_1_6_1_n113), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_1_n39) );
  INV_X1 npu_inst_pe_1_6_1_U81 ( .A(npu_inst_pe_1_6_1_n39), .ZN(
        npu_inst_pe_1_6_1_n106) );
  AND2_X1 npu_inst_pe_1_6_1_U80 ( .A1(npu_inst_pe_1_6_1_N93), .A2(npu_inst_n36), .ZN(npu_inst_int_data_y_6__1__0_) );
  NAND2_X1 npu_inst_pe_1_6_1_U79 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_1_n60), .ZN(npu_inst_pe_1_6_1_n74) );
  OAI21_X1 npu_inst_pe_1_6_1_U78 ( .B1(npu_inst_pe_1_6_1_n63), .B2(
        npu_inst_pe_1_6_1_n60), .A(npu_inst_pe_1_6_1_n74), .ZN(
        npu_inst_pe_1_6_1_n97) );
  NAND2_X1 npu_inst_pe_1_6_1_U77 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_1_n60), .ZN(npu_inst_pe_1_6_1_n73) );
  OAI21_X1 npu_inst_pe_1_6_1_U76 ( .B1(npu_inst_pe_1_6_1_n61), .B2(
        npu_inst_pe_1_6_1_n60), .A(npu_inst_pe_1_6_1_n73), .ZN(
        npu_inst_pe_1_6_1_n96) );
  NAND2_X1 npu_inst_pe_1_6_1_U75 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_1_n56), .ZN(npu_inst_pe_1_6_1_n72) );
  OAI21_X1 npu_inst_pe_1_6_1_U74 ( .B1(npu_inst_pe_1_6_1_n63), .B2(
        npu_inst_pe_1_6_1_n56), .A(npu_inst_pe_1_6_1_n72), .ZN(
        npu_inst_pe_1_6_1_n95) );
  NAND2_X1 npu_inst_pe_1_6_1_U73 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_1_n56), .ZN(npu_inst_pe_1_6_1_n71) );
  OAI21_X1 npu_inst_pe_1_6_1_U72 ( .B1(npu_inst_pe_1_6_1_n61), .B2(
        npu_inst_pe_1_6_1_n56), .A(npu_inst_pe_1_6_1_n71), .ZN(
        npu_inst_pe_1_6_1_n94) );
  NAND2_X1 npu_inst_pe_1_6_1_U71 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_1_n52), .ZN(npu_inst_pe_1_6_1_n70) );
  OAI21_X1 npu_inst_pe_1_6_1_U70 ( .B1(npu_inst_pe_1_6_1_n63), .B2(
        npu_inst_pe_1_6_1_n52), .A(npu_inst_pe_1_6_1_n70), .ZN(
        npu_inst_pe_1_6_1_n93) );
  NAND2_X1 npu_inst_pe_1_6_1_U69 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_1_n52), .ZN(npu_inst_pe_1_6_1_n69) );
  OAI21_X1 npu_inst_pe_1_6_1_U68 ( .B1(npu_inst_pe_1_6_1_n61), .B2(
        npu_inst_pe_1_6_1_n52), .A(npu_inst_pe_1_6_1_n69), .ZN(
        npu_inst_pe_1_6_1_n92) );
  NAND2_X1 npu_inst_pe_1_6_1_U67 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_1_n48), .ZN(npu_inst_pe_1_6_1_n68) );
  OAI21_X1 npu_inst_pe_1_6_1_U66 ( .B1(npu_inst_pe_1_6_1_n63), .B2(
        npu_inst_pe_1_6_1_n48), .A(npu_inst_pe_1_6_1_n68), .ZN(
        npu_inst_pe_1_6_1_n91) );
  NAND2_X1 npu_inst_pe_1_6_1_U65 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_1_n48), .ZN(npu_inst_pe_1_6_1_n67) );
  OAI21_X1 npu_inst_pe_1_6_1_U64 ( .B1(npu_inst_pe_1_6_1_n61), .B2(
        npu_inst_pe_1_6_1_n48), .A(npu_inst_pe_1_6_1_n67), .ZN(
        npu_inst_pe_1_6_1_n90) );
  NAND2_X1 npu_inst_pe_1_6_1_U63 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_1_n44), .ZN(npu_inst_pe_1_6_1_n66) );
  OAI21_X1 npu_inst_pe_1_6_1_U62 ( .B1(npu_inst_pe_1_6_1_n63), .B2(
        npu_inst_pe_1_6_1_n44), .A(npu_inst_pe_1_6_1_n66), .ZN(
        npu_inst_pe_1_6_1_n89) );
  NAND2_X1 npu_inst_pe_1_6_1_U61 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_1_n44), .ZN(npu_inst_pe_1_6_1_n65) );
  OAI21_X1 npu_inst_pe_1_6_1_U60 ( .B1(npu_inst_pe_1_6_1_n61), .B2(
        npu_inst_pe_1_6_1_n44), .A(npu_inst_pe_1_6_1_n65), .ZN(
        npu_inst_pe_1_6_1_n88) );
  NAND2_X1 npu_inst_pe_1_6_1_U59 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_1_n40), .ZN(npu_inst_pe_1_6_1_n64) );
  OAI21_X1 npu_inst_pe_1_6_1_U58 ( .B1(npu_inst_pe_1_6_1_n63), .B2(
        npu_inst_pe_1_6_1_n40), .A(npu_inst_pe_1_6_1_n64), .ZN(
        npu_inst_pe_1_6_1_n87) );
  NAND2_X1 npu_inst_pe_1_6_1_U57 ( .A1(npu_inst_pe_1_6_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_1_n40), .ZN(npu_inst_pe_1_6_1_n62) );
  OAI21_X1 npu_inst_pe_1_6_1_U56 ( .B1(npu_inst_pe_1_6_1_n61), .B2(
        npu_inst_pe_1_6_1_n40), .A(npu_inst_pe_1_6_1_n62), .ZN(
        npu_inst_pe_1_6_1_n86) );
  AOI22_X1 npu_inst_pe_1_6_1_U55 ( .A1(npu_inst_pe_1_6_1_n38), .A2(
        npu_inst_int_data_y_7__1__0_), .B1(npu_inst_pe_1_6_1_n113), .B2(
        npu_inst_pe_1_6_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_1_n37) );
  INV_X1 npu_inst_pe_1_6_1_U54 ( .A(npu_inst_pe_1_6_1_n37), .ZN(
        npu_inst_pe_1_6_1_n112) );
  AND2_X1 npu_inst_pe_1_6_1_U53 ( .A1(npu_inst_n36), .A2(npu_inst_pe_1_6_1_N94), .ZN(npu_inst_int_data_y_6__1__1_) );
  AOI222_X1 npu_inst_pe_1_6_1_U52 ( .A1(npu_inst_int_data_res_7__1__0_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N73), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N65), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n84) );
  INV_X1 npu_inst_pe_1_6_1_U51 ( .A(npu_inst_pe_1_6_1_n84), .ZN(
        npu_inst_pe_1_6_1_n100) );
  AOI222_X1 npu_inst_pe_1_6_1_U50 ( .A1(npu_inst_pe_1_6_1_n1), .A2(
        npu_inst_int_data_res_7__1__7_), .B1(npu_inst_pe_1_6_1_N80), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N72), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n75) );
  INV_X1 npu_inst_pe_1_6_1_U49 ( .A(npu_inst_pe_1_6_1_n75), .ZN(
        npu_inst_pe_1_6_1_n32) );
  AOI222_X1 npu_inst_pe_1_6_1_U48 ( .A1(npu_inst_int_data_res_7__1__1_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N74), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N66), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n83) );
  INV_X1 npu_inst_pe_1_6_1_U47 ( .A(npu_inst_pe_1_6_1_n83), .ZN(
        npu_inst_pe_1_6_1_n99) );
  AOI222_X1 npu_inst_pe_1_6_1_U46 ( .A1(npu_inst_int_data_res_7__1__3_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N76), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N68), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n81) );
  INV_X1 npu_inst_pe_1_6_1_U45 ( .A(npu_inst_pe_1_6_1_n81), .ZN(
        npu_inst_pe_1_6_1_n36) );
  AOI222_X1 npu_inst_pe_1_6_1_U44 ( .A1(npu_inst_int_data_res_7__1__4_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N77), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N69), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n80) );
  INV_X1 npu_inst_pe_1_6_1_U43 ( .A(npu_inst_pe_1_6_1_n80), .ZN(
        npu_inst_pe_1_6_1_n35) );
  AOI222_X1 npu_inst_pe_1_6_1_U42 ( .A1(npu_inst_int_data_res_7__1__5_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N78), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N70), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n79) );
  INV_X1 npu_inst_pe_1_6_1_U41 ( .A(npu_inst_pe_1_6_1_n79), .ZN(
        npu_inst_pe_1_6_1_n34) );
  AOI222_X1 npu_inst_pe_1_6_1_U40 ( .A1(npu_inst_int_data_res_7__1__6_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N79), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N71), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n78) );
  INV_X1 npu_inst_pe_1_6_1_U39 ( .A(npu_inst_pe_1_6_1_n78), .ZN(
        npu_inst_pe_1_6_1_n33) );
  AND2_X1 npu_inst_pe_1_6_1_U38 ( .A1(npu_inst_int_data_x_6__1__1_), .A2(
        npu_inst_pe_1_6_1_int_q_weight_1_), .ZN(npu_inst_pe_1_6_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_1_U37 ( .A1(npu_inst_int_data_x_6__1__0_), .A2(
        npu_inst_pe_1_6_1_int_q_weight_1_), .ZN(npu_inst_pe_1_6_1_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_6_1_U36 ( .A(npu_inst_pe_1_6_1_int_data_1_), .ZN(
        npu_inst_pe_1_6_1_n13) );
  NOR3_X1 npu_inst_pe_1_6_1_U35 ( .A1(npu_inst_pe_1_6_1_n26), .A2(npu_inst_n36), .A3(npu_inst_int_ckg[14]), .ZN(npu_inst_pe_1_6_1_n85) );
  OR2_X1 npu_inst_pe_1_6_1_U34 ( .A1(npu_inst_pe_1_6_1_n85), .A2(
        npu_inst_pe_1_6_1_n1), .ZN(npu_inst_pe_1_6_1_N84) );
  AOI222_X1 npu_inst_pe_1_6_1_U33 ( .A1(npu_inst_int_data_res_7__1__2_), .A2(
        npu_inst_pe_1_6_1_n1), .B1(npu_inst_pe_1_6_1_N75), .B2(
        npu_inst_pe_1_6_1_n76), .C1(npu_inst_pe_1_6_1_N67), .C2(
        npu_inst_pe_1_6_1_n77), .ZN(npu_inst_pe_1_6_1_n82) );
  INV_X1 npu_inst_pe_1_6_1_U32 ( .A(npu_inst_pe_1_6_1_n82), .ZN(
        npu_inst_pe_1_6_1_n98) );
  AOI22_X1 npu_inst_pe_1_6_1_U31 ( .A1(npu_inst_n36), .A2(
        npu_inst_int_data_y_7__1__1_), .B1(npu_inst_pe_1_6_1_n2), .B2(
        npu_inst_int_data_x_6__2__1_), .ZN(npu_inst_pe_1_6_1_n63) );
  AOI22_X1 npu_inst_pe_1_6_1_U30 ( .A1(npu_inst_n36), .A2(
        npu_inst_int_data_y_7__1__0_), .B1(npu_inst_pe_1_6_1_n2), .B2(
        npu_inst_int_data_x_6__2__0_), .ZN(npu_inst_pe_1_6_1_n61) );
  INV_X1 npu_inst_pe_1_6_1_U29 ( .A(npu_inst_pe_1_6_1_int_data_0_), .ZN(
        npu_inst_pe_1_6_1_n12) );
  INV_X1 npu_inst_pe_1_6_1_U28 ( .A(npu_inst_n50), .ZN(npu_inst_pe_1_6_1_n4)
         );
  OR3_X1 npu_inst_pe_1_6_1_U27 ( .A1(npu_inst_pe_1_6_1_n5), .A2(
        npu_inst_pe_1_6_1_n7), .A3(npu_inst_pe_1_6_1_n4), .ZN(
        npu_inst_pe_1_6_1_n56) );
  OR3_X1 npu_inst_pe_1_6_1_U26 ( .A1(npu_inst_pe_1_6_1_n4), .A2(
        npu_inst_pe_1_6_1_n7), .A3(npu_inst_pe_1_6_1_n6), .ZN(
        npu_inst_pe_1_6_1_n48) );
  INV_X1 npu_inst_pe_1_6_1_U25 ( .A(npu_inst_pe_1_6_1_n4), .ZN(
        npu_inst_pe_1_6_1_n3) );
  OR3_X1 npu_inst_pe_1_6_1_U24 ( .A1(npu_inst_pe_1_6_1_n3), .A2(
        npu_inst_pe_1_6_1_n7), .A3(npu_inst_pe_1_6_1_n6), .ZN(
        npu_inst_pe_1_6_1_n52) );
  OR3_X1 npu_inst_pe_1_6_1_U23 ( .A1(npu_inst_pe_1_6_1_n5), .A2(
        npu_inst_pe_1_6_1_n7), .A3(npu_inst_pe_1_6_1_n3), .ZN(
        npu_inst_pe_1_6_1_n60) );
  BUF_X1 npu_inst_pe_1_6_1_U22 ( .A(npu_inst_n15), .Z(npu_inst_pe_1_6_1_n1) );
  NOR2_X1 npu_inst_pe_1_6_1_U21 ( .A1(npu_inst_pe_1_6_1_n60), .A2(
        npu_inst_pe_1_6_1_n2), .ZN(npu_inst_pe_1_6_1_n58) );
  NOR2_X1 npu_inst_pe_1_6_1_U20 ( .A1(npu_inst_pe_1_6_1_n56), .A2(
        npu_inst_pe_1_6_1_n2), .ZN(npu_inst_pe_1_6_1_n54) );
  NOR2_X1 npu_inst_pe_1_6_1_U19 ( .A1(npu_inst_pe_1_6_1_n52), .A2(
        npu_inst_pe_1_6_1_n2), .ZN(npu_inst_pe_1_6_1_n50) );
  NOR2_X1 npu_inst_pe_1_6_1_U18 ( .A1(npu_inst_pe_1_6_1_n48), .A2(
        npu_inst_pe_1_6_1_n2), .ZN(npu_inst_pe_1_6_1_n46) );
  NOR2_X1 npu_inst_pe_1_6_1_U17 ( .A1(npu_inst_pe_1_6_1_n40), .A2(
        npu_inst_pe_1_6_1_n2), .ZN(npu_inst_pe_1_6_1_n38) );
  NOR2_X1 npu_inst_pe_1_6_1_U16 ( .A1(npu_inst_pe_1_6_1_n44), .A2(
        npu_inst_pe_1_6_1_n2), .ZN(npu_inst_pe_1_6_1_n42) );
  BUF_X1 npu_inst_pe_1_6_1_U15 ( .A(npu_inst_n77), .Z(npu_inst_pe_1_6_1_n7) );
  INV_X1 npu_inst_pe_1_6_1_U14 ( .A(npu_inst_n105), .ZN(npu_inst_pe_1_6_1_n11)
         );
  INV_X1 npu_inst_pe_1_6_1_U13 ( .A(npu_inst_pe_1_6_1_n38), .ZN(
        npu_inst_pe_1_6_1_n113) );
  INV_X1 npu_inst_pe_1_6_1_U12 ( .A(npu_inst_pe_1_6_1_n58), .ZN(
        npu_inst_pe_1_6_1_n118) );
  INV_X1 npu_inst_pe_1_6_1_U11 ( .A(npu_inst_pe_1_6_1_n54), .ZN(
        npu_inst_pe_1_6_1_n117) );
  INV_X1 npu_inst_pe_1_6_1_U10 ( .A(npu_inst_pe_1_6_1_n50), .ZN(
        npu_inst_pe_1_6_1_n116) );
  INV_X1 npu_inst_pe_1_6_1_U9 ( .A(npu_inst_pe_1_6_1_n46), .ZN(
        npu_inst_pe_1_6_1_n115) );
  INV_X1 npu_inst_pe_1_6_1_U8 ( .A(npu_inst_pe_1_6_1_n42), .ZN(
        npu_inst_pe_1_6_1_n114) );
  BUF_X1 npu_inst_pe_1_6_1_U7 ( .A(npu_inst_pe_1_6_1_n11), .Z(
        npu_inst_pe_1_6_1_n10) );
  BUF_X1 npu_inst_pe_1_6_1_U6 ( .A(npu_inst_pe_1_6_1_n11), .Z(
        npu_inst_pe_1_6_1_n9) );
  BUF_X1 npu_inst_pe_1_6_1_U5 ( .A(npu_inst_pe_1_6_1_n11), .Z(
        npu_inst_pe_1_6_1_n8) );
  NOR2_X1 npu_inst_pe_1_6_1_U4 ( .A1(npu_inst_pe_1_6_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_1_n1), .ZN(npu_inst_pe_1_6_1_n76) );
  NOR2_X1 npu_inst_pe_1_6_1_U3 ( .A1(npu_inst_pe_1_6_1_n27), .A2(
        npu_inst_pe_1_6_1_n1), .ZN(npu_inst_pe_1_6_1_n77) );
  FA_X1 npu_inst_pe_1_6_1_sub_77_U2_1 ( .A(npu_inst_int_data_res_6__1__1_), 
        .B(npu_inst_pe_1_6_1_n13), .CI(npu_inst_pe_1_6_1_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_6_1_sub_77_carry_2_), .S(npu_inst_pe_1_6_1_N66) );
  FA_X1 npu_inst_pe_1_6_1_add_79_U1_1 ( .A(npu_inst_int_data_res_6__1__1_), 
        .B(npu_inst_pe_1_6_1_int_data_1_), .CI(
        npu_inst_pe_1_6_1_add_79_carry_1_), .CO(
        npu_inst_pe_1_6_1_add_79_carry_2_), .S(npu_inst_pe_1_6_1_N74) );
  NAND3_X1 npu_inst_pe_1_6_1_U101 ( .A1(npu_inst_pe_1_6_1_n4), .A2(
        npu_inst_pe_1_6_1_n6), .A3(npu_inst_pe_1_6_1_n7), .ZN(
        npu_inst_pe_1_6_1_n44) );
  NAND3_X1 npu_inst_pe_1_6_1_U100 ( .A1(npu_inst_pe_1_6_1_n3), .A2(
        npu_inst_pe_1_6_1_n6), .A3(npu_inst_pe_1_6_1_n7), .ZN(
        npu_inst_pe_1_6_1_n40) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_1_n33), .CK(
        npu_inst_pe_1_6_1_net3351), .RN(npu_inst_pe_1_6_1_n8), .Q(
        npu_inst_int_data_res_6__1__6_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_1_n34), .CK(
        npu_inst_pe_1_6_1_net3351), .RN(npu_inst_pe_1_6_1_n8), .Q(
        npu_inst_int_data_res_6__1__5_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_1_n35), .CK(
        npu_inst_pe_1_6_1_net3351), .RN(npu_inst_pe_1_6_1_n8), .Q(
        npu_inst_int_data_res_6__1__4_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_1_n36), .CK(
        npu_inst_pe_1_6_1_net3351), .RN(npu_inst_pe_1_6_1_n8), .Q(
        npu_inst_int_data_res_6__1__3_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_1_n98), .CK(
        npu_inst_pe_1_6_1_net3351), .RN(npu_inst_pe_1_6_1_n8), .Q(
        npu_inst_int_data_res_6__1__2_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_1_n99), .CK(
        npu_inst_pe_1_6_1_net3351), .RN(npu_inst_pe_1_6_1_n8), .Q(
        npu_inst_int_data_res_6__1__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_1_n32), .CK(
        npu_inst_pe_1_6_1_net3351), .RN(npu_inst_pe_1_6_1_n8), .Q(
        npu_inst_int_data_res_6__1__7_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_1_n100), 
        .CK(npu_inst_pe_1_6_1_net3351), .RN(npu_inst_pe_1_6_1_n8), .Q(
        npu_inst_int_data_res_6__1__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_weight_reg_0_ ( .D(npu_inst_n91), .CK(
        npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n8), .Q(
        npu_inst_pe_1_6_1_int_q_weight_0_), .QN(npu_inst_pe_1_6_1_n27) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_weight_reg_1_ ( .D(npu_inst_n97), .CK(
        npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n8), .Q(
        npu_inst_pe_1_6_1_int_q_weight_1_), .QN(npu_inst_pe_1_6_1_n26) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_1_n112), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n8), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_1_n106), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n8), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_1_n111), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_1_n105), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_1_n110), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_1_n104), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_1_n109), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_1_n103), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_1_n108), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_1_n102), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_1_n107), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_1_n101), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_1_n86), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_1_n87), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n9), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_1_n88), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_1_n89), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_1_n90), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_1_n91), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_1_n92), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_1_n93), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_1_n94), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_1_n95), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_1_n96), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_1_n97), 
        .CK(npu_inst_pe_1_6_1_net3357), .RN(npu_inst_pe_1_6_1_n10), .Q(
        npu_inst_pe_1_6_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_1_net3351) );
  CLKGATETST_X1 npu_inst_pe_1_6_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n44), .SE(1'b0), .GCK(npu_inst_pe_1_6_1_net3357) );
  MUX2_X1 npu_inst_pe_1_6_2_U153 ( .A(npu_inst_pe_1_6_2_n31), .B(
        npu_inst_pe_1_6_2_n28), .S(npu_inst_pe_1_6_2_n7), .Z(
        npu_inst_pe_1_6_2_N93) );
  MUX2_X1 npu_inst_pe_1_6_2_U152 ( .A(npu_inst_pe_1_6_2_n30), .B(
        npu_inst_pe_1_6_2_n29), .S(npu_inst_pe_1_6_2_n5), .Z(
        npu_inst_pe_1_6_2_n31) );
  MUX2_X1 npu_inst_pe_1_6_2_U151 ( .A(npu_inst_pe_1_6_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_2_n3), .Z(
        npu_inst_pe_1_6_2_n30) );
  MUX2_X1 npu_inst_pe_1_6_2_U150 ( .A(npu_inst_pe_1_6_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_2_n3), .Z(
        npu_inst_pe_1_6_2_n29) );
  MUX2_X1 npu_inst_pe_1_6_2_U149 ( .A(npu_inst_pe_1_6_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_2_n3), .Z(
        npu_inst_pe_1_6_2_n28) );
  MUX2_X1 npu_inst_pe_1_6_2_U148 ( .A(npu_inst_pe_1_6_2_n25), .B(
        npu_inst_pe_1_6_2_n22), .S(npu_inst_pe_1_6_2_n7), .Z(
        npu_inst_pe_1_6_2_N94) );
  MUX2_X1 npu_inst_pe_1_6_2_U147 ( .A(npu_inst_pe_1_6_2_n24), .B(
        npu_inst_pe_1_6_2_n23), .S(npu_inst_pe_1_6_2_n5), .Z(
        npu_inst_pe_1_6_2_n25) );
  MUX2_X1 npu_inst_pe_1_6_2_U146 ( .A(npu_inst_pe_1_6_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_2_n3), .Z(
        npu_inst_pe_1_6_2_n24) );
  MUX2_X1 npu_inst_pe_1_6_2_U145 ( .A(npu_inst_pe_1_6_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_2_n3), .Z(
        npu_inst_pe_1_6_2_n23) );
  MUX2_X1 npu_inst_pe_1_6_2_U144 ( .A(npu_inst_pe_1_6_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_2_n3), .Z(
        npu_inst_pe_1_6_2_n22) );
  MUX2_X1 npu_inst_pe_1_6_2_U143 ( .A(npu_inst_pe_1_6_2_n21), .B(
        npu_inst_pe_1_6_2_n18), .S(npu_inst_pe_1_6_2_n7), .Z(
        npu_inst_int_data_x_6__2__1_) );
  MUX2_X1 npu_inst_pe_1_6_2_U142 ( .A(npu_inst_pe_1_6_2_n20), .B(
        npu_inst_pe_1_6_2_n19), .S(npu_inst_pe_1_6_2_n5), .Z(
        npu_inst_pe_1_6_2_n21) );
  MUX2_X1 npu_inst_pe_1_6_2_U141 ( .A(npu_inst_pe_1_6_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_2_n3), .Z(
        npu_inst_pe_1_6_2_n20) );
  MUX2_X1 npu_inst_pe_1_6_2_U140 ( .A(npu_inst_pe_1_6_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_2_n3), .Z(
        npu_inst_pe_1_6_2_n19) );
  MUX2_X1 npu_inst_pe_1_6_2_U139 ( .A(npu_inst_pe_1_6_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_2_n3), .Z(
        npu_inst_pe_1_6_2_n18) );
  MUX2_X1 npu_inst_pe_1_6_2_U138 ( .A(npu_inst_pe_1_6_2_n17), .B(
        npu_inst_pe_1_6_2_n14), .S(npu_inst_pe_1_6_2_n7), .Z(
        npu_inst_int_data_x_6__2__0_) );
  MUX2_X1 npu_inst_pe_1_6_2_U137 ( .A(npu_inst_pe_1_6_2_n16), .B(
        npu_inst_pe_1_6_2_n15), .S(npu_inst_pe_1_6_2_n5), .Z(
        npu_inst_pe_1_6_2_n17) );
  MUX2_X1 npu_inst_pe_1_6_2_U136 ( .A(npu_inst_pe_1_6_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_2_n3), .Z(
        npu_inst_pe_1_6_2_n16) );
  MUX2_X1 npu_inst_pe_1_6_2_U135 ( .A(npu_inst_pe_1_6_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_2_n3), .Z(
        npu_inst_pe_1_6_2_n15) );
  MUX2_X1 npu_inst_pe_1_6_2_U134 ( .A(npu_inst_pe_1_6_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_2_n3), .Z(
        npu_inst_pe_1_6_2_n14) );
  XOR2_X1 npu_inst_pe_1_6_2_U133 ( .A(npu_inst_pe_1_6_2_int_data_0_), .B(
        npu_inst_int_data_res_6__2__0_), .Z(npu_inst_pe_1_6_2_N73) );
  AND2_X1 npu_inst_pe_1_6_2_U132 ( .A1(npu_inst_int_data_res_6__2__0_), .A2(
        npu_inst_pe_1_6_2_int_data_0_), .ZN(npu_inst_pe_1_6_2_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_2_U131 ( .A(npu_inst_int_data_res_6__2__0_), .B(
        npu_inst_pe_1_6_2_n12), .ZN(npu_inst_pe_1_6_2_N65) );
  OR2_X1 npu_inst_pe_1_6_2_U130 ( .A1(npu_inst_pe_1_6_2_n12), .A2(
        npu_inst_int_data_res_6__2__0_), .ZN(npu_inst_pe_1_6_2_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_2_U129 ( .A(npu_inst_int_data_res_6__2__2_), .B(
        npu_inst_pe_1_6_2_add_79_carry_2_), .Z(npu_inst_pe_1_6_2_N75) );
  AND2_X1 npu_inst_pe_1_6_2_U128 ( .A1(npu_inst_pe_1_6_2_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_6__2__2_), .ZN(
        npu_inst_pe_1_6_2_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_2_U127 ( .A(npu_inst_int_data_res_6__2__3_), .B(
        npu_inst_pe_1_6_2_add_79_carry_3_), .Z(npu_inst_pe_1_6_2_N76) );
  AND2_X1 npu_inst_pe_1_6_2_U126 ( .A1(npu_inst_pe_1_6_2_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_6__2__3_), .ZN(
        npu_inst_pe_1_6_2_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_2_U125 ( .A(npu_inst_int_data_res_6__2__4_), .B(
        npu_inst_pe_1_6_2_add_79_carry_4_), .Z(npu_inst_pe_1_6_2_N77) );
  AND2_X1 npu_inst_pe_1_6_2_U124 ( .A1(npu_inst_pe_1_6_2_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_6__2__4_), .ZN(
        npu_inst_pe_1_6_2_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_2_U123 ( .A(npu_inst_int_data_res_6__2__5_), .B(
        npu_inst_pe_1_6_2_add_79_carry_5_), .Z(npu_inst_pe_1_6_2_N78) );
  AND2_X1 npu_inst_pe_1_6_2_U122 ( .A1(npu_inst_pe_1_6_2_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_6__2__5_), .ZN(
        npu_inst_pe_1_6_2_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_2_U121 ( .A(npu_inst_int_data_res_6__2__6_), .B(
        npu_inst_pe_1_6_2_add_79_carry_6_), .Z(npu_inst_pe_1_6_2_N79) );
  AND2_X1 npu_inst_pe_1_6_2_U120 ( .A1(npu_inst_pe_1_6_2_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_6__2__6_), .ZN(
        npu_inst_pe_1_6_2_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_2_U119 ( .A(npu_inst_int_data_res_6__2__7_), .B(
        npu_inst_pe_1_6_2_add_79_carry_7_), .Z(npu_inst_pe_1_6_2_N80) );
  XNOR2_X1 npu_inst_pe_1_6_2_U118 ( .A(npu_inst_pe_1_6_2_sub_77_carry_2_), .B(
        npu_inst_int_data_res_6__2__2_), .ZN(npu_inst_pe_1_6_2_N67) );
  OR2_X1 npu_inst_pe_1_6_2_U117 ( .A1(npu_inst_int_data_res_6__2__2_), .A2(
        npu_inst_pe_1_6_2_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_6_2_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_2_U116 ( .A(npu_inst_pe_1_6_2_sub_77_carry_3_), .B(
        npu_inst_int_data_res_6__2__3_), .ZN(npu_inst_pe_1_6_2_N68) );
  OR2_X1 npu_inst_pe_1_6_2_U115 ( .A1(npu_inst_int_data_res_6__2__3_), .A2(
        npu_inst_pe_1_6_2_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_6_2_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_2_U114 ( .A(npu_inst_pe_1_6_2_sub_77_carry_4_), .B(
        npu_inst_int_data_res_6__2__4_), .ZN(npu_inst_pe_1_6_2_N69) );
  OR2_X1 npu_inst_pe_1_6_2_U113 ( .A1(npu_inst_int_data_res_6__2__4_), .A2(
        npu_inst_pe_1_6_2_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_6_2_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_2_U112 ( .A(npu_inst_pe_1_6_2_sub_77_carry_5_), .B(
        npu_inst_int_data_res_6__2__5_), .ZN(npu_inst_pe_1_6_2_N70) );
  OR2_X1 npu_inst_pe_1_6_2_U111 ( .A1(npu_inst_int_data_res_6__2__5_), .A2(
        npu_inst_pe_1_6_2_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_6_2_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_2_U110 ( .A(npu_inst_pe_1_6_2_sub_77_carry_6_), .B(
        npu_inst_int_data_res_6__2__6_), .ZN(npu_inst_pe_1_6_2_N71) );
  OR2_X1 npu_inst_pe_1_6_2_U109 ( .A1(npu_inst_int_data_res_6__2__6_), .A2(
        npu_inst_pe_1_6_2_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_6_2_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_2_U108 ( .A(npu_inst_int_data_res_6__2__7_), .B(
        npu_inst_pe_1_6_2_sub_77_carry_7_), .ZN(npu_inst_pe_1_6_2_N72) );
  INV_X1 npu_inst_pe_1_6_2_U107 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_6_2_n6)
         );
  INV_X1 npu_inst_pe_1_6_2_U106 ( .A(npu_inst_pe_1_6_2_n6), .ZN(
        npu_inst_pe_1_6_2_n5) );
  INV_X1 npu_inst_pe_1_6_2_U105 ( .A(npu_inst_n35), .ZN(npu_inst_pe_1_6_2_n2)
         );
  AOI22_X1 npu_inst_pe_1_6_2_U104 ( .A1(npu_inst_int_data_y_7__2__0_), .A2(
        npu_inst_pe_1_6_2_n58), .B1(npu_inst_pe_1_6_2_n118), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_2_n57) );
  INV_X1 npu_inst_pe_1_6_2_U103 ( .A(npu_inst_pe_1_6_2_n57), .ZN(
        npu_inst_pe_1_6_2_n107) );
  AOI22_X1 npu_inst_pe_1_6_2_U102 ( .A1(npu_inst_int_data_y_7__2__0_), .A2(
        npu_inst_pe_1_6_2_n54), .B1(npu_inst_pe_1_6_2_n117), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_2_n53) );
  INV_X1 npu_inst_pe_1_6_2_U99 ( .A(npu_inst_pe_1_6_2_n53), .ZN(
        npu_inst_pe_1_6_2_n108) );
  AOI22_X1 npu_inst_pe_1_6_2_U98 ( .A1(npu_inst_int_data_y_7__2__0_), .A2(
        npu_inst_pe_1_6_2_n50), .B1(npu_inst_pe_1_6_2_n116), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_2_n49) );
  INV_X1 npu_inst_pe_1_6_2_U97 ( .A(npu_inst_pe_1_6_2_n49), .ZN(
        npu_inst_pe_1_6_2_n109) );
  AOI22_X1 npu_inst_pe_1_6_2_U96 ( .A1(npu_inst_int_data_y_7__2__0_), .A2(
        npu_inst_pe_1_6_2_n46), .B1(npu_inst_pe_1_6_2_n115), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_2_n45) );
  INV_X1 npu_inst_pe_1_6_2_U95 ( .A(npu_inst_pe_1_6_2_n45), .ZN(
        npu_inst_pe_1_6_2_n110) );
  AOI22_X1 npu_inst_pe_1_6_2_U94 ( .A1(npu_inst_int_data_y_7__2__0_), .A2(
        npu_inst_pe_1_6_2_n42), .B1(npu_inst_pe_1_6_2_n114), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_2_n41) );
  INV_X1 npu_inst_pe_1_6_2_U93 ( .A(npu_inst_pe_1_6_2_n41), .ZN(
        npu_inst_pe_1_6_2_n111) );
  AOI22_X1 npu_inst_pe_1_6_2_U92 ( .A1(npu_inst_int_data_y_7__2__1_), .A2(
        npu_inst_pe_1_6_2_n58), .B1(npu_inst_pe_1_6_2_n118), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_2_n59) );
  INV_X1 npu_inst_pe_1_6_2_U91 ( .A(npu_inst_pe_1_6_2_n59), .ZN(
        npu_inst_pe_1_6_2_n101) );
  AOI22_X1 npu_inst_pe_1_6_2_U90 ( .A1(npu_inst_int_data_y_7__2__1_), .A2(
        npu_inst_pe_1_6_2_n54), .B1(npu_inst_pe_1_6_2_n117), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_2_n55) );
  INV_X1 npu_inst_pe_1_6_2_U89 ( .A(npu_inst_pe_1_6_2_n55), .ZN(
        npu_inst_pe_1_6_2_n102) );
  AOI22_X1 npu_inst_pe_1_6_2_U88 ( .A1(npu_inst_int_data_y_7__2__1_), .A2(
        npu_inst_pe_1_6_2_n50), .B1(npu_inst_pe_1_6_2_n116), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_2_n51) );
  INV_X1 npu_inst_pe_1_6_2_U87 ( .A(npu_inst_pe_1_6_2_n51), .ZN(
        npu_inst_pe_1_6_2_n103) );
  AOI22_X1 npu_inst_pe_1_6_2_U86 ( .A1(npu_inst_int_data_y_7__2__1_), .A2(
        npu_inst_pe_1_6_2_n46), .B1(npu_inst_pe_1_6_2_n115), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_2_n47) );
  INV_X1 npu_inst_pe_1_6_2_U85 ( .A(npu_inst_pe_1_6_2_n47), .ZN(
        npu_inst_pe_1_6_2_n104) );
  AOI22_X1 npu_inst_pe_1_6_2_U84 ( .A1(npu_inst_int_data_y_7__2__1_), .A2(
        npu_inst_pe_1_6_2_n42), .B1(npu_inst_pe_1_6_2_n114), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_2_n43) );
  INV_X1 npu_inst_pe_1_6_2_U83 ( .A(npu_inst_pe_1_6_2_n43), .ZN(
        npu_inst_pe_1_6_2_n105) );
  AOI22_X1 npu_inst_pe_1_6_2_U82 ( .A1(npu_inst_pe_1_6_2_n38), .A2(
        npu_inst_int_data_y_7__2__1_), .B1(npu_inst_pe_1_6_2_n113), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_2_n39) );
  INV_X1 npu_inst_pe_1_6_2_U81 ( .A(npu_inst_pe_1_6_2_n39), .ZN(
        npu_inst_pe_1_6_2_n106) );
  AND2_X1 npu_inst_pe_1_6_2_U80 ( .A1(npu_inst_pe_1_6_2_N93), .A2(npu_inst_n35), .ZN(npu_inst_int_data_y_6__2__0_) );
  NAND2_X1 npu_inst_pe_1_6_2_U79 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_2_n60), .ZN(npu_inst_pe_1_6_2_n74) );
  OAI21_X1 npu_inst_pe_1_6_2_U78 ( .B1(npu_inst_pe_1_6_2_n63), .B2(
        npu_inst_pe_1_6_2_n60), .A(npu_inst_pe_1_6_2_n74), .ZN(
        npu_inst_pe_1_6_2_n97) );
  NAND2_X1 npu_inst_pe_1_6_2_U77 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_2_n60), .ZN(npu_inst_pe_1_6_2_n73) );
  OAI21_X1 npu_inst_pe_1_6_2_U76 ( .B1(npu_inst_pe_1_6_2_n61), .B2(
        npu_inst_pe_1_6_2_n60), .A(npu_inst_pe_1_6_2_n73), .ZN(
        npu_inst_pe_1_6_2_n96) );
  NAND2_X1 npu_inst_pe_1_6_2_U75 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_2_n56), .ZN(npu_inst_pe_1_6_2_n72) );
  OAI21_X1 npu_inst_pe_1_6_2_U74 ( .B1(npu_inst_pe_1_6_2_n63), .B2(
        npu_inst_pe_1_6_2_n56), .A(npu_inst_pe_1_6_2_n72), .ZN(
        npu_inst_pe_1_6_2_n95) );
  NAND2_X1 npu_inst_pe_1_6_2_U73 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_2_n56), .ZN(npu_inst_pe_1_6_2_n71) );
  OAI21_X1 npu_inst_pe_1_6_2_U72 ( .B1(npu_inst_pe_1_6_2_n61), .B2(
        npu_inst_pe_1_6_2_n56), .A(npu_inst_pe_1_6_2_n71), .ZN(
        npu_inst_pe_1_6_2_n94) );
  NAND2_X1 npu_inst_pe_1_6_2_U71 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_2_n52), .ZN(npu_inst_pe_1_6_2_n70) );
  OAI21_X1 npu_inst_pe_1_6_2_U70 ( .B1(npu_inst_pe_1_6_2_n63), .B2(
        npu_inst_pe_1_6_2_n52), .A(npu_inst_pe_1_6_2_n70), .ZN(
        npu_inst_pe_1_6_2_n93) );
  NAND2_X1 npu_inst_pe_1_6_2_U69 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_2_n52), .ZN(npu_inst_pe_1_6_2_n69) );
  OAI21_X1 npu_inst_pe_1_6_2_U68 ( .B1(npu_inst_pe_1_6_2_n61), .B2(
        npu_inst_pe_1_6_2_n52), .A(npu_inst_pe_1_6_2_n69), .ZN(
        npu_inst_pe_1_6_2_n92) );
  NAND2_X1 npu_inst_pe_1_6_2_U67 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_2_n48), .ZN(npu_inst_pe_1_6_2_n68) );
  OAI21_X1 npu_inst_pe_1_6_2_U66 ( .B1(npu_inst_pe_1_6_2_n63), .B2(
        npu_inst_pe_1_6_2_n48), .A(npu_inst_pe_1_6_2_n68), .ZN(
        npu_inst_pe_1_6_2_n91) );
  NAND2_X1 npu_inst_pe_1_6_2_U65 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_2_n48), .ZN(npu_inst_pe_1_6_2_n67) );
  OAI21_X1 npu_inst_pe_1_6_2_U64 ( .B1(npu_inst_pe_1_6_2_n61), .B2(
        npu_inst_pe_1_6_2_n48), .A(npu_inst_pe_1_6_2_n67), .ZN(
        npu_inst_pe_1_6_2_n90) );
  NAND2_X1 npu_inst_pe_1_6_2_U63 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_2_n44), .ZN(npu_inst_pe_1_6_2_n66) );
  OAI21_X1 npu_inst_pe_1_6_2_U62 ( .B1(npu_inst_pe_1_6_2_n63), .B2(
        npu_inst_pe_1_6_2_n44), .A(npu_inst_pe_1_6_2_n66), .ZN(
        npu_inst_pe_1_6_2_n89) );
  NAND2_X1 npu_inst_pe_1_6_2_U61 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_2_n44), .ZN(npu_inst_pe_1_6_2_n65) );
  OAI21_X1 npu_inst_pe_1_6_2_U60 ( .B1(npu_inst_pe_1_6_2_n61), .B2(
        npu_inst_pe_1_6_2_n44), .A(npu_inst_pe_1_6_2_n65), .ZN(
        npu_inst_pe_1_6_2_n88) );
  NAND2_X1 npu_inst_pe_1_6_2_U59 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_2_n40), .ZN(npu_inst_pe_1_6_2_n64) );
  OAI21_X1 npu_inst_pe_1_6_2_U58 ( .B1(npu_inst_pe_1_6_2_n63), .B2(
        npu_inst_pe_1_6_2_n40), .A(npu_inst_pe_1_6_2_n64), .ZN(
        npu_inst_pe_1_6_2_n87) );
  NAND2_X1 npu_inst_pe_1_6_2_U57 ( .A1(npu_inst_pe_1_6_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_2_n40), .ZN(npu_inst_pe_1_6_2_n62) );
  OAI21_X1 npu_inst_pe_1_6_2_U56 ( .B1(npu_inst_pe_1_6_2_n61), .B2(
        npu_inst_pe_1_6_2_n40), .A(npu_inst_pe_1_6_2_n62), .ZN(
        npu_inst_pe_1_6_2_n86) );
  AOI22_X1 npu_inst_pe_1_6_2_U55 ( .A1(npu_inst_pe_1_6_2_n38), .A2(
        npu_inst_int_data_y_7__2__0_), .B1(npu_inst_pe_1_6_2_n113), .B2(
        npu_inst_pe_1_6_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_2_n37) );
  INV_X1 npu_inst_pe_1_6_2_U54 ( .A(npu_inst_pe_1_6_2_n37), .ZN(
        npu_inst_pe_1_6_2_n112) );
  AND2_X1 npu_inst_pe_1_6_2_U53 ( .A1(npu_inst_n35), .A2(npu_inst_pe_1_6_2_N94), .ZN(npu_inst_int_data_y_6__2__1_) );
  AOI222_X1 npu_inst_pe_1_6_2_U52 ( .A1(npu_inst_int_data_res_7__2__0_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N73), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N65), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n84) );
  INV_X1 npu_inst_pe_1_6_2_U51 ( .A(npu_inst_pe_1_6_2_n84), .ZN(
        npu_inst_pe_1_6_2_n100) );
  AOI222_X1 npu_inst_pe_1_6_2_U50 ( .A1(npu_inst_pe_1_6_2_n1), .A2(
        npu_inst_int_data_res_7__2__7_), .B1(npu_inst_pe_1_6_2_N80), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N72), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n75) );
  INV_X1 npu_inst_pe_1_6_2_U49 ( .A(npu_inst_pe_1_6_2_n75), .ZN(
        npu_inst_pe_1_6_2_n32) );
  AOI222_X1 npu_inst_pe_1_6_2_U48 ( .A1(npu_inst_int_data_res_7__2__1_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N74), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N66), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n83) );
  INV_X1 npu_inst_pe_1_6_2_U47 ( .A(npu_inst_pe_1_6_2_n83), .ZN(
        npu_inst_pe_1_6_2_n99) );
  AOI222_X1 npu_inst_pe_1_6_2_U46 ( .A1(npu_inst_int_data_res_7__2__3_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N76), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N68), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n81) );
  INV_X1 npu_inst_pe_1_6_2_U45 ( .A(npu_inst_pe_1_6_2_n81), .ZN(
        npu_inst_pe_1_6_2_n36) );
  AOI222_X1 npu_inst_pe_1_6_2_U44 ( .A1(npu_inst_int_data_res_7__2__4_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N77), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N69), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n80) );
  INV_X1 npu_inst_pe_1_6_2_U43 ( .A(npu_inst_pe_1_6_2_n80), .ZN(
        npu_inst_pe_1_6_2_n35) );
  AOI222_X1 npu_inst_pe_1_6_2_U42 ( .A1(npu_inst_int_data_res_7__2__5_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N78), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N70), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n79) );
  INV_X1 npu_inst_pe_1_6_2_U41 ( .A(npu_inst_pe_1_6_2_n79), .ZN(
        npu_inst_pe_1_6_2_n34) );
  AOI222_X1 npu_inst_pe_1_6_2_U40 ( .A1(npu_inst_int_data_res_7__2__6_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N79), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N71), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n78) );
  INV_X1 npu_inst_pe_1_6_2_U39 ( .A(npu_inst_pe_1_6_2_n78), .ZN(
        npu_inst_pe_1_6_2_n33) );
  AND2_X1 npu_inst_pe_1_6_2_U38 ( .A1(npu_inst_int_data_x_6__2__1_), .A2(
        npu_inst_pe_1_6_2_int_q_weight_1_), .ZN(npu_inst_pe_1_6_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_2_U37 ( .A1(npu_inst_int_data_x_6__2__0_), .A2(
        npu_inst_pe_1_6_2_int_q_weight_1_), .ZN(npu_inst_pe_1_6_2_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_6_2_U36 ( .A(npu_inst_pe_1_6_2_int_data_1_), .ZN(
        npu_inst_pe_1_6_2_n13) );
  NOR3_X1 npu_inst_pe_1_6_2_U35 ( .A1(npu_inst_pe_1_6_2_n26), .A2(npu_inst_n35), .A3(npu_inst_int_ckg[13]), .ZN(npu_inst_pe_1_6_2_n85) );
  OR2_X1 npu_inst_pe_1_6_2_U34 ( .A1(npu_inst_pe_1_6_2_n85), .A2(
        npu_inst_pe_1_6_2_n1), .ZN(npu_inst_pe_1_6_2_N84) );
  AOI222_X1 npu_inst_pe_1_6_2_U33 ( .A1(npu_inst_int_data_res_7__2__2_), .A2(
        npu_inst_pe_1_6_2_n1), .B1(npu_inst_pe_1_6_2_N75), .B2(
        npu_inst_pe_1_6_2_n76), .C1(npu_inst_pe_1_6_2_N67), .C2(
        npu_inst_pe_1_6_2_n77), .ZN(npu_inst_pe_1_6_2_n82) );
  INV_X1 npu_inst_pe_1_6_2_U32 ( .A(npu_inst_pe_1_6_2_n82), .ZN(
        npu_inst_pe_1_6_2_n98) );
  AOI22_X1 npu_inst_pe_1_6_2_U31 ( .A1(npu_inst_n35), .A2(
        npu_inst_int_data_y_7__2__1_), .B1(npu_inst_pe_1_6_2_n2), .B2(
        npu_inst_int_data_x_6__3__1_), .ZN(npu_inst_pe_1_6_2_n63) );
  AOI22_X1 npu_inst_pe_1_6_2_U30 ( .A1(npu_inst_n35), .A2(
        npu_inst_int_data_y_7__2__0_), .B1(npu_inst_pe_1_6_2_n2), .B2(
        npu_inst_int_data_x_6__3__0_), .ZN(npu_inst_pe_1_6_2_n61) );
  INV_X1 npu_inst_pe_1_6_2_U29 ( .A(npu_inst_pe_1_6_2_int_data_0_), .ZN(
        npu_inst_pe_1_6_2_n12) );
  INV_X1 npu_inst_pe_1_6_2_U28 ( .A(npu_inst_n50), .ZN(npu_inst_pe_1_6_2_n4)
         );
  OR3_X1 npu_inst_pe_1_6_2_U27 ( .A1(npu_inst_pe_1_6_2_n5), .A2(
        npu_inst_pe_1_6_2_n7), .A3(npu_inst_pe_1_6_2_n4), .ZN(
        npu_inst_pe_1_6_2_n56) );
  OR3_X1 npu_inst_pe_1_6_2_U26 ( .A1(npu_inst_pe_1_6_2_n4), .A2(
        npu_inst_pe_1_6_2_n7), .A3(npu_inst_pe_1_6_2_n6), .ZN(
        npu_inst_pe_1_6_2_n48) );
  INV_X1 npu_inst_pe_1_6_2_U25 ( .A(npu_inst_pe_1_6_2_n4), .ZN(
        npu_inst_pe_1_6_2_n3) );
  OR3_X1 npu_inst_pe_1_6_2_U24 ( .A1(npu_inst_pe_1_6_2_n3), .A2(
        npu_inst_pe_1_6_2_n7), .A3(npu_inst_pe_1_6_2_n6), .ZN(
        npu_inst_pe_1_6_2_n52) );
  OR3_X1 npu_inst_pe_1_6_2_U23 ( .A1(npu_inst_pe_1_6_2_n5), .A2(
        npu_inst_pe_1_6_2_n7), .A3(npu_inst_pe_1_6_2_n3), .ZN(
        npu_inst_pe_1_6_2_n60) );
  BUF_X1 npu_inst_pe_1_6_2_U22 ( .A(npu_inst_n15), .Z(npu_inst_pe_1_6_2_n1) );
  NOR2_X1 npu_inst_pe_1_6_2_U21 ( .A1(npu_inst_pe_1_6_2_n60), .A2(
        npu_inst_pe_1_6_2_n2), .ZN(npu_inst_pe_1_6_2_n58) );
  NOR2_X1 npu_inst_pe_1_6_2_U20 ( .A1(npu_inst_pe_1_6_2_n56), .A2(
        npu_inst_pe_1_6_2_n2), .ZN(npu_inst_pe_1_6_2_n54) );
  NOR2_X1 npu_inst_pe_1_6_2_U19 ( .A1(npu_inst_pe_1_6_2_n52), .A2(
        npu_inst_pe_1_6_2_n2), .ZN(npu_inst_pe_1_6_2_n50) );
  NOR2_X1 npu_inst_pe_1_6_2_U18 ( .A1(npu_inst_pe_1_6_2_n48), .A2(
        npu_inst_pe_1_6_2_n2), .ZN(npu_inst_pe_1_6_2_n46) );
  NOR2_X1 npu_inst_pe_1_6_2_U17 ( .A1(npu_inst_pe_1_6_2_n40), .A2(
        npu_inst_pe_1_6_2_n2), .ZN(npu_inst_pe_1_6_2_n38) );
  NOR2_X1 npu_inst_pe_1_6_2_U16 ( .A1(npu_inst_pe_1_6_2_n44), .A2(
        npu_inst_pe_1_6_2_n2), .ZN(npu_inst_pe_1_6_2_n42) );
  BUF_X1 npu_inst_pe_1_6_2_U15 ( .A(npu_inst_n77), .Z(npu_inst_pe_1_6_2_n7) );
  INV_X1 npu_inst_pe_1_6_2_U14 ( .A(npu_inst_n105), .ZN(npu_inst_pe_1_6_2_n11)
         );
  INV_X1 npu_inst_pe_1_6_2_U13 ( .A(npu_inst_pe_1_6_2_n38), .ZN(
        npu_inst_pe_1_6_2_n113) );
  INV_X1 npu_inst_pe_1_6_2_U12 ( .A(npu_inst_pe_1_6_2_n58), .ZN(
        npu_inst_pe_1_6_2_n118) );
  INV_X1 npu_inst_pe_1_6_2_U11 ( .A(npu_inst_pe_1_6_2_n54), .ZN(
        npu_inst_pe_1_6_2_n117) );
  INV_X1 npu_inst_pe_1_6_2_U10 ( .A(npu_inst_pe_1_6_2_n50), .ZN(
        npu_inst_pe_1_6_2_n116) );
  INV_X1 npu_inst_pe_1_6_2_U9 ( .A(npu_inst_pe_1_6_2_n46), .ZN(
        npu_inst_pe_1_6_2_n115) );
  INV_X1 npu_inst_pe_1_6_2_U8 ( .A(npu_inst_pe_1_6_2_n42), .ZN(
        npu_inst_pe_1_6_2_n114) );
  BUF_X1 npu_inst_pe_1_6_2_U7 ( .A(npu_inst_pe_1_6_2_n11), .Z(
        npu_inst_pe_1_6_2_n10) );
  BUF_X1 npu_inst_pe_1_6_2_U6 ( .A(npu_inst_pe_1_6_2_n11), .Z(
        npu_inst_pe_1_6_2_n9) );
  BUF_X1 npu_inst_pe_1_6_2_U5 ( .A(npu_inst_pe_1_6_2_n11), .Z(
        npu_inst_pe_1_6_2_n8) );
  NOR2_X1 npu_inst_pe_1_6_2_U4 ( .A1(npu_inst_pe_1_6_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_2_n1), .ZN(npu_inst_pe_1_6_2_n76) );
  NOR2_X1 npu_inst_pe_1_6_2_U3 ( .A1(npu_inst_pe_1_6_2_n27), .A2(
        npu_inst_pe_1_6_2_n1), .ZN(npu_inst_pe_1_6_2_n77) );
  FA_X1 npu_inst_pe_1_6_2_sub_77_U2_1 ( .A(npu_inst_int_data_res_6__2__1_), 
        .B(npu_inst_pe_1_6_2_n13), .CI(npu_inst_pe_1_6_2_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_6_2_sub_77_carry_2_), .S(npu_inst_pe_1_6_2_N66) );
  FA_X1 npu_inst_pe_1_6_2_add_79_U1_1 ( .A(npu_inst_int_data_res_6__2__1_), 
        .B(npu_inst_pe_1_6_2_int_data_1_), .CI(
        npu_inst_pe_1_6_2_add_79_carry_1_), .CO(
        npu_inst_pe_1_6_2_add_79_carry_2_), .S(npu_inst_pe_1_6_2_N74) );
  NAND3_X1 npu_inst_pe_1_6_2_U101 ( .A1(npu_inst_pe_1_6_2_n4), .A2(
        npu_inst_pe_1_6_2_n6), .A3(npu_inst_pe_1_6_2_n7), .ZN(
        npu_inst_pe_1_6_2_n44) );
  NAND3_X1 npu_inst_pe_1_6_2_U100 ( .A1(npu_inst_pe_1_6_2_n3), .A2(
        npu_inst_pe_1_6_2_n6), .A3(npu_inst_pe_1_6_2_n7), .ZN(
        npu_inst_pe_1_6_2_n40) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_2_n33), .CK(
        npu_inst_pe_1_6_2_net3328), .RN(npu_inst_pe_1_6_2_n8), .Q(
        npu_inst_int_data_res_6__2__6_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_2_n34), .CK(
        npu_inst_pe_1_6_2_net3328), .RN(npu_inst_pe_1_6_2_n8), .Q(
        npu_inst_int_data_res_6__2__5_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_2_n35), .CK(
        npu_inst_pe_1_6_2_net3328), .RN(npu_inst_pe_1_6_2_n8), .Q(
        npu_inst_int_data_res_6__2__4_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_2_n36), .CK(
        npu_inst_pe_1_6_2_net3328), .RN(npu_inst_pe_1_6_2_n8), .Q(
        npu_inst_int_data_res_6__2__3_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_2_n98), .CK(
        npu_inst_pe_1_6_2_net3328), .RN(npu_inst_pe_1_6_2_n8), .Q(
        npu_inst_int_data_res_6__2__2_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_2_n99), .CK(
        npu_inst_pe_1_6_2_net3328), .RN(npu_inst_pe_1_6_2_n8), .Q(
        npu_inst_int_data_res_6__2__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_2_n32), .CK(
        npu_inst_pe_1_6_2_net3328), .RN(npu_inst_pe_1_6_2_n8), .Q(
        npu_inst_int_data_res_6__2__7_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_2_n100), 
        .CK(npu_inst_pe_1_6_2_net3328), .RN(npu_inst_pe_1_6_2_n8), .Q(
        npu_inst_int_data_res_6__2__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_weight_reg_0_ ( .D(npu_inst_n91), .CK(
        npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n8), .Q(
        npu_inst_pe_1_6_2_int_q_weight_0_), .QN(npu_inst_pe_1_6_2_n27) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_weight_reg_1_ ( .D(npu_inst_n97), .CK(
        npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n8), .Q(
        npu_inst_pe_1_6_2_int_q_weight_1_), .QN(npu_inst_pe_1_6_2_n26) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_2_n112), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n8), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_2_n106), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n8), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_2_n111), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_2_n105), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_2_n110), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_2_n104), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_2_n109), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_2_n103), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_2_n108), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_2_n102), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_2_n107), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_2_n101), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_2_n86), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_2_n87), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n9), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_2_n88), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_2_n89), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_2_n90), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_2_n91), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_2_n92), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_2_n93), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_2_n94), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_2_n95), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_2_n96), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_2_n97), 
        .CK(npu_inst_pe_1_6_2_net3334), .RN(npu_inst_pe_1_6_2_n10), .Q(
        npu_inst_pe_1_6_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_2_net3328) );
  CLKGATETST_X1 npu_inst_pe_1_6_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n44), .SE(1'b0), .GCK(npu_inst_pe_1_6_2_net3334) );
  MUX2_X1 npu_inst_pe_1_6_3_U153 ( .A(npu_inst_pe_1_6_3_n31), .B(
        npu_inst_pe_1_6_3_n28), .S(npu_inst_pe_1_6_3_n7), .Z(
        npu_inst_pe_1_6_3_N93) );
  MUX2_X1 npu_inst_pe_1_6_3_U152 ( .A(npu_inst_pe_1_6_3_n30), .B(
        npu_inst_pe_1_6_3_n29), .S(npu_inst_pe_1_6_3_n5), .Z(
        npu_inst_pe_1_6_3_n31) );
  MUX2_X1 npu_inst_pe_1_6_3_U151 ( .A(npu_inst_pe_1_6_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_3_n3), .Z(
        npu_inst_pe_1_6_3_n30) );
  MUX2_X1 npu_inst_pe_1_6_3_U150 ( .A(npu_inst_pe_1_6_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_3_n3), .Z(
        npu_inst_pe_1_6_3_n29) );
  MUX2_X1 npu_inst_pe_1_6_3_U149 ( .A(npu_inst_pe_1_6_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_3_n3), .Z(
        npu_inst_pe_1_6_3_n28) );
  MUX2_X1 npu_inst_pe_1_6_3_U148 ( .A(npu_inst_pe_1_6_3_n25), .B(
        npu_inst_pe_1_6_3_n22), .S(npu_inst_pe_1_6_3_n7), .Z(
        npu_inst_pe_1_6_3_N94) );
  MUX2_X1 npu_inst_pe_1_6_3_U147 ( .A(npu_inst_pe_1_6_3_n24), .B(
        npu_inst_pe_1_6_3_n23), .S(npu_inst_pe_1_6_3_n5), .Z(
        npu_inst_pe_1_6_3_n25) );
  MUX2_X1 npu_inst_pe_1_6_3_U146 ( .A(npu_inst_pe_1_6_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_3_n3), .Z(
        npu_inst_pe_1_6_3_n24) );
  MUX2_X1 npu_inst_pe_1_6_3_U145 ( .A(npu_inst_pe_1_6_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_3_n3), .Z(
        npu_inst_pe_1_6_3_n23) );
  MUX2_X1 npu_inst_pe_1_6_3_U144 ( .A(npu_inst_pe_1_6_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_3_n3), .Z(
        npu_inst_pe_1_6_3_n22) );
  MUX2_X1 npu_inst_pe_1_6_3_U143 ( .A(npu_inst_pe_1_6_3_n21), .B(
        npu_inst_pe_1_6_3_n18), .S(npu_inst_pe_1_6_3_n7), .Z(
        npu_inst_int_data_x_6__3__1_) );
  MUX2_X1 npu_inst_pe_1_6_3_U142 ( .A(npu_inst_pe_1_6_3_n20), .B(
        npu_inst_pe_1_6_3_n19), .S(npu_inst_pe_1_6_3_n5), .Z(
        npu_inst_pe_1_6_3_n21) );
  MUX2_X1 npu_inst_pe_1_6_3_U141 ( .A(npu_inst_pe_1_6_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_3_n3), .Z(
        npu_inst_pe_1_6_3_n20) );
  MUX2_X1 npu_inst_pe_1_6_3_U140 ( .A(npu_inst_pe_1_6_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_3_n3), .Z(
        npu_inst_pe_1_6_3_n19) );
  MUX2_X1 npu_inst_pe_1_6_3_U139 ( .A(npu_inst_pe_1_6_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_3_n3), .Z(
        npu_inst_pe_1_6_3_n18) );
  MUX2_X1 npu_inst_pe_1_6_3_U138 ( .A(npu_inst_pe_1_6_3_n17), .B(
        npu_inst_pe_1_6_3_n14), .S(npu_inst_pe_1_6_3_n7), .Z(
        npu_inst_int_data_x_6__3__0_) );
  MUX2_X1 npu_inst_pe_1_6_3_U137 ( .A(npu_inst_pe_1_6_3_n16), .B(
        npu_inst_pe_1_6_3_n15), .S(npu_inst_pe_1_6_3_n5), .Z(
        npu_inst_pe_1_6_3_n17) );
  MUX2_X1 npu_inst_pe_1_6_3_U136 ( .A(npu_inst_pe_1_6_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_3_n3), .Z(
        npu_inst_pe_1_6_3_n16) );
  MUX2_X1 npu_inst_pe_1_6_3_U135 ( .A(npu_inst_pe_1_6_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_3_n3), .Z(
        npu_inst_pe_1_6_3_n15) );
  MUX2_X1 npu_inst_pe_1_6_3_U134 ( .A(npu_inst_pe_1_6_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_3_n3), .Z(
        npu_inst_pe_1_6_3_n14) );
  XOR2_X1 npu_inst_pe_1_6_3_U133 ( .A(npu_inst_pe_1_6_3_int_data_0_), .B(
        npu_inst_int_data_res_6__3__0_), .Z(npu_inst_pe_1_6_3_N73) );
  AND2_X1 npu_inst_pe_1_6_3_U132 ( .A1(npu_inst_int_data_res_6__3__0_), .A2(
        npu_inst_pe_1_6_3_int_data_0_), .ZN(npu_inst_pe_1_6_3_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_3_U131 ( .A(npu_inst_int_data_res_6__3__0_), .B(
        npu_inst_pe_1_6_3_n12), .ZN(npu_inst_pe_1_6_3_N65) );
  OR2_X1 npu_inst_pe_1_6_3_U130 ( .A1(npu_inst_pe_1_6_3_n12), .A2(
        npu_inst_int_data_res_6__3__0_), .ZN(npu_inst_pe_1_6_3_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_3_U129 ( .A(npu_inst_int_data_res_6__3__2_), .B(
        npu_inst_pe_1_6_3_add_79_carry_2_), .Z(npu_inst_pe_1_6_3_N75) );
  AND2_X1 npu_inst_pe_1_6_3_U128 ( .A1(npu_inst_pe_1_6_3_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_6__3__2_), .ZN(
        npu_inst_pe_1_6_3_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_3_U127 ( .A(npu_inst_int_data_res_6__3__3_), .B(
        npu_inst_pe_1_6_3_add_79_carry_3_), .Z(npu_inst_pe_1_6_3_N76) );
  AND2_X1 npu_inst_pe_1_6_3_U126 ( .A1(npu_inst_pe_1_6_3_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_6__3__3_), .ZN(
        npu_inst_pe_1_6_3_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_3_U125 ( .A(npu_inst_int_data_res_6__3__4_), .B(
        npu_inst_pe_1_6_3_add_79_carry_4_), .Z(npu_inst_pe_1_6_3_N77) );
  AND2_X1 npu_inst_pe_1_6_3_U124 ( .A1(npu_inst_pe_1_6_3_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_6__3__4_), .ZN(
        npu_inst_pe_1_6_3_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_3_U123 ( .A(npu_inst_int_data_res_6__3__5_), .B(
        npu_inst_pe_1_6_3_add_79_carry_5_), .Z(npu_inst_pe_1_6_3_N78) );
  AND2_X1 npu_inst_pe_1_6_3_U122 ( .A1(npu_inst_pe_1_6_3_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_6__3__5_), .ZN(
        npu_inst_pe_1_6_3_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_3_U121 ( .A(npu_inst_int_data_res_6__3__6_), .B(
        npu_inst_pe_1_6_3_add_79_carry_6_), .Z(npu_inst_pe_1_6_3_N79) );
  AND2_X1 npu_inst_pe_1_6_3_U120 ( .A1(npu_inst_pe_1_6_3_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_6__3__6_), .ZN(
        npu_inst_pe_1_6_3_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_3_U119 ( .A(npu_inst_int_data_res_6__3__7_), .B(
        npu_inst_pe_1_6_3_add_79_carry_7_), .Z(npu_inst_pe_1_6_3_N80) );
  XNOR2_X1 npu_inst_pe_1_6_3_U118 ( .A(npu_inst_pe_1_6_3_sub_77_carry_2_), .B(
        npu_inst_int_data_res_6__3__2_), .ZN(npu_inst_pe_1_6_3_N67) );
  OR2_X1 npu_inst_pe_1_6_3_U117 ( .A1(npu_inst_int_data_res_6__3__2_), .A2(
        npu_inst_pe_1_6_3_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_6_3_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_3_U116 ( .A(npu_inst_pe_1_6_3_sub_77_carry_3_), .B(
        npu_inst_int_data_res_6__3__3_), .ZN(npu_inst_pe_1_6_3_N68) );
  OR2_X1 npu_inst_pe_1_6_3_U115 ( .A1(npu_inst_int_data_res_6__3__3_), .A2(
        npu_inst_pe_1_6_3_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_6_3_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_3_U114 ( .A(npu_inst_pe_1_6_3_sub_77_carry_4_), .B(
        npu_inst_int_data_res_6__3__4_), .ZN(npu_inst_pe_1_6_3_N69) );
  OR2_X1 npu_inst_pe_1_6_3_U113 ( .A1(npu_inst_int_data_res_6__3__4_), .A2(
        npu_inst_pe_1_6_3_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_6_3_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_3_U112 ( .A(npu_inst_pe_1_6_3_sub_77_carry_5_), .B(
        npu_inst_int_data_res_6__3__5_), .ZN(npu_inst_pe_1_6_3_N70) );
  OR2_X1 npu_inst_pe_1_6_3_U111 ( .A1(npu_inst_int_data_res_6__3__5_), .A2(
        npu_inst_pe_1_6_3_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_6_3_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_3_U110 ( .A(npu_inst_pe_1_6_3_sub_77_carry_6_), .B(
        npu_inst_int_data_res_6__3__6_), .ZN(npu_inst_pe_1_6_3_N71) );
  OR2_X1 npu_inst_pe_1_6_3_U109 ( .A1(npu_inst_int_data_res_6__3__6_), .A2(
        npu_inst_pe_1_6_3_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_6_3_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_3_U108 ( .A(npu_inst_int_data_res_6__3__7_), .B(
        npu_inst_pe_1_6_3_sub_77_carry_7_), .ZN(npu_inst_pe_1_6_3_N72) );
  INV_X1 npu_inst_pe_1_6_3_U107 ( .A(npu_inst_n58), .ZN(npu_inst_pe_1_6_3_n6)
         );
  INV_X1 npu_inst_pe_1_6_3_U106 ( .A(npu_inst_pe_1_6_3_n6), .ZN(
        npu_inst_pe_1_6_3_n5) );
  INV_X1 npu_inst_pe_1_6_3_U105 ( .A(npu_inst_n35), .ZN(npu_inst_pe_1_6_3_n2)
         );
  AOI22_X1 npu_inst_pe_1_6_3_U104 ( .A1(npu_inst_int_data_y_7__3__0_), .A2(
        npu_inst_pe_1_6_3_n58), .B1(npu_inst_pe_1_6_3_n118), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_3_n57) );
  INV_X1 npu_inst_pe_1_6_3_U103 ( .A(npu_inst_pe_1_6_3_n57), .ZN(
        npu_inst_pe_1_6_3_n107) );
  AOI22_X1 npu_inst_pe_1_6_3_U102 ( .A1(npu_inst_int_data_y_7__3__0_), .A2(
        npu_inst_pe_1_6_3_n54), .B1(npu_inst_pe_1_6_3_n117), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_3_n53) );
  INV_X1 npu_inst_pe_1_6_3_U99 ( .A(npu_inst_pe_1_6_3_n53), .ZN(
        npu_inst_pe_1_6_3_n108) );
  AOI22_X1 npu_inst_pe_1_6_3_U98 ( .A1(npu_inst_int_data_y_7__3__0_), .A2(
        npu_inst_pe_1_6_3_n50), .B1(npu_inst_pe_1_6_3_n116), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_3_n49) );
  INV_X1 npu_inst_pe_1_6_3_U97 ( .A(npu_inst_pe_1_6_3_n49), .ZN(
        npu_inst_pe_1_6_3_n109) );
  AOI22_X1 npu_inst_pe_1_6_3_U96 ( .A1(npu_inst_int_data_y_7__3__0_), .A2(
        npu_inst_pe_1_6_3_n46), .B1(npu_inst_pe_1_6_3_n115), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_3_n45) );
  INV_X1 npu_inst_pe_1_6_3_U95 ( .A(npu_inst_pe_1_6_3_n45), .ZN(
        npu_inst_pe_1_6_3_n110) );
  AOI22_X1 npu_inst_pe_1_6_3_U94 ( .A1(npu_inst_int_data_y_7__3__0_), .A2(
        npu_inst_pe_1_6_3_n42), .B1(npu_inst_pe_1_6_3_n114), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_3_n41) );
  INV_X1 npu_inst_pe_1_6_3_U93 ( .A(npu_inst_pe_1_6_3_n41), .ZN(
        npu_inst_pe_1_6_3_n111) );
  AOI22_X1 npu_inst_pe_1_6_3_U92 ( .A1(npu_inst_int_data_y_7__3__1_), .A2(
        npu_inst_pe_1_6_3_n58), .B1(npu_inst_pe_1_6_3_n118), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_3_n59) );
  INV_X1 npu_inst_pe_1_6_3_U91 ( .A(npu_inst_pe_1_6_3_n59), .ZN(
        npu_inst_pe_1_6_3_n101) );
  AOI22_X1 npu_inst_pe_1_6_3_U90 ( .A1(npu_inst_int_data_y_7__3__1_), .A2(
        npu_inst_pe_1_6_3_n54), .B1(npu_inst_pe_1_6_3_n117), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_3_n55) );
  INV_X1 npu_inst_pe_1_6_3_U89 ( .A(npu_inst_pe_1_6_3_n55), .ZN(
        npu_inst_pe_1_6_3_n102) );
  AOI22_X1 npu_inst_pe_1_6_3_U88 ( .A1(npu_inst_int_data_y_7__3__1_), .A2(
        npu_inst_pe_1_6_3_n50), .B1(npu_inst_pe_1_6_3_n116), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_3_n51) );
  INV_X1 npu_inst_pe_1_6_3_U87 ( .A(npu_inst_pe_1_6_3_n51), .ZN(
        npu_inst_pe_1_6_3_n103) );
  AOI22_X1 npu_inst_pe_1_6_3_U86 ( .A1(npu_inst_int_data_y_7__3__1_), .A2(
        npu_inst_pe_1_6_3_n46), .B1(npu_inst_pe_1_6_3_n115), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_3_n47) );
  INV_X1 npu_inst_pe_1_6_3_U85 ( .A(npu_inst_pe_1_6_3_n47), .ZN(
        npu_inst_pe_1_6_3_n104) );
  AOI22_X1 npu_inst_pe_1_6_3_U84 ( .A1(npu_inst_int_data_y_7__3__1_), .A2(
        npu_inst_pe_1_6_3_n42), .B1(npu_inst_pe_1_6_3_n114), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_3_n43) );
  INV_X1 npu_inst_pe_1_6_3_U83 ( .A(npu_inst_pe_1_6_3_n43), .ZN(
        npu_inst_pe_1_6_3_n105) );
  AOI22_X1 npu_inst_pe_1_6_3_U82 ( .A1(npu_inst_pe_1_6_3_n38), .A2(
        npu_inst_int_data_y_7__3__1_), .B1(npu_inst_pe_1_6_3_n113), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_3_n39) );
  INV_X1 npu_inst_pe_1_6_3_U81 ( .A(npu_inst_pe_1_6_3_n39), .ZN(
        npu_inst_pe_1_6_3_n106) );
  AND2_X1 npu_inst_pe_1_6_3_U80 ( .A1(npu_inst_pe_1_6_3_N93), .A2(npu_inst_n35), .ZN(npu_inst_int_data_y_6__3__0_) );
  NAND2_X1 npu_inst_pe_1_6_3_U79 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_3_n60), .ZN(npu_inst_pe_1_6_3_n74) );
  OAI21_X1 npu_inst_pe_1_6_3_U78 ( .B1(npu_inst_pe_1_6_3_n63), .B2(
        npu_inst_pe_1_6_3_n60), .A(npu_inst_pe_1_6_3_n74), .ZN(
        npu_inst_pe_1_6_3_n97) );
  NAND2_X1 npu_inst_pe_1_6_3_U77 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_3_n60), .ZN(npu_inst_pe_1_6_3_n73) );
  OAI21_X1 npu_inst_pe_1_6_3_U76 ( .B1(npu_inst_pe_1_6_3_n61), .B2(
        npu_inst_pe_1_6_3_n60), .A(npu_inst_pe_1_6_3_n73), .ZN(
        npu_inst_pe_1_6_3_n96) );
  NAND2_X1 npu_inst_pe_1_6_3_U75 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_3_n56), .ZN(npu_inst_pe_1_6_3_n72) );
  OAI21_X1 npu_inst_pe_1_6_3_U74 ( .B1(npu_inst_pe_1_6_3_n63), .B2(
        npu_inst_pe_1_6_3_n56), .A(npu_inst_pe_1_6_3_n72), .ZN(
        npu_inst_pe_1_6_3_n95) );
  NAND2_X1 npu_inst_pe_1_6_3_U73 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_3_n56), .ZN(npu_inst_pe_1_6_3_n71) );
  OAI21_X1 npu_inst_pe_1_6_3_U72 ( .B1(npu_inst_pe_1_6_3_n61), .B2(
        npu_inst_pe_1_6_3_n56), .A(npu_inst_pe_1_6_3_n71), .ZN(
        npu_inst_pe_1_6_3_n94) );
  NAND2_X1 npu_inst_pe_1_6_3_U71 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_3_n52), .ZN(npu_inst_pe_1_6_3_n70) );
  OAI21_X1 npu_inst_pe_1_6_3_U70 ( .B1(npu_inst_pe_1_6_3_n63), .B2(
        npu_inst_pe_1_6_3_n52), .A(npu_inst_pe_1_6_3_n70), .ZN(
        npu_inst_pe_1_6_3_n93) );
  NAND2_X1 npu_inst_pe_1_6_3_U69 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_3_n52), .ZN(npu_inst_pe_1_6_3_n69) );
  OAI21_X1 npu_inst_pe_1_6_3_U68 ( .B1(npu_inst_pe_1_6_3_n61), .B2(
        npu_inst_pe_1_6_3_n52), .A(npu_inst_pe_1_6_3_n69), .ZN(
        npu_inst_pe_1_6_3_n92) );
  NAND2_X1 npu_inst_pe_1_6_3_U67 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_3_n48), .ZN(npu_inst_pe_1_6_3_n68) );
  OAI21_X1 npu_inst_pe_1_6_3_U66 ( .B1(npu_inst_pe_1_6_3_n63), .B2(
        npu_inst_pe_1_6_3_n48), .A(npu_inst_pe_1_6_3_n68), .ZN(
        npu_inst_pe_1_6_3_n91) );
  NAND2_X1 npu_inst_pe_1_6_3_U65 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_3_n48), .ZN(npu_inst_pe_1_6_3_n67) );
  OAI21_X1 npu_inst_pe_1_6_3_U64 ( .B1(npu_inst_pe_1_6_3_n61), .B2(
        npu_inst_pe_1_6_3_n48), .A(npu_inst_pe_1_6_3_n67), .ZN(
        npu_inst_pe_1_6_3_n90) );
  NAND2_X1 npu_inst_pe_1_6_3_U63 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_3_n44), .ZN(npu_inst_pe_1_6_3_n66) );
  OAI21_X1 npu_inst_pe_1_6_3_U62 ( .B1(npu_inst_pe_1_6_3_n63), .B2(
        npu_inst_pe_1_6_3_n44), .A(npu_inst_pe_1_6_3_n66), .ZN(
        npu_inst_pe_1_6_3_n89) );
  NAND2_X1 npu_inst_pe_1_6_3_U61 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_3_n44), .ZN(npu_inst_pe_1_6_3_n65) );
  OAI21_X1 npu_inst_pe_1_6_3_U60 ( .B1(npu_inst_pe_1_6_3_n61), .B2(
        npu_inst_pe_1_6_3_n44), .A(npu_inst_pe_1_6_3_n65), .ZN(
        npu_inst_pe_1_6_3_n88) );
  NAND2_X1 npu_inst_pe_1_6_3_U59 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_3_n40), .ZN(npu_inst_pe_1_6_3_n64) );
  OAI21_X1 npu_inst_pe_1_6_3_U58 ( .B1(npu_inst_pe_1_6_3_n63), .B2(
        npu_inst_pe_1_6_3_n40), .A(npu_inst_pe_1_6_3_n64), .ZN(
        npu_inst_pe_1_6_3_n87) );
  NAND2_X1 npu_inst_pe_1_6_3_U57 ( .A1(npu_inst_pe_1_6_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_3_n40), .ZN(npu_inst_pe_1_6_3_n62) );
  OAI21_X1 npu_inst_pe_1_6_3_U56 ( .B1(npu_inst_pe_1_6_3_n61), .B2(
        npu_inst_pe_1_6_3_n40), .A(npu_inst_pe_1_6_3_n62), .ZN(
        npu_inst_pe_1_6_3_n86) );
  AOI22_X1 npu_inst_pe_1_6_3_U55 ( .A1(npu_inst_pe_1_6_3_n38), .A2(
        npu_inst_int_data_y_7__3__0_), .B1(npu_inst_pe_1_6_3_n113), .B2(
        npu_inst_pe_1_6_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_3_n37) );
  INV_X1 npu_inst_pe_1_6_3_U54 ( .A(npu_inst_pe_1_6_3_n37), .ZN(
        npu_inst_pe_1_6_3_n112) );
  AND2_X1 npu_inst_pe_1_6_3_U53 ( .A1(npu_inst_n35), .A2(npu_inst_pe_1_6_3_N94), .ZN(npu_inst_int_data_y_6__3__1_) );
  AOI222_X1 npu_inst_pe_1_6_3_U52 ( .A1(npu_inst_int_data_res_7__3__0_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N73), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N65), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n84) );
  INV_X1 npu_inst_pe_1_6_3_U51 ( .A(npu_inst_pe_1_6_3_n84), .ZN(
        npu_inst_pe_1_6_3_n100) );
  AOI222_X1 npu_inst_pe_1_6_3_U50 ( .A1(npu_inst_pe_1_6_3_n1), .A2(
        npu_inst_int_data_res_7__3__7_), .B1(npu_inst_pe_1_6_3_N80), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N72), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n75) );
  INV_X1 npu_inst_pe_1_6_3_U49 ( .A(npu_inst_pe_1_6_3_n75), .ZN(
        npu_inst_pe_1_6_3_n32) );
  AOI222_X1 npu_inst_pe_1_6_3_U48 ( .A1(npu_inst_int_data_res_7__3__1_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N74), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N66), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n83) );
  INV_X1 npu_inst_pe_1_6_3_U47 ( .A(npu_inst_pe_1_6_3_n83), .ZN(
        npu_inst_pe_1_6_3_n99) );
  AOI222_X1 npu_inst_pe_1_6_3_U46 ( .A1(npu_inst_int_data_res_7__3__3_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N76), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N68), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n81) );
  INV_X1 npu_inst_pe_1_6_3_U45 ( .A(npu_inst_pe_1_6_3_n81), .ZN(
        npu_inst_pe_1_6_3_n36) );
  AOI222_X1 npu_inst_pe_1_6_3_U44 ( .A1(npu_inst_int_data_res_7__3__4_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N77), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N69), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n80) );
  INV_X1 npu_inst_pe_1_6_3_U43 ( .A(npu_inst_pe_1_6_3_n80), .ZN(
        npu_inst_pe_1_6_3_n35) );
  AOI222_X1 npu_inst_pe_1_6_3_U42 ( .A1(npu_inst_int_data_res_7__3__5_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N78), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N70), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n79) );
  INV_X1 npu_inst_pe_1_6_3_U41 ( .A(npu_inst_pe_1_6_3_n79), .ZN(
        npu_inst_pe_1_6_3_n34) );
  AOI222_X1 npu_inst_pe_1_6_3_U40 ( .A1(npu_inst_int_data_res_7__3__6_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N79), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N71), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n78) );
  INV_X1 npu_inst_pe_1_6_3_U39 ( .A(npu_inst_pe_1_6_3_n78), .ZN(
        npu_inst_pe_1_6_3_n33) );
  AND2_X1 npu_inst_pe_1_6_3_U38 ( .A1(npu_inst_int_data_x_6__3__1_), .A2(
        npu_inst_pe_1_6_3_int_q_weight_1_), .ZN(npu_inst_pe_1_6_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_3_U37 ( .A1(npu_inst_int_data_x_6__3__0_), .A2(
        npu_inst_pe_1_6_3_int_q_weight_1_), .ZN(npu_inst_pe_1_6_3_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_6_3_U36 ( .A(npu_inst_pe_1_6_3_int_data_1_), .ZN(
        npu_inst_pe_1_6_3_n13) );
  NOR3_X1 npu_inst_pe_1_6_3_U35 ( .A1(npu_inst_pe_1_6_3_n26), .A2(npu_inst_n35), .A3(npu_inst_int_ckg[12]), .ZN(npu_inst_pe_1_6_3_n85) );
  OR2_X1 npu_inst_pe_1_6_3_U34 ( .A1(npu_inst_pe_1_6_3_n85), .A2(
        npu_inst_pe_1_6_3_n1), .ZN(npu_inst_pe_1_6_3_N84) );
  AOI222_X1 npu_inst_pe_1_6_3_U33 ( .A1(npu_inst_int_data_res_7__3__2_), .A2(
        npu_inst_pe_1_6_3_n1), .B1(npu_inst_pe_1_6_3_N75), .B2(
        npu_inst_pe_1_6_3_n76), .C1(npu_inst_pe_1_6_3_N67), .C2(
        npu_inst_pe_1_6_3_n77), .ZN(npu_inst_pe_1_6_3_n82) );
  INV_X1 npu_inst_pe_1_6_3_U32 ( .A(npu_inst_pe_1_6_3_n82), .ZN(
        npu_inst_pe_1_6_3_n98) );
  AOI22_X1 npu_inst_pe_1_6_3_U31 ( .A1(npu_inst_n35), .A2(
        npu_inst_int_data_y_7__3__1_), .B1(npu_inst_pe_1_6_3_n2), .B2(
        npu_inst_int_data_x_6__4__1_), .ZN(npu_inst_pe_1_6_3_n63) );
  AOI22_X1 npu_inst_pe_1_6_3_U30 ( .A1(npu_inst_n35), .A2(
        npu_inst_int_data_y_7__3__0_), .B1(npu_inst_pe_1_6_3_n2), .B2(
        npu_inst_int_data_x_6__4__0_), .ZN(npu_inst_pe_1_6_3_n61) );
  INV_X1 npu_inst_pe_1_6_3_U29 ( .A(npu_inst_pe_1_6_3_int_data_0_), .ZN(
        npu_inst_pe_1_6_3_n12) );
  INV_X1 npu_inst_pe_1_6_3_U28 ( .A(npu_inst_n50), .ZN(npu_inst_pe_1_6_3_n4)
         );
  OR3_X1 npu_inst_pe_1_6_3_U27 ( .A1(npu_inst_pe_1_6_3_n5), .A2(
        npu_inst_pe_1_6_3_n7), .A3(npu_inst_pe_1_6_3_n4), .ZN(
        npu_inst_pe_1_6_3_n56) );
  OR3_X1 npu_inst_pe_1_6_3_U26 ( .A1(npu_inst_pe_1_6_3_n4), .A2(
        npu_inst_pe_1_6_3_n7), .A3(npu_inst_pe_1_6_3_n6), .ZN(
        npu_inst_pe_1_6_3_n48) );
  INV_X1 npu_inst_pe_1_6_3_U25 ( .A(npu_inst_pe_1_6_3_n4), .ZN(
        npu_inst_pe_1_6_3_n3) );
  OR3_X1 npu_inst_pe_1_6_3_U24 ( .A1(npu_inst_pe_1_6_3_n3), .A2(
        npu_inst_pe_1_6_3_n7), .A3(npu_inst_pe_1_6_3_n6), .ZN(
        npu_inst_pe_1_6_3_n52) );
  OR3_X1 npu_inst_pe_1_6_3_U23 ( .A1(npu_inst_pe_1_6_3_n5), .A2(
        npu_inst_pe_1_6_3_n7), .A3(npu_inst_pe_1_6_3_n3), .ZN(
        npu_inst_pe_1_6_3_n60) );
  BUF_X1 npu_inst_pe_1_6_3_U22 ( .A(npu_inst_n15), .Z(npu_inst_pe_1_6_3_n1) );
  NOR2_X1 npu_inst_pe_1_6_3_U21 ( .A1(npu_inst_pe_1_6_3_n60), .A2(
        npu_inst_pe_1_6_3_n2), .ZN(npu_inst_pe_1_6_3_n58) );
  NOR2_X1 npu_inst_pe_1_6_3_U20 ( .A1(npu_inst_pe_1_6_3_n56), .A2(
        npu_inst_pe_1_6_3_n2), .ZN(npu_inst_pe_1_6_3_n54) );
  NOR2_X1 npu_inst_pe_1_6_3_U19 ( .A1(npu_inst_pe_1_6_3_n52), .A2(
        npu_inst_pe_1_6_3_n2), .ZN(npu_inst_pe_1_6_3_n50) );
  NOR2_X1 npu_inst_pe_1_6_3_U18 ( .A1(npu_inst_pe_1_6_3_n48), .A2(
        npu_inst_pe_1_6_3_n2), .ZN(npu_inst_pe_1_6_3_n46) );
  NOR2_X1 npu_inst_pe_1_6_3_U17 ( .A1(npu_inst_pe_1_6_3_n40), .A2(
        npu_inst_pe_1_6_3_n2), .ZN(npu_inst_pe_1_6_3_n38) );
  NOR2_X1 npu_inst_pe_1_6_3_U16 ( .A1(npu_inst_pe_1_6_3_n44), .A2(
        npu_inst_pe_1_6_3_n2), .ZN(npu_inst_pe_1_6_3_n42) );
  BUF_X1 npu_inst_pe_1_6_3_U15 ( .A(npu_inst_n77), .Z(npu_inst_pe_1_6_3_n7) );
  INV_X1 npu_inst_pe_1_6_3_U14 ( .A(npu_inst_n105), .ZN(npu_inst_pe_1_6_3_n11)
         );
  INV_X1 npu_inst_pe_1_6_3_U13 ( .A(npu_inst_pe_1_6_3_n38), .ZN(
        npu_inst_pe_1_6_3_n113) );
  INV_X1 npu_inst_pe_1_6_3_U12 ( .A(npu_inst_pe_1_6_3_n58), .ZN(
        npu_inst_pe_1_6_3_n118) );
  INV_X1 npu_inst_pe_1_6_3_U11 ( .A(npu_inst_pe_1_6_3_n54), .ZN(
        npu_inst_pe_1_6_3_n117) );
  INV_X1 npu_inst_pe_1_6_3_U10 ( .A(npu_inst_pe_1_6_3_n50), .ZN(
        npu_inst_pe_1_6_3_n116) );
  INV_X1 npu_inst_pe_1_6_3_U9 ( .A(npu_inst_pe_1_6_3_n46), .ZN(
        npu_inst_pe_1_6_3_n115) );
  INV_X1 npu_inst_pe_1_6_3_U8 ( .A(npu_inst_pe_1_6_3_n42), .ZN(
        npu_inst_pe_1_6_3_n114) );
  BUF_X1 npu_inst_pe_1_6_3_U7 ( .A(npu_inst_pe_1_6_3_n11), .Z(
        npu_inst_pe_1_6_3_n10) );
  BUF_X1 npu_inst_pe_1_6_3_U6 ( .A(npu_inst_pe_1_6_3_n11), .Z(
        npu_inst_pe_1_6_3_n9) );
  BUF_X1 npu_inst_pe_1_6_3_U5 ( .A(npu_inst_pe_1_6_3_n11), .Z(
        npu_inst_pe_1_6_3_n8) );
  NOR2_X1 npu_inst_pe_1_6_3_U4 ( .A1(npu_inst_pe_1_6_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_3_n1), .ZN(npu_inst_pe_1_6_3_n76) );
  NOR2_X1 npu_inst_pe_1_6_3_U3 ( .A1(npu_inst_pe_1_6_3_n27), .A2(
        npu_inst_pe_1_6_3_n1), .ZN(npu_inst_pe_1_6_3_n77) );
  FA_X1 npu_inst_pe_1_6_3_sub_77_U2_1 ( .A(npu_inst_int_data_res_6__3__1_), 
        .B(npu_inst_pe_1_6_3_n13), .CI(npu_inst_pe_1_6_3_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_6_3_sub_77_carry_2_), .S(npu_inst_pe_1_6_3_N66) );
  FA_X1 npu_inst_pe_1_6_3_add_79_U1_1 ( .A(npu_inst_int_data_res_6__3__1_), 
        .B(npu_inst_pe_1_6_3_int_data_1_), .CI(
        npu_inst_pe_1_6_3_add_79_carry_1_), .CO(
        npu_inst_pe_1_6_3_add_79_carry_2_), .S(npu_inst_pe_1_6_3_N74) );
  NAND3_X1 npu_inst_pe_1_6_3_U101 ( .A1(npu_inst_pe_1_6_3_n4), .A2(
        npu_inst_pe_1_6_3_n6), .A3(npu_inst_pe_1_6_3_n7), .ZN(
        npu_inst_pe_1_6_3_n44) );
  NAND3_X1 npu_inst_pe_1_6_3_U100 ( .A1(npu_inst_pe_1_6_3_n3), .A2(
        npu_inst_pe_1_6_3_n6), .A3(npu_inst_pe_1_6_3_n7), .ZN(
        npu_inst_pe_1_6_3_n40) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_3_n33), .CK(
        npu_inst_pe_1_6_3_net3305), .RN(npu_inst_pe_1_6_3_n8), .Q(
        npu_inst_int_data_res_6__3__6_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_3_n34), .CK(
        npu_inst_pe_1_6_3_net3305), .RN(npu_inst_pe_1_6_3_n8), .Q(
        npu_inst_int_data_res_6__3__5_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_3_n35), .CK(
        npu_inst_pe_1_6_3_net3305), .RN(npu_inst_pe_1_6_3_n8), .Q(
        npu_inst_int_data_res_6__3__4_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_3_n36), .CK(
        npu_inst_pe_1_6_3_net3305), .RN(npu_inst_pe_1_6_3_n8), .Q(
        npu_inst_int_data_res_6__3__3_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_3_n98), .CK(
        npu_inst_pe_1_6_3_net3305), .RN(npu_inst_pe_1_6_3_n8), .Q(
        npu_inst_int_data_res_6__3__2_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_3_n99), .CK(
        npu_inst_pe_1_6_3_net3305), .RN(npu_inst_pe_1_6_3_n8), .Q(
        npu_inst_int_data_res_6__3__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_3_n32), .CK(
        npu_inst_pe_1_6_3_net3305), .RN(npu_inst_pe_1_6_3_n8), .Q(
        npu_inst_int_data_res_6__3__7_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_3_n100), 
        .CK(npu_inst_pe_1_6_3_net3305), .RN(npu_inst_pe_1_6_3_n8), .Q(
        npu_inst_int_data_res_6__3__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_weight_reg_0_ ( .D(npu_inst_n91), .CK(
        npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n8), .Q(
        npu_inst_pe_1_6_3_int_q_weight_0_), .QN(npu_inst_pe_1_6_3_n27) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_weight_reg_1_ ( .D(npu_inst_n97), .CK(
        npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n8), .Q(
        npu_inst_pe_1_6_3_int_q_weight_1_), .QN(npu_inst_pe_1_6_3_n26) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_3_n112), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n8), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_3_n106), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n8), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_3_n111), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_3_n105), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_3_n110), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_3_n104), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_3_n109), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_3_n103), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_3_n108), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_3_n102), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_3_n107), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_3_n101), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_3_n86), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_3_n87), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n9), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_3_n88), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_3_n89), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_3_n90), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_3_n91), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_3_n92), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_3_n93), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_3_n94), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_3_n95), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_3_n96), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_3_n97), 
        .CK(npu_inst_pe_1_6_3_net3311), .RN(npu_inst_pe_1_6_3_n10), .Q(
        npu_inst_pe_1_6_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_3_net3305) );
  CLKGATETST_X1 npu_inst_pe_1_6_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n44), .SE(1'b0), .GCK(npu_inst_pe_1_6_3_net3311) );
  MUX2_X1 npu_inst_pe_1_6_4_U152 ( .A(npu_inst_pe_1_6_4_n30), .B(
        npu_inst_pe_1_6_4_n25), .S(npu_inst_pe_1_6_4_n6), .Z(
        npu_inst_pe_1_6_4_N93) );
  MUX2_X1 npu_inst_pe_1_6_4_U151 ( .A(npu_inst_pe_1_6_4_n29), .B(
        npu_inst_pe_1_6_4_n28), .S(npu_inst_n57), .Z(npu_inst_pe_1_6_4_n30) );
  MUX2_X1 npu_inst_pe_1_6_4_U150 ( .A(npu_inst_pe_1_6_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_4_n3), .Z(
        npu_inst_pe_1_6_4_n29) );
  MUX2_X1 npu_inst_pe_1_6_4_U149 ( .A(npu_inst_pe_1_6_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_4_n3), .Z(
        npu_inst_pe_1_6_4_n28) );
  MUX2_X1 npu_inst_pe_1_6_4_U148 ( .A(npu_inst_pe_1_6_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_4_n3), .Z(
        npu_inst_pe_1_6_4_n25) );
  MUX2_X1 npu_inst_pe_1_6_4_U147 ( .A(npu_inst_pe_1_6_4_n24), .B(
        npu_inst_pe_1_6_4_n21), .S(npu_inst_pe_1_6_4_n6), .Z(
        npu_inst_pe_1_6_4_N94) );
  MUX2_X1 npu_inst_pe_1_6_4_U146 ( .A(npu_inst_pe_1_6_4_n23), .B(
        npu_inst_pe_1_6_4_n22), .S(npu_inst_n57), .Z(npu_inst_pe_1_6_4_n24) );
  MUX2_X1 npu_inst_pe_1_6_4_U145 ( .A(npu_inst_pe_1_6_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_4_n3), .Z(
        npu_inst_pe_1_6_4_n23) );
  MUX2_X1 npu_inst_pe_1_6_4_U144 ( .A(npu_inst_pe_1_6_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_4_n3), .Z(
        npu_inst_pe_1_6_4_n22) );
  MUX2_X1 npu_inst_pe_1_6_4_U143 ( .A(npu_inst_pe_1_6_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_4_n3), .Z(
        npu_inst_pe_1_6_4_n21) );
  MUX2_X1 npu_inst_pe_1_6_4_U142 ( .A(npu_inst_pe_1_6_4_n20), .B(
        npu_inst_pe_1_6_4_n17), .S(npu_inst_pe_1_6_4_n6), .Z(
        npu_inst_int_data_x_6__4__1_) );
  MUX2_X1 npu_inst_pe_1_6_4_U141 ( .A(npu_inst_pe_1_6_4_n19), .B(
        npu_inst_pe_1_6_4_n18), .S(npu_inst_n57), .Z(npu_inst_pe_1_6_4_n20) );
  MUX2_X1 npu_inst_pe_1_6_4_U140 ( .A(npu_inst_pe_1_6_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_4_n3), .Z(
        npu_inst_pe_1_6_4_n19) );
  MUX2_X1 npu_inst_pe_1_6_4_U139 ( .A(npu_inst_pe_1_6_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_4_n3), .Z(
        npu_inst_pe_1_6_4_n18) );
  MUX2_X1 npu_inst_pe_1_6_4_U138 ( .A(npu_inst_pe_1_6_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_4_n3), .Z(
        npu_inst_pe_1_6_4_n17) );
  MUX2_X1 npu_inst_pe_1_6_4_U137 ( .A(npu_inst_pe_1_6_4_n16), .B(
        npu_inst_pe_1_6_4_n13), .S(npu_inst_pe_1_6_4_n6), .Z(
        npu_inst_int_data_x_6__4__0_) );
  MUX2_X1 npu_inst_pe_1_6_4_U136 ( .A(npu_inst_pe_1_6_4_n15), .B(
        npu_inst_pe_1_6_4_n14), .S(npu_inst_n57), .Z(npu_inst_pe_1_6_4_n16) );
  MUX2_X1 npu_inst_pe_1_6_4_U135 ( .A(npu_inst_pe_1_6_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_4_n3), .Z(
        npu_inst_pe_1_6_4_n15) );
  MUX2_X1 npu_inst_pe_1_6_4_U134 ( .A(npu_inst_pe_1_6_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_4_n3), .Z(
        npu_inst_pe_1_6_4_n14) );
  MUX2_X1 npu_inst_pe_1_6_4_U133 ( .A(npu_inst_pe_1_6_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_4_n3), .Z(
        npu_inst_pe_1_6_4_n13) );
  XOR2_X1 npu_inst_pe_1_6_4_U132 ( .A(npu_inst_pe_1_6_4_int_data_0_), .B(
        npu_inst_int_data_res_6__4__0_), .Z(npu_inst_pe_1_6_4_N73) );
  AND2_X1 npu_inst_pe_1_6_4_U131 ( .A1(npu_inst_int_data_res_6__4__0_), .A2(
        npu_inst_pe_1_6_4_int_data_0_), .ZN(npu_inst_pe_1_6_4_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_4_U130 ( .A(npu_inst_int_data_res_6__4__0_), .B(
        npu_inst_pe_1_6_4_n11), .ZN(npu_inst_pe_1_6_4_N65) );
  OR2_X1 npu_inst_pe_1_6_4_U129 ( .A1(npu_inst_pe_1_6_4_n11), .A2(
        npu_inst_int_data_res_6__4__0_), .ZN(npu_inst_pe_1_6_4_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_4_U128 ( .A(npu_inst_int_data_res_6__4__2_), .B(
        npu_inst_pe_1_6_4_add_79_carry_2_), .Z(npu_inst_pe_1_6_4_N75) );
  AND2_X1 npu_inst_pe_1_6_4_U127 ( .A1(npu_inst_pe_1_6_4_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_6__4__2_), .ZN(
        npu_inst_pe_1_6_4_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_4_U126 ( .A(npu_inst_int_data_res_6__4__3_), .B(
        npu_inst_pe_1_6_4_add_79_carry_3_), .Z(npu_inst_pe_1_6_4_N76) );
  AND2_X1 npu_inst_pe_1_6_4_U125 ( .A1(npu_inst_pe_1_6_4_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_6__4__3_), .ZN(
        npu_inst_pe_1_6_4_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_4_U124 ( .A(npu_inst_int_data_res_6__4__4_), .B(
        npu_inst_pe_1_6_4_add_79_carry_4_), .Z(npu_inst_pe_1_6_4_N77) );
  AND2_X1 npu_inst_pe_1_6_4_U123 ( .A1(npu_inst_pe_1_6_4_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_6__4__4_), .ZN(
        npu_inst_pe_1_6_4_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_4_U122 ( .A(npu_inst_int_data_res_6__4__5_), .B(
        npu_inst_pe_1_6_4_add_79_carry_5_), .Z(npu_inst_pe_1_6_4_N78) );
  AND2_X1 npu_inst_pe_1_6_4_U121 ( .A1(npu_inst_pe_1_6_4_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_6__4__5_), .ZN(
        npu_inst_pe_1_6_4_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_4_U120 ( .A(npu_inst_int_data_res_6__4__6_), .B(
        npu_inst_pe_1_6_4_add_79_carry_6_), .Z(npu_inst_pe_1_6_4_N79) );
  AND2_X1 npu_inst_pe_1_6_4_U119 ( .A1(npu_inst_pe_1_6_4_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_6__4__6_), .ZN(
        npu_inst_pe_1_6_4_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_4_U118 ( .A(npu_inst_int_data_res_6__4__7_), .B(
        npu_inst_pe_1_6_4_add_79_carry_7_), .Z(npu_inst_pe_1_6_4_N80) );
  XNOR2_X1 npu_inst_pe_1_6_4_U117 ( .A(npu_inst_pe_1_6_4_sub_77_carry_2_), .B(
        npu_inst_int_data_res_6__4__2_), .ZN(npu_inst_pe_1_6_4_N67) );
  OR2_X1 npu_inst_pe_1_6_4_U116 ( .A1(npu_inst_int_data_res_6__4__2_), .A2(
        npu_inst_pe_1_6_4_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_6_4_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_4_U115 ( .A(npu_inst_pe_1_6_4_sub_77_carry_3_), .B(
        npu_inst_int_data_res_6__4__3_), .ZN(npu_inst_pe_1_6_4_N68) );
  OR2_X1 npu_inst_pe_1_6_4_U114 ( .A1(npu_inst_int_data_res_6__4__3_), .A2(
        npu_inst_pe_1_6_4_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_6_4_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_4_U113 ( .A(npu_inst_pe_1_6_4_sub_77_carry_4_), .B(
        npu_inst_int_data_res_6__4__4_), .ZN(npu_inst_pe_1_6_4_N69) );
  OR2_X1 npu_inst_pe_1_6_4_U112 ( .A1(npu_inst_int_data_res_6__4__4_), .A2(
        npu_inst_pe_1_6_4_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_6_4_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_4_U111 ( .A(npu_inst_pe_1_6_4_sub_77_carry_5_), .B(
        npu_inst_int_data_res_6__4__5_), .ZN(npu_inst_pe_1_6_4_N70) );
  OR2_X1 npu_inst_pe_1_6_4_U110 ( .A1(npu_inst_int_data_res_6__4__5_), .A2(
        npu_inst_pe_1_6_4_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_6_4_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_4_U109 ( .A(npu_inst_pe_1_6_4_sub_77_carry_6_), .B(
        npu_inst_int_data_res_6__4__6_), .ZN(npu_inst_pe_1_6_4_N71) );
  OR2_X1 npu_inst_pe_1_6_4_U108 ( .A1(npu_inst_int_data_res_6__4__6_), .A2(
        npu_inst_pe_1_6_4_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_6_4_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_4_U107 ( .A(npu_inst_int_data_res_6__4__7_), .B(
        npu_inst_pe_1_6_4_sub_77_carry_7_), .ZN(npu_inst_pe_1_6_4_N72) );
  INV_X1 npu_inst_pe_1_6_4_U106 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_6_4_n5)
         );
  INV_X1 npu_inst_pe_1_6_4_U105 ( .A(npu_inst_n35), .ZN(npu_inst_pe_1_6_4_n2)
         );
  AOI22_X1 npu_inst_pe_1_6_4_U104 ( .A1(npu_inst_int_data_y_7__4__0_), .A2(
        npu_inst_pe_1_6_4_n58), .B1(npu_inst_pe_1_6_4_n117), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_4_n57) );
  INV_X1 npu_inst_pe_1_6_4_U103 ( .A(npu_inst_pe_1_6_4_n57), .ZN(
        npu_inst_pe_1_6_4_n106) );
  AOI22_X1 npu_inst_pe_1_6_4_U102 ( .A1(npu_inst_int_data_y_7__4__0_), .A2(
        npu_inst_pe_1_6_4_n54), .B1(npu_inst_pe_1_6_4_n116), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_4_n53) );
  INV_X1 npu_inst_pe_1_6_4_U99 ( .A(npu_inst_pe_1_6_4_n53), .ZN(
        npu_inst_pe_1_6_4_n107) );
  AOI22_X1 npu_inst_pe_1_6_4_U98 ( .A1(npu_inst_int_data_y_7__4__0_), .A2(
        npu_inst_pe_1_6_4_n50), .B1(npu_inst_pe_1_6_4_n115), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_4_n49) );
  INV_X1 npu_inst_pe_1_6_4_U97 ( .A(npu_inst_pe_1_6_4_n49), .ZN(
        npu_inst_pe_1_6_4_n108) );
  AOI22_X1 npu_inst_pe_1_6_4_U96 ( .A1(npu_inst_int_data_y_7__4__0_), .A2(
        npu_inst_pe_1_6_4_n46), .B1(npu_inst_pe_1_6_4_n114), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_4_n45) );
  INV_X1 npu_inst_pe_1_6_4_U95 ( .A(npu_inst_pe_1_6_4_n45), .ZN(
        npu_inst_pe_1_6_4_n109) );
  AOI22_X1 npu_inst_pe_1_6_4_U94 ( .A1(npu_inst_int_data_y_7__4__0_), .A2(
        npu_inst_pe_1_6_4_n42), .B1(npu_inst_pe_1_6_4_n113), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_4_n41) );
  INV_X1 npu_inst_pe_1_6_4_U93 ( .A(npu_inst_pe_1_6_4_n41), .ZN(
        npu_inst_pe_1_6_4_n110) );
  AOI22_X1 npu_inst_pe_1_6_4_U92 ( .A1(npu_inst_int_data_y_7__4__1_), .A2(
        npu_inst_pe_1_6_4_n58), .B1(npu_inst_pe_1_6_4_n117), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_4_n59) );
  INV_X1 npu_inst_pe_1_6_4_U91 ( .A(npu_inst_pe_1_6_4_n59), .ZN(
        npu_inst_pe_1_6_4_n100) );
  AOI22_X1 npu_inst_pe_1_6_4_U90 ( .A1(npu_inst_int_data_y_7__4__1_), .A2(
        npu_inst_pe_1_6_4_n54), .B1(npu_inst_pe_1_6_4_n116), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_4_n55) );
  INV_X1 npu_inst_pe_1_6_4_U89 ( .A(npu_inst_pe_1_6_4_n55), .ZN(
        npu_inst_pe_1_6_4_n101) );
  AOI22_X1 npu_inst_pe_1_6_4_U88 ( .A1(npu_inst_int_data_y_7__4__1_), .A2(
        npu_inst_pe_1_6_4_n50), .B1(npu_inst_pe_1_6_4_n115), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_4_n51) );
  INV_X1 npu_inst_pe_1_6_4_U87 ( .A(npu_inst_pe_1_6_4_n51), .ZN(
        npu_inst_pe_1_6_4_n102) );
  AOI22_X1 npu_inst_pe_1_6_4_U86 ( .A1(npu_inst_int_data_y_7__4__1_), .A2(
        npu_inst_pe_1_6_4_n46), .B1(npu_inst_pe_1_6_4_n114), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_4_n47) );
  INV_X1 npu_inst_pe_1_6_4_U85 ( .A(npu_inst_pe_1_6_4_n47), .ZN(
        npu_inst_pe_1_6_4_n103) );
  AOI22_X1 npu_inst_pe_1_6_4_U84 ( .A1(npu_inst_int_data_y_7__4__1_), .A2(
        npu_inst_pe_1_6_4_n42), .B1(npu_inst_pe_1_6_4_n113), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_4_n43) );
  INV_X1 npu_inst_pe_1_6_4_U83 ( .A(npu_inst_pe_1_6_4_n43), .ZN(
        npu_inst_pe_1_6_4_n104) );
  AOI22_X1 npu_inst_pe_1_6_4_U82 ( .A1(npu_inst_pe_1_6_4_n38), .A2(
        npu_inst_int_data_y_7__4__1_), .B1(npu_inst_pe_1_6_4_n112), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_4_n39) );
  INV_X1 npu_inst_pe_1_6_4_U81 ( .A(npu_inst_pe_1_6_4_n39), .ZN(
        npu_inst_pe_1_6_4_n105) );
  AND2_X1 npu_inst_pe_1_6_4_U80 ( .A1(npu_inst_pe_1_6_4_N93), .A2(npu_inst_n35), .ZN(npu_inst_int_data_y_6__4__0_) );
  NAND2_X1 npu_inst_pe_1_6_4_U79 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_4_n60), .ZN(npu_inst_pe_1_6_4_n74) );
  OAI21_X1 npu_inst_pe_1_6_4_U78 ( .B1(npu_inst_pe_1_6_4_n63), .B2(
        npu_inst_pe_1_6_4_n60), .A(npu_inst_pe_1_6_4_n74), .ZN(
        npu_inst_pe_1_6_4_n97) );
  NAND2_X1 npu_inst_pe_1_6_4_U77 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_4_n60), .ZN(npu_inst_pe_1_6_4_n73) );
  OAI21_X1 npu_inst_pe_1_6_4_U76 ( .B1(npu_inst_pe_1_6_4_n61), .B2(
        npu_inst_pe_1_6_4_n60), .A(npu_inst_pe_1_6_4_n73), .ZN(
        npu_inst_pe_1_6_4_n96) );
  NAND2_X1 npu_inst_pe_1_6_4_U75 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_4_n56), .ZN(npu_inst_pe_1_6_4_n72) );
  OAI21_X1 npu_inst_pe_1_6_4_U74 ( .B1(npu_inst_pe_1_6_4_n63), .B2(
        npu_inst_pe_1_6_4_n56), .A(npu_inst_pe_1_6_4_n72), .ZN(
        npu_inst_pe_1_6_4_n95) );
  NAND2_X1 npu_inst_pe_1_6_4_U73 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_4_n56), .ZN(npu_inst_pe_1_6_4_n71) );
  OAI21_X1 npu_inst_pe_1_6_4_U72 ( .B1(npu_inst_pe_1_6_4_n61), .B2(
        npu_inst_pe_1_6_4_n56), .A(npu_inst_pe_1_6_4_n71), .ZN(
        npu_inst_pe_1_6_4_n94) );
  NAND2_X1 npu_inst_pe_1_6_4_U71 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_4_n52), .ZN(npu_inst_pe_1_6_4_n70) );
  OAI21_X1 npu_inst_pe_1_6_4_U70 ( .B1(npu_inst_pe_1_6_4_n63), .B2(
        npu_inst_pe_1_6_4_n52), .A(npu_inst_pe_1_6_4_n70), .ZN(
        npu_inst_pe_1_6_4_n93) );
  NAND2_X1 npu_inst_pe_1_6_4_U69 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_4_n52), .ZN(npu_inst_pe_1_6_4_n69) );
  OAI21_X1 npu_inst_pe_1_6_4_U68 ( .B1(npu_inst_pe_1_6_4_n61), .B2(
        npu_inst_pe_1_6_4_n52), .A(npu_inst_pe_1_6_4_n69), .ZN(
        npu_inst_pe_1_6_4_n92) );
  NAND2_X1 npu_inst_pe_1_6_4_U67 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_4_n48), .ZN(npu_inst_pe_1_6_4_n68) );
  OAI21_X1 npu_inst_pe_1_6_4_U66 ( .B1(npu_inst_pe_1_6_4_n63), .B2(
        npu_inst_pe_1_6_4_n48), .A(npu_inst_pe_1_6_4_n68), .ZN(
        npu_inst_pe_1_6_4_n91) );
  NAND2_X1 npu_inst_pe_1_6_4_U65 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_4_n48), .ZN(npu_inst_pe_1_6_4_n67) );
  OAI21_X1 npu_inst_pe_1_6_4_U64 ( .B1(npu_inst_pe_1_6_4_n61), .B2(
        npu_inst_pe_1_6_4_n48), .A(npu_inst_pe_1_6_4_n67), .ZN(
        npu_inst_pe_1_6_4_n90) );
  NAND2_X1 npu_inst_pe_1_6_4_U63 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_4_n44), .ZN(npu_inst_pe_1_6_4_n66) );
  OAI21_X1 npu_inst_pe_1_6_4_U62 ( .B1(npu_inst_pe_1_6_4_n63), .B2(
        npu_inst_pe_1_6_4_n44), .A(npu_inst_pe_1_6_4_n66), .ZN(
        npu_inst_pe_1_6_4_n89) );
  NAND2_X1 npu_inst_pe_1_6_4_U61 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_4_n44), .ZN(npu_inst_pe_1_6_4_n65) );
  OAI21_X1 npu_inst_pe_1_6_4_U60 ( .B1(npu_inst_pe_1_6_4_n61), .B2(
        npu_inst_pe_1_6_4_n44), .A(npu_inst_pe_1_6_4_n65), .ZN(
        npu_inst_pe_1_6_4_n88) );
  NAND2_X1 npu_inst_pe_1_6_4_U59 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_4_n40), .ZN(npu_inst_pe_1_6_4_n64) );
  OAI21_X1 npu_inst_pe_1_6_4_U58 ( .B1(npu_inst_pe_1_6_4_n63), .B2(
        npu_inst_pe_1_6_4_n40), .A(npu_inst_pe_1_6_4_n64), .ZN(
        npu_inst_pe_1_6_4_n87) );
  NAND2_X1 npu_inst_pe_1_6_4_U57 ( .A1(npu_inst_pe_1_6_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_4_n40), .ZN(npu_inst_pe_1_6_4_n62) );
  OAI21_X1 npu_inst_pe_1_6_4_U56 ( .B1(npu_inst_pe_1_6_4_n61), .B2(
        npu_inst_pe_1_6_4_n40), .A(npu_inst_pe_1_6_4_n62), .ZN(
        npu_inst_pe_1_6_4_n86) );
  AOI22_X1 npu_inst_pe_1_6_4_U55 ( .A1(npu_inst_pe_1_6_4_n38), .A2(
        npu_inst_int_data_y_7__4__0_), .B1(npu_inst_pe_1_6_4_n112), .B2(
        npu_inst_pe_1_6_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_4_n37) );
  INV_X1 npu_inst_pe_1_6_4_U54 ( .A(npu_inst_pe_1_6_4_n37), .ZN(
        npu_inst_pe_1_6_4_n111) );
  AND2_X1 npu_inst_pe_1_6_4_U53 ( .A1(npu_inst_n35), .A2(npu_inst_pe_1_6_4_N94), .ZN(npu_inst_int_data_y_6__4__1_) );
  AOI222_X1 npu_inst_pe_1_6_4_U52 ( .A1(npu_inst_int_data_res_7__4__0_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N73), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N65), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n84) );
  INV_X1 npu_inst_pe_1_6_4_U51 ( .A(npu_inst_pe_1_6_4_n84), .ZN(
        npu_inst_pe_1_6_4_n99) );
  AOI222_X1 npu_inst_pe_1_6_4_U50 ( .A1(npu_inst_pe_1_6_4_n1), .A2(
        npu_inst_int_data_res_7__4__7_), .B1(npu_inst_pe_1_6_4_N80), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N72), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n75) );
  INV_X1 npu_inst_pe_1_6_4_U49 ( .A(npu_inst_pe_1_6_4_n75), .ZN(
        npu_inst_pe_1_6_4_n31) );
  AOI222_X1 npu_inst_pe_1_6_4_U48 ( .A1(npu_inst_int_data_res_7__4__1_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N74), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N66), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n83) );
  INV_X1 npu_inst_pe_1_6_4_U47 ( .A(npu_inst_pe_1_6_4_n83), .ZN(
        npu_inst_pe_1_6_4_n98) );
  AOI222_X1 npu_inst_pe_1_6_4_U46 ( .A1(npu_inst_int_data_res_7__4__3_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N76), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N68), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n81) );
  INV_X1 npu_inst_pe_1_6_4_U45 ( .A(npu_inst_pe_1_6_4_n81), .ZN(
        npu_inst_pe_1_6_4_n35) );
  AOI222_X1 npu_inst_pe_1_6_4_U44 ( .A1(npu_inst_int_data_res_7__4__4_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N77), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N69), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n80) );
  INV_X1 npu_inst_pe_1_6_4_U43 ( .A(npu_inst_pe_1_6_4_n80), .ZN(
        npu_inst_pe_1_6_4_n34) );
  AOI222_X1 npu_inst_pe_1_6_4_U42 ( .A1(npu_inst_int_data_res_7__4__5_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N78), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N70), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n79) );
  INV_X1 npu_inst_pe_1_6_4_U41 ( .A(npu_inst_pe_1_6_4_n79), .ZN(
        npu_inst_pe_1_6_4_n33) );
  AOI222_X1 npu_inst_pe_1_6_4_U40 ( .A1(npu_inst_int_data_res_7__4__6_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N79), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N71), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n78) );
  INV_X1 npu_inst_pe_1_6_4_U39 ( .A(npu_inst_pe_1_6_4_n78), .ZN(
        npu_inst_pe_1_6_4_n32) );
  AND2_X1 npu_inst_pe_1_6_4_U38 ( .A1(npu_inst_int_data_x_6__4__1_), .A2(
        npu_inst_pe_1_6_4_int_q_weight_1_), .ZN(npu_inst_pe_1_6_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_4_U37 ( .A1(npu_inst_int_data_x_6__4__0_), .A2(
        npu_inst_pe_1_6_4_int_q_weight_1_), .ZN(npu_inst_pe_1_6_4_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_6_4_U36 ( .A(npu_inst_pe_1_6_4_int_data_1_), .ZN(
        npu_inst_pe_1_6_4_n12) );
  NOR3_X1 npu_inst_pe_1_6_4_U35 ( .A1(npu_inst_pe_1_6_4_n26), .A2(npu_inst_n35), .A3(npu_inst_int_ckg[11]), .ZN(npu_inst_pe_1_6_4_n85) );
  OR2_X1 npu_inst_pe_1_6_4_U34 ( .A1(npu_inst_pe_1_6_4_n85), .A2(
        npu_inst_pe_1_6_4_n1), .ZN(npu_inst_pe_1_6_4_N84) );
  AOI222_X1 npu_inst_pe_1_6_4_U33 ( .A1(npu_inst_int_data_res_7__4__2_), .A2(
        npu_inst_pe_1_6_4_n1), .B1(npu_inst_pe_1_6_4_N75), .B2(
        npu_inst_pe_1_6_4_n76), .C1(npu_inst_pe_1_6_4_N67), .C2(
        npu_inst_pe_1_6_4_n77), .ZN(npu_inst_pe_1_6_4_n82) );
  INV_X1 npu_inst_pe_1_6_4_U32 ( .A(npu_inst_pe_1_6_4_n82), .ZN(
        npu_inst_pe_1_6_4_n36) );
  AOI22_X1 npu_inst_pe_1_6_4_U31 ( .A1(npu_inst_n35), .A2(
        npu_inst_int_data_y_7__4__1_), .B1(npu_inst_pe_1_6_4_n2), .B2(
        npu_inst_int_data_x_6__5__1_), .ZN(npu_inst_pe_1_6_4_n63) );
  AOI22_X1 npu_inst_pe_1_6_4_U30 ( .A1(npu_inst_n35), .A2(
        npu_inst_int_data_y_7__4__0_), .B1(npu_inst_pe_1_6_4_n2), .B2(
        npu_inst_int_data_x_6__5__0_), .ZN(npu_inst_pe_1_6_4_n61) );
  INV_X1 npu_inst_pe_1_6_4_U29 ( .A(npu_inst_pe_1_6_4_int_data_0_), .ZN(
        npu_inst_pe_1_6_4_n11) );
  INV_X1 npu_inst_pe_1_6_4_U28 ( .A(npu_inst_n49), .ZN(npu_inst_pe_1_6_4_n4)
         );
  OR3_X1 npu_inst_pe_1_6_4_U27 ( .A1(npu_inst_n57), .A2(npu_inst_pe_1_6_4_n6), 
        .A3(npu_inst_pe_1_6_4_n4), .ZN(npu_inst_pe_1_6_4_n56) );
  OR3_X1 npu_inst_pe_1_6_4_U26 ( .A1(npu_inst_pe_1_6_4_n4), .A2(
        npu_inst_pe_1_6_4_n6), .A3(npu_inst_pe_1_6_4_n5), .ZN(
        npu_inst_pe_1_6_4_n48) );
  INV_X1 npu_inst_pe_1_6_4_U25 ( .A(npu_inst_pe_1_6_4_n4), .ZN(
        npu_inst_pe_1_6_4_n3) );
  OR3_X1 npu_inst_pe_1_6_4_U24 ( .A1(npu_inst_pe_1_6_4_n3), .A2(
        npu_inst_pe_1_6_4_n6), .A3(npu_inst_pe_1_6_4_n5), .ZN(
        npu_inst_pe_1_6_4_n52) );
  OR3_X1 npu_inst_pe_1_6_4_U23 ( .A1(npu_inst_n57), .A2(npu_inst_pe_1_6_4_n6), 
        .A3(npu_inst_pe_1_6_4_n3), .ZN(npu_inst_pe_1_6_4_n60) );
  BUF_X1 npu_inst_pe_1_6_4_U22 ( .A(npu_inst_n14), .Z(npu_inst_pe_1_6_4_n1) );
  NOR2_X1 npu_inst_pe_1_6_4_U21 ( .A1(npu_inst_pe_1_6_4_n60), .A2(
        npu_inst_pe_1_6_4_n2), .ZN(npu_inst_pe_1_6_4_n58) );
  NOR2_X1 npu_inst_pe_1_6_4_U20 ( .A1(npu_inst_pe_1_6_4_n56), .A2(
        npu_inst_pe_1_6_4_n2), .ZN(npu_inst_pe_1_6_4_n54) );
  NOR2_X1 npu_inst_pe_1_6_4_U19 ( .A1(npu_inst_pe_1_6_4_n52), .A2(
        npu_inst_pe_1_6_4_n2), .ZN(npu_inst_pe_1_6_4_n50) );
  NOR2_X1 npu_inst_pe_1_6_4_U18 ( .A1(npu_inst_pe_1_6_4_n48), .A2(
        npu_inst_pe_1_6_4_n2), .ZN(npu_inst_pe_1_6_4_n46) );
  NOR2_X1 npu_inst_pe_1_6_4_U17 ( .A1(npu_inst_pe_1_6_4_n40), .A2(
        npu_inst_pe_1_6_4_n2), .ZN(npu_inst_pe_1_6_4_n38) );
  NOR2_X1 npu_inst_pe_1_6_4_U16 ( .A1(npu_inst_pe_1_6_4_n44), .A2(
        npu_inst_pe_1_6_4_n2), .ZN(npu_inst_pe_1_6_4_n42) );
  BUF_X1 npu_inst_pe_1_6_4_U15 ( .A(npu_inst_n76), .Z(npu_inst_pe_1_6_4_n6) );
  INV_X1 npu_inst_pe_1_6_4_U14 ( .A(npu_inst_n104), .ZN(npu_inst_pe_1_6_4_n10)
         );
  INV_X1 npu_inst_pe_1_6_4_U13 ( .A(npu_inst_pe_1_6_4_n38), .ZN(
        npu_inst_pe_1_6_4_n112) );
  INV_X1 npu_inst_pe_1_6_4_U12 ( .A(npu_inst_pe_1_6_4_n58), .ZN(
        npu_inst_pe_1_6_4_n117) );
  INV_X1 npu_inst_pe_1_6_4_U11 ( .A(npu_inst_pe_1_6_4_n54), .ZN(
        npu_inst_pe_1_6_4_n116) );
  INV_X1 npu_inst_pe_1_6_4_U10 ( .A(npu_inst_pe_1_6_4_n50), .ZN(
        npu_inst_pe_1_6_4_n115) );
  INV_X1 npu_inst_pe_1_6_4_U9 ( .A(npu_inst_pe_1_6_4_n46), .ZN(
        npu_inst_pe_1_6_4_n114) );
  INV_X1 npu_inst_pe_1_6_4_U8 ( .A(npu_inst_pe_1_6_4_n42), .ZN(
        npu_inst_pe_1_6_4_n113) );
  BUF_X1 npu_inst_pe_1_6_4_U7 ( .A(npu_inst_pe_1_6_4_n10), .Z(
        npu_inst_pe_1_6_4_n9) );
  BUF_X1 npu_inst_pe_1_6_4_U6 ( .A(npu_inst_pe_1_6_4_n10), .Z(
        npu_inst_pe_1_6_4_n8) );
  BUF_X1 npu_inst_pe_1_6_4_U5 ( .A(npu_inst_pe_1_6_4_n10), .Z(
        npu_inst_pe_1_6_4_n7) );
  NOR2_X1 npu_inst_pe_1_6_4_U4 ( .A1(npu_inst_pe_1_6_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_4_n1), .ZN(npu_inst_pe_1_6_4_n76) );
  NOR2_X1 npu_inst_pe_1_6_4_U3 ( .A1(npu_inst_pe_1_6_4_n27), .A2(
        npu_inst_pe_1_6_4_n1), .ZN(npu_inst_pe_1_6_4_n77) );
  FA_X1 npu_inst_pe_1_6_4_sub_77_U2_1 ( .A(npu_inst_int_data_res_6__4__1_), 
        .B(npu_inst_pe_1_6_4_n12), .CI(npu_inst_pe_1_6_4_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_6_4_sub_77_carry_2_), .S(npu_inst_pe_1_6_4_N66) );
  FA_X1 npu_inst_pe_1_6_4_add_79_U1_1 ( .A(npu_inst_int_data_res_6__4__1_), 
        .B(npu_inst_pe_1_6_4_int_data_1_), .CI(
        npu_inst_pe_1_6_4_add_79_carry_1_), .CO(
        npu_inst_pe_1_6_4_add_79_carry_2_), .S(npu_inst_pe_1_6_4_N74) );
  NAND3_X1 npu_inst_pe_1_6_4_U101 ( .A1(npu_inst_pe_1_6_4_n4), .A2(
        npu_inst_pe_1_6_4_n5), .A3(npu_inst_pe_1_6_4_n6), .ZN(
        npu_inst_pe_1_6_4_n44) );
  NAND3_X1 npu_inst_pe_1_6_4_U100 ( .A1(npu_inst_pe_1_6_4_n3), .A2(
        npu_inst_pe_1_6_4_n5), .A3(npu_inst_pe_1_6_4_n6), .ZN(
        npu_inst_pe_1_6_4_n40) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_4_n32), .CK(
        npu_inst_pe_1_6_4_net3282), .RN(npu_inst_pe_1_6_4_n7), .Q(
        npu_inst_int_data_res_6__4__6_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_4_n33), .CK(
        npu_inst_pe_1_6_4_net3282), .RN(npu_inst_pe_1_6_4_n7), .Q(
        npu_inst_int_data_res_6__4__5_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_4_n34), .CK(
        npu_inst_pe_1_6_4_net3282), .RN(npu_inst_pe_1_6_4_n7), .Q(
        npu_inst_int_data_res_6__4__4_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_4_n35), .CK(
        npu_inst_pe_1_6_4_net3282), .RN(npu_inst_pe_1_6_4_n7), .Q(
        npu_inst_int_data_res_6__4__3_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_4_n36), .CK(
        npu_inst_pe_1_6_4_net3282), .RN(npu_inst_pe_1_6_4_n7), .Q(
        npu_inst_int_data_res_6__4__2_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_4_n98), .CK(
        npu_inst_pe_1_6_4_net3282), .RN(npu_inst_pe_1_6_4_n7), .Q(
        npu_inst_int_data_res_6__4__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_4_n31), .CK(
        npu_inst_pe_1_6_4_net3282), .RN(npu_inst_pe_1_6_4_n7), .Q(
        npu_inst_int_data_res_6__4__7_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_4_n99), .CK(
        npu_inst_pe_1_6_4_net3282), .RN(npu_inst_pe_1_6_4_n7), .Q(
        npu_inst_int_data_res_6__4__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_weight_reg_0_ ( .D(npu_inst_n90), .CK(
        npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n7), .Q(
        npu_inst_pe_1_6_4_int_q_weight_0_), .QN(npu_inst_pe_1_6_4_n27) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_weight_reg_1_ ( .D(npu_inst_n96), .CK(
        npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n7), .Q(
        npu_inst_pe_1_6_4_int_q_weight_1_), .QN(npu_inst_pe_1_6_4_n26) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_4_n111), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n7), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_4_n105), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n7), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_4_n110), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_4_n104), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_4_n109), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_4_n103), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_4_n108), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_4_n102), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_4_n107), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_4_n101), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_4_n106), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_4_n100), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_4_n86), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_4_n87), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n8), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_4_n88), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_4_n89), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_4_n90), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_4_n91), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_4_n92), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_4_n93), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_4_n94), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_4_n95), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_4_n96), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_4_n97), 
        .CK(npu_inst_pe_1_6_4_net3288), .RN(npu_inst_pe_1_6_4_n9), .Q(
        npu_inst_pe_1_6_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_4_net3282) );
  CLKGATETST_X1 npu_inst_pe_1_6_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n44), .SE(1'b0), .GCK(npu_inst_pe_1_6_4_net3288) );
  MUX2_X1 npu_inst_pe_1_6_5_U153 ( .A(npu_inst_pe_1_6_5_n31), .B(
        npu_inst_pe_1_6_5_n28), .S(npu_inst_pe_1_6_5_n7), .Z(
        npu_inst_pe_1_6_5_N93) );
  MUX2_X1 npu_inst_pe_1_6_5_U152 ( .A(npu_inst_pe_1_6_5_n30), .B(
        npu_inst_pe_1_6_5_n29), .S(npu_inst_pe_1_6_5_n5), .Z(
        npu_inst_pe_1_6_5_n31) );
  MUX2_X1 npu_inst_pe_1_6_5_U151 ( .A(npu_inst_pe_1_6_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_5_n3), .Z(
        npu_inst_pe_1_6_5_n30) );
  MUX2_X1 npu_inst_pe_1_6_5_U150 ( .A(npu_inst_pe_1_6_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_5_n3), .Z(
        npu_inst_pe_1_6_5_n29) );
  MUX2_X1 npu_inst_pe_1_6_5_U149 ( .A(npu_inst_pe_1_6_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_5_n3), .Z(
        npu_inst_pe_1_6_5_n28) );
  MUX2_X1 npu_inst_pe_1_6_5_U148 ( .A(npu_inst_pe_1_6_5_n25), .B(
        npu_inst_pe_1_6_5_n22), .S(npu_inst_pe_1_6_5_n7), .Z(
        npu_inst_pe_1_6_5_N94) );
  MUX2_X1 npu_inst_pe_1_6_5_U147 ( .A(npu_inst_pe_1_6_5_n24), .B(
        npu_inst_pe_1_6_5_n23), .S(npu_inst_pe_1_6_5_n5), .Z(
        npu_inst_pe_1_6_5_n25) );
  MUX2_X1 npu_inst_pe_1_6_5_U146 ( .A(npu_inst_pe_1_6_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_5_n3), .Z(
        npu_inst_pe_1_6_5_n24) );
  MUX2_X1 npu_inst_pe_1_6_5_U145 ( .A(npu_inst_pe_1_6_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_5_n3), .Z(
        npu_inst_pe_1_6_5_n23) );
  MUX2_X1 npu_inst_pe_1_6_5_U144 ( .A(npu_inst_pe_1_6_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_5_n3), .Z(
        npu_inst_pe_1_6_5_n22) );
  MUX2_X1 npu_inst_pe_1_6_5_U143 ( .A(npu_inst_pe_1_6_5_n21), .B(
        npu_inst_pe_1_6_5_n18), .S(npu_inst_pe_1_6_5_n7), .Z(
        npu_inst_int_data_x_6__5__1_) );
  MUX2_X1 npu_inst_pe_1_6_5_U142 ( .A(npu_inst_pe_1_6_5_n20), .B(
        npu_inst_pe_1_6_5_n19), .S(npu_inst_pe_1_6_5_n5), .Z(
        npu_inst_pe_1_6_5_n21) );
  MUX2_X1 npu_inst_pe_1_6_5_U141 ( .A(npu_inst_pe_1_6_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_5_n3), .Z(
        npu_inst_pe_1_6_5_n20) );
  MUX2_X1 npu_inst_pe_1_6_5_U140 ( .A(npu_inst_pe_1_6_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_5_n3), .Z(
        npu_inst_pe_1_6_5_n19) );
  MUX2_X1 npu_inst_pe_1_6_5_U139 ( .A(npu_inst_pe_1_6_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_5_n3), .Z(
        npu_inst_pe_1_6_5_n18) );
  MUX2_X1 npu_inst_pe_1_6_5_U138 ( .A(npu_inst_pe_1_6_5_n17), .B(
        npu_inst_pe_1_6_5_n14), .S(npu_inst_pe_1_6_5_n7), .Z(
        npu_inst_int_data_x_6__5__0_) );
  MUX2_X1 npu_inst_pe_1_6_5_U137 ( .A(npu_inst_pe_1_6_5_n16), .B(
        npu_inst_pe_1_6_5_n15), .S(npu_inst_pe_1_6_5_n5), .Z(
        npu_inst_pe_1_6_5_n17) );
  MUX2_X1 npu_inst_pe_1_6_5_U136 ( .A(npu_inst_pe_1_6_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_5_n3), .Z(
        npu_inst_pe_1_6_5_n16) );
  MUX2_X1 npu_inst_pe_1_6_5_U135 ( .A(npu_inst_pe_1_6_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_5_n3), .Z(
        npu_inst_pe_1_6_5_n15) );
  MUX2_X1 npu_inst_pe_1_6_5_U134 ( .A(npu_inst_pe_1_6_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_5_n3), .Z(
        npu_inst_pe_1_6_5_n14) );
  XOR2_X1 npu_inst_pe_1_6_5_U133 ( .A(npu_inst_pe_1_6_5_int_data_0_), .B(
        npu_inst_int_data_res_6__5__0_), .Z(npu_inst_pe_1_6_5_N73) );
  AND2_X1 npu_inst_pe_1_6_5_U132 ( .A1(npu_inst_int_data_res_6__5__0_), .A2(
        npu_inst_pe_1_6_5_int_data_0_), .ZN(npu_inst_pe_1_6_5_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_5_U131 ( .A(npu_inst_int_data_res_6__5__0_), .B(
        npu_inst_pe_1_6_5_n12), .ZN(npu_inst_pe_1_6_5_N65) );
  OR2_X1 npu_inst_pe_1_6_5_U130 ( .A1(npu_inst_pe_1_6_5_n12), .A2(
        npu_inst_int_data_res_6__5__0_), .ZN(npu_inst_pe_1_6_5_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_5_U129 ( .A(npu_inst_int_data_res_6__5__2_), .B(
        npu_inst_pe_1_6_5_add_79_carry_2_), .Z(npu_inst_pe_1_6_5_N75) );
  AND2_X1 npu_inst_pe_1_6_5_U128 ( .A1(npu_inst_pe_1_6_5_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_6__5__2_), .ZN(
        npu_inst_pe_1_6_5_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_5_U127 ( .A(npu_inst_int_data_res_6__5__3_), .B(
        npu_inst_pe_1_6_5_add_79_carry_3_), .Z(npu_inst_pe_1_6_5_N76) );
  AND2_X1 npu_inst_pe_1_6_5_U126 ( .A1(npu_inst_pe_1_6_5_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_6__5__3_), .ZN(
        npu_inst_pe_1_6_5_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_5_U125 ( .A(npu_inst_int_data_res_6__5__4_), .B(
        npu_inst_pe_1_6_5_add_79_carry_4_), .Z(npu_inst_pe_1_6_5_N77) );
  AND2_X1 npu_inst_pe_1_6_5_U124 ( .A1(npu_inst_pe_1_6_5_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_6__5__4_), .ZN(
        npu_inst_pe_1_6_5_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_5_U123 ( .A(npu_inst_int_data_res_6__5__5_), .B(
        npu_inst_pe_1_6_5_add_79_carry_5_), .Z(npu_inst_pe_1_6_5_N78) );
  AND2_X1 npu_inst_pe_1_6_5_U122 ( .A1(npu_inst_pe_1_6_5_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_6__5__5_), .ZN(
        npu_inst_pe_1_6_5_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_5_U121 ( .A(npu_inst_int_data_res_6__5__6_), .B(
        npu_inst_pe_1_6_5_add_79_carry_6_), .Z(npu_inst_pe_1_6_5_N79) );
  AND2_X1 npu_inst_pe_1_6_5_U120 ( .A1(npu_inst_pe_1_6_5_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_6__5__6_), .ZN(
        npu_inst_pe_1_6_5_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_5_U119 ( .A(npu_inst_int_data_res_6__5__7_), .B(
        npu_inst_pe_1_6_5_add_79_carry_7_), .Z(npu_inst_pe_1_6_5_N80) );
  XNOR2_X1 npu_inst_pe_1_6_5_U118 ( .A(npu_inst_pe_1_6_5_sub_77_carry_2_), .B(
        npu_inst_int_data_res_6__5__2_), .ZN(npu_inst_pe_1_6_5_N67) );
  OR2_X1 npu_inst_pe_1_6_5_U117 ( .A1(npu_inst_int_data_res_6__5__2_), .A2(
        npu_inst_pe_1_6_5_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_6_5_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_5_U116 ( .A(npu_inst_pe_1_6_5_sub_77_carry_3_), .B(
        npu_inst_int_data_res_6__5__3_), .ZN(npu_inst_pe_1_6_5_N68) );
  OR2_X1 npu_inst_pe_1_6_5_U115 ( .A1(npu_inst_int_data_res_6__5__3_), .A2(
        npu_inst_pe_1_6_5_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_6_5_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_5_U114 ( .A(npu_inst_pe_1_6_5_sub_77_carry_4_), .B(
        npu_inst_int_data_res_6__5__4_), .ZN(npu_inst_pe_1_6_5_N69) );
  OR2_X1 npu_inst_pe_1_6_5_U113 ( .A1(npu_inst_int_data_res_6__5__4_), .A2(
        npu_inst_pe_1_6_5_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_6_5_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_5_U112 ( .A(npu_inst_pe_1_6_5_sub_77_carry_5_), .B(
        npu_inst_int_data_res_6__5__5_), .ZN(npu_inst_pe_1_6_5_N70) );
  OR2_X1 npu_inst_pe_1_6_5_U111 ( .A1(npu_inst_int_data_res_6__5__5_), .A2(
        npu_inst_pe_1_6_5_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_6_5_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_5_U110 ( .A(npu_inst_pe_1_6_5_sub_77_carry_6_), .B(
        npu_inst_int_data_res_6__5__6_), .ZN(npu_inst_pe_1_6_5_N71) );
  OR2_X1 npu_inst_pe_1_6_5_U109 ( .A1(npu_inst_int_data_res_6__5__6_), .A2(
        npu_inst_pe_1_6_5_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_6_5_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_5_U108 ( .A(npu_inst_int_data_res_6__5__7_), .B(
        npu_inst_pe_1_6_5_sub_77_carry_7_), .ZN(npu_inst_pe_1_6_5_N72) );
  INV_X1 npu_inst_pe_1_6_5_U107 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_6_5_n6)
         );
  INV_X1 npu_inst_pe_1_6_5_U106 ( .A(npu_inst_pe_1_6_5_n6), .ZN(
        npu_inst_pe_1_6_5_n5) );
  INV_X1 npu_inst_pe_1_6_5_U105 ( .A(npu_inst_n35), .ZN(npu_inst_pe_1_6_5_n2)
         );
  AOI22_X1 npu_inst_pe_1_6_5_U104 ( .A1(npu_inst_int_data_y_7__5__0_), .A2(
        npu_inst_pe_1_6_5_n58), .B1(npu_inst_pe_1_6_5_n118), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_5_n57) );
  INV_X1 npu_inst_pe_1_6_5_U103 ( .A(npu_inst_pe_1_6_5_n57), .ZN(
        npu_inst_pe_1_6_5_n107) );
  AOI22_X1 npu_inst_pe_1_6_5_U102 ( .A1(npu_inst_int_data_y_7__5__0_), .A2(
        npu_inst_pe_1_6_5_n54), .B1(npu_inst_pe_1_6_5_n117), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_5_n53) );
  INV_X1 npu_inst_pe_1_6_5_U99 ( .A(npu_inst_pe_1_6_5_n53), .ZN(
        npu_inst_pe_1_6_5_n108) );
  AOI22_X1 npu_inst_pe_1_6_5_U98 ( .A1(npu_inst_int_data_y_7__5__0_), .A2(
        npu_inst_pe_1_6_5_n50), .B1(npu_inst_pe_1_6_5_n116), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_5_n49) );
  INV_X1 npu_inst_pe_1_6_5_U97 ( .A(npu_inst_pe_1_6_5_n49), .ZN(
        npu_inst_pe_1_6_5_n109) );
  AOI22_X1 npu_inst_pe_1_6_5_U96 ( .A1(npu_inst_int_data_y_7__5__0_), .A2(
        npu_inst_pe_1_6_5_n46), .B1(npu_inst_pe_1_6_5_n115), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_5_n45) );
  INV_X1 npu_inst_pe_1_6_5_U95 ( .A(npu_inst_pe_1_6_5_n45), .ZN(
        npu_inst_pe_1_6_5_n110) );
  AOI22_X1 npu_inst_pe_1_6_5_U94 ( .A1(npu_inst_int_data_y_7__5__0_), .A2(
        npu_inst_pe_1_6_5_n42), .B1(npu_inst_pe_1_6_5_n114), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_5_n41) );
  INV_X1 npu_inst_pe_1_6_5_U93 ( .A(npu_inst_pe_1_6_5_n41), .ZN(
        npu_inst_pe_1_6_5_n111) );
  AOI22_X1 npu_inst_pe_1_6_5_U92 ( .A1(npu_inst_int_data_y_7__5__1_), .A2(
        npu_inst_pe_1_6_5_n58), .B1(npu_inst_pe_1_6_5_n118), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_5_n59) );
  INV_X1 npu_inst_pe_1_6_5_U91 ( .A(npu_inst_pe_1_6_5_n59), .ZN(
        npu_inst_pe_1_6_5_n101) );
  AOI22_X1 npu_inst_pe_1_6_5_U90 ( .A1(npu_inst_int_data_y_7__5__1_), .A2(
        npu_inst_pe_1_6_5_n54), .B1(npu_inst_pe_1_6_5_n117), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_5_n55) );
  INV_X1 npu_inst_pe_1_6_5_U89 ( .A(npu_inst_pe_1_6_5_n55), .ZN(
        npu_inst_pe_1_6_5_n102) );
  AOI22_X1 npu_inst_pe_1_6_5_U88 ( .A1(npu_inst_int_data_y_7__5__1_), .A2(
        npu_inst_pe_1_6_5_n50), .B1(npu_inst_pe_1_6_5_n116), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_5_n51) );
  INV_X1 npu_inst_pe_1_6_5_U87 ( .A(npu_inst_pe_1_6_5_n51), .ZN(
        npu_inst_pe_1_6_5_n103) );
  AOI22_X1 npu_inst_pe_1_6_5_U86 ( .A1(npu_inst_int_data_y_7__5__1_), .A2(
        npu_inst_pe_1_6_5_n46), .B1(npu_inst_pe_1_6_5_n115), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_5_n47) );
  INV_X1 npu_inst_pe_1_6_5_U85 ( .A(npu_inst_pe_1_6_5_n47), .ZN(
        npu_inst_pe_1_6_5_n104) );
  AOI22_X1 npu_inst_pe_1_6_5_U84 ( .A1(npu_inst_int_data_y_7__5__1_), .A2(
        npu_inst_pe_1_6_5_n42), .B1(npu_inst_pe_1_6_5_n114), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_5_n43) );
  INV_X1 npu_inst_pe_1_6_5_U83 ( .A(npu_inst_pe_1_6_5_n43), .ZN(
        npu_inst_pe_1_6_5_n105) );
  AOI22_X1 npu_inst_pe_1_6_5_U82 ( .A1(npu_inst_pe_1_6_5_n38), .A2(
        npu_inst_int_data_y_7__5__1_), .B1(npu_inst_pe_1_6_5_n113), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_5_n39) );
  INV_X1 npu_inst_pe_1_6_5_U81 ( .A(npu_inst_pe_1_6_5_n39), .ZN(
        npu_inst_pe_1_6_5_n106) );
  AND2_X1 npu_inst_pe_1_6_5_U80 ( .A1(npu_inst_pe_1_6_5_N93), .A2(npu_inst_n35), .ZN(npu_inst_int_data_y_6__5__0_) );
  NAND2_X1 npu_inst_pe_1_6_5_U79 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_5_n60), .ZN(npu_inst_pe_1_6_5_n74) );
  OAI21_X1 npu_inst_pe_1_6_5_U78 ( .B1(npu_inst_pe_1_6_5_n63), .B2(
        npu_inst_pe_1_6_5_n60), .A(npu_inst_pe_1_6_5_n74), .ZN(
        npu_inst_pe_1_6_5_n97) );
  NAND2_X1 npu_inst_pe_1_6_5_U77 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_5_n60), .ZN(npu_inst_pe_1_6_5_n73) );
  OAI21_X1 npu_inst_pe_1_6_5_U76 ( .B1(npu_inst_pe_1_6_5_n61), .B2(
        npu_inst_pe_1_6_5_n60), .A(npu_inst_pe_1_6_5_n73), .ZN(
        npu_inst_pe_1_6_5_n96) );
  NAND2_X1 npu_inst_pe_1_6_5_U75 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_5_n56), .ZN(npu_inst_pe_1_6_5_n72) );
  OAI21_X1 npu_inst_pe_1_6_5_U74 ( .B1(npu_inst_pe_1_6_5_n63), .B2(
        npu_inst_pe_1_6_5_n56), .A(npu_inst_pe_1_6_5_n72), .ZN(
        npu_inst_pe_1_6_5_n95) );
  NAND2_X1 npu_inst_pe_1_6_5_U73 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_5_n56), .ZN(npu_inst_pe_1_6_5_n71) );
  OAI21_X1 npu_inst_pe_1_6_5_U72 ( .B1(npu_inst_pe_1_6_5_n61), .B2(
        npu_inst_pe_1_6_5_n56), .A(npu_inst_pe_1_6_5_n71), .ZN(
        npu_inst_pe_1_6_5_n94) );
  NAND2_X1 npu_inst_pe_1_6_5_U71 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_5_n52), .ZN(npu_inst_pe_1_6_5_n70) );
  OAI21_X1 npu_inst_pe_1_6_5_U70 ( .B1(npu_inst_pe_1_6_5_n63), .B2(
        npu_inst_pe_1_6_5_n52), .A(npu_inst_pe_1_6_5_n70), .ZN(
        npu_inst_pe_1_6_5_n93) );
  NAND2_X1 npu_inst_pe_1_6_5_U69 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_5_n52), .ZN(npu_inst_pe_1_6_5_n69) );
  OAI21_X1 npu_inst_pe_1_6_5_U68 ( .B1(npu_inst_pe_1_6_5_n61), .B2(
        npu_inst_pe_1_6_5_n52), .A(npu_inst_pe_1_6_5_n69), .ZN(
        npu_inst_pe_1_6_5_n92) );
  NAND2_X1 npu_inst_pe_1_6_5_U67 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_5_n48), .ZN(npu_inst_pe_1_6_5_n68) );
  OAI21_X1 npu_inst_pe_1_6_5_U66 ( .B1(npu_inst_pe_1_6_5_n63), .B2(
        npu_inst_pe_1_6_5_n48), .A(npu_inst_pe_1_6_5_n68), .ZN(
        npu_inst_pe_1_6_5_n91) );
  NAND2_X1 npu_inst_pe_1_6_5_U65 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_5_n48), .ZN(npu_inst_pe_1_6_5_n67) );
  OAI21_X1 npu_inst_pe_1_6_5_U64 ( .B1(npu_inst_pe_1_6_5_n61), .B2(
        npu_inst_pe_1_6_5_n48), .A(npu_inst_pe_1_6_5_n67), .ZN(
        npu_inst_pe_1_6_5_n90) );
  NAND2_X1 npu_inst_pe_1_6_5_U63 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_5_n44), .ZN(npu_inst_pe_1_6_5_n66) );
  OAI21_X1 npu_inst_pe_1_6_5_U62 ( .B1(npu_inst_pe_1_6_5_n63), .B2(
        npu_inst_pe_1_6_5_n44), .A(npu_inst_pe_1_6_5_n66), .ZN(
        npu_inst_pe_1_6_5_n89) );
  NAND2_X1 npu_inst_pe_1_6_5_U61 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_5_n44), .ZN(npu_inst_pe_1_6_5_n65) );
  OAI21_X1 npu_inst_pe_1_6_5_U60 ( .B1(npu_inst_pe_1_6_5_n61), .B2(
        npu_inst_pe_1_6_5_n44), .A(npu_inst_pe_1_6_5_n65), .ZN(
        npu_inst_pe_1_6_5_n88) );
  NAND2_X1 npu_inst_pe_1_6_5_U59 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_5_n40), .ZN(npu_inst_pe_1_6_5_n64) );
  OAI21_X1 npu_inst_pe_1_6_5_U58 ( .B1(npu_inst_pe_1_6_5_n63), .B2(
        npu_inst_pe_1_6_5_n40), .A(npu_inst_pe_1_6_5_n64), .ZN(
        npu_inst_pe_1_6_5_n87) );
  NAND2_X1 npu_inst_pe_1_6_5_U57 ( .A1(npu_inst_pe_1_6_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_5_n40), .ZN(npu_inst_pe_1_6_5_n62) );
  OAI21_X1 npu_inst_pe_1_6_5_U56 ( .B1(npu_inst_pe_1_6_5_n61), .B2(
        npu_inst_pe_1_6_5_n40), .A(npu_inst_pe_1_6_5_n62), .ZN(
        npu_inst_pe_1_6_5_n86) );
  AOI22_X1 npu_inst_pe_1_6_5_U55 ( .A1(npu_inst_pe_1_6_5_n38), .A2(
        npu_inst_int_data_y_7__5__0_), .B1(npu_inst_pe_1_6_5_n113), .B2(
        npu_inst_pe_1_6_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_5_n37) );
  INV_X1 npu_inst_pe_1_6_5_U54 ( .A(npu_inst_pe_1_6_5_n37), .ZN(
        npu_inst_pe_1_6_5_n112) );
  AND2_X1 npu_inst_pe_1_6_5_U53 ( .A1(npu_inst_n35), .A2(npu_inst_pe_1_6_5_N94), .ZN(npu_inst_int_data_y_6__5__1_) );
  AOI222_X1 npu_inst_pe_1_6_5_U52 ( .A1(npu_inst_int_data_res_7__5__0_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N73), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N65), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n84) );
  INV_X1 npu_inst_pe_1_6_5_U51 ( .A(npu_inst_pe_1_6_5_n84), .ZN(
        npu_inst_pe_1_6_5_n100) );
  AOI222_X1 npu_inst_pe_1_6_5_U50 ( .A1(npu_inst_pe_1_6_5_n1), .A2(
        npu_inst_int_data_res_7__5__7_), .B1(npu_inst_pe_1_6_5_N80), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N72), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n75) );
  INV_X1 npu_inst_pe_1_6_5_U49 ( .A(npu_inst_pe_1_6_5_n75), .ZN(
        npu_inst_pe_1_6_5_n32) );
  AOI222_X1 npu_inst_pe_1_6_5_U48 ( .A1(npu_inst_int_data_res_7__5__1_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N74), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N66), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n83) );
  INV_X1 npu_inst_pe_1_6_5_U47 ( .A(npu_inst_pe_1_6_5_n83), .ZN(
        npu_inst_pe_1_6_5_n99) );
  AOI222_X1 npu_inst_pe_1_6_5_U46 ( .A1(npu_inst_int_data_res_7__5__3_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N76), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N68), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n81) );
  INV_X1 npu_inst_pe_1_6_5_U45 ( .A(npu_inst_pe_1_6_5_n81), .ZN(
        npu_inst_pe_1_6_5_n36) );
  AOI222_X1 npu_inst_pe_1_6_5_U44 ( .A1(npu_inst_int_data_res_7__5__4_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N77), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N69), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n80) );
  INV_X1 npu_inst_pe_1_6_5_U43 ( .A(npu_inst_pe_1_6_5_n80), .ZN(
        npu_inst_pe_1_6_5_n35) );
  AOI222_X1 npu_inst_pe_1_6_5_U42 ( .A1(npu_inst_int_data_res_7__5__5_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N78), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N70), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n79) );
  INV_X1 npu_inst_pe_1_6_5_U41 ( .A(npu_inst_pe_1_6_5_n79), .ZN(
        npu_inst_pe_1_6_5_n34) );
  AOI222_X1 npu_inst_pe_1_6_5_U40 ( .A1(npu_inst_int_data_res_7__5__6_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N79), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N71), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n78) );
  INV_X1 npu_inst_pe_1_6_5_U39 ( .A(npu_inst_pe_1_6_5_n78), .ZN(
        npu_inst_pe_1_6_5_n33) );
  AND2_X1 npu_inst_pe_1_6_5_U38 ( .A1(npu_inst_int_data_x_6__5__1_), .A2(
        npu_inst_pe_1_6_5_int_q_weight_1_), .ZN(npu_inst_pe_1_6_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_5_U37 ( .A1(npu_inst_int_data_x_6__5__0_), .A2(
        npu_inst_pe_1_6_5_int_q_weight_1_), .ZN(npu_inst_pe_1_6_5_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_6_5_U36 ( .A(npu_inst_pe_1_6_5_int_data_1_), .ZN(
        npu_inst_pe_1_6_5_n13) );
  NOR3_X1 npu_inst_pe_1_6_5_U35 ( .A1(npu_inst_pe_1_6_5_n26), .A2(npu_inst_n35), .A3(npu_inst_int_ckg[10]), .ZN(npu_inst_pe_1_6_5_n85) );
  OR2_X1 npu_inst_pe_1_6_5_U34 ( .A1(npu_inst_pe_1_6_5_n85), .A2(
        npu_inst_pe_1_6_5_n1), .ZN(npu_inst_pe_1_6_5_N84) );
  AOI222_X1 npu_inst_pe_1_6_5_U33 ( .A1(npu_inst_int_data_res_7__5__2_), .A2(
        npu_inst_pe_1_6_5_n1), .B1(npu_inst_pe_1_6_5_N75), .B2(
        npu_inst_pe_1_6_5_n76), .C1(npu_inst_pe_1_6_5_N67), .C2(
        npu_inst_pe_1_6_5_n77), .ZN(npu_inst_pe_1_6_5_n82) );
  INV_X1 npu_inst_pe_1_6_5_U32 ( .A(npu_inst_pe_1_6_5_n82), .ZN(
        npu_inst_pe_1_6_5_n98) );
  AOI22_X1 npu_inst_pe_1_6_5_U31 ( .A1(npu_inst_n35), .A2(
        npu_inst_int_data_y_7__5__1_), .B1(npu_inst_pe_1_6_5_n2), .B2(
        npu_inst_int_data_x_6__6__1_), .ZN(npu_inst_pe_1_6_5_n63) );
  AOI22_X1 npu_inst_pe_1_6_5_U30 ( .A1(npu_inst_n35), .A2(
        npu_inst_int_data_y_7__5__0_), .B1(npu_inst_pe_1_6_5_n2), .B2(
        npu_inst_int_data_x_6__6__0_), .ZN(npu_inst_pe_1_6_5_n61) );
  INV_X1 npu_inst_pe_1_6_5_U29 ( .A(npu_inst_pe_1_6_5_int_data_0_), .ZN(
        npu_inst_pe_1_6_5_n12) );
  INV_X1 npu_inst_pe_1_6_5_U28 ( .A(npu_inst_n49), .ZN(npu_inst_pe_1_6_5_n4)
         );
  OR3_X1 npu_inst_pe_1_6_5_U27 ( .A1(npu_inst_pe_1_6_5_n5), .A2(
        npu_inst_pe_1_6_5_n7), .A3(npu_inst_pe_1_6_5_n4), .ZN(
        npu_inst_pe_1_6_5_n56) );
  OR3_X1 npu_inst_pe_1_6_5_U26 ( .A1(npu_inst_pe_1_6_5_n4), .A2(
        npu_inst_pe_1_6_5_n7), .A3(npu_inst_pe_1_6_5_n6), .ZN(
        npu_inst_pe_1_6_5_n48) );
  INV_X1 npu_inst_pe_1_6_5_U25 ( .A(npu_inst_pe_1_6_5_n4), .ZN(
        npu_inst_pe_1_6_5_n3) );
  OR3_X1 npu_inst_pe_1_6_5_U24 ( .A1(npu_inst_pe_1_6_5_n3), .A2(
        npu_inst_pe_1_6_5_n7), .A3(npu_inst_pe_1_6_5_n6), .ZN(
        npu_inst_pe_1_6_5_n52) );
  OR3_X1 npu_inst_pe_1_6_5_U23 ( .A1(npu_inst_pe_1_6_5_n5), .A2(
        npu_inst_pe_1_6_5_n7), .A3(npu_inst_pe_1_6_5_n3), .ZN(
        npu_inst_pe_1_6_5_n60) );
  BUF_X1 npu_inst_pe_1_6_5_U22 ( .A(npu_inst_n14), .Z(npu_inst_pe_1_6_5_n1) );
  NOR2_X1 npu_inst_pe_1_6_5_U21 ( .A1(npu_inst_pe_1_6_5_n60), .A2(
        npu_inst_pe_1_6_5_n2), .ZN(npu_inst_pe_1_6_5_n58) );
  NOR2_X1 npu_inst_pe_1_6_5_U20 ( .A1(npu_inst_pe_1_6_5_n56), .A2(
        npu_inst_pe_1_6_5_n2), .ZN(npu_inst_pe_1_6_5_n54) );
  NOR2_X1 npu_inst_pe_1_6_5_U19 ( .A1(npu_inst_pe_1_6_5_n52), .A2(
        npu_inst_pe_1_6_5_n2), .ZN(npu_inst_pe_1_6_5_n50) );
  NOR2_X1 npu_inst_pe_1_6_5_U18 ( .A1(npu_inst_pe_1_6_5_n48), .A2(
        npu_inst_pe_1_6_5_n2), .ZN(npu_inst_pe_1_6_5_n46) );
  NOR2_X1 npu_inst_pe_1_6_5_U17 ( .A1(npu_inst_pe_1_6_5_n40), .A2(
        npu_inst_pe_1_6_5_n2), .ZN(npu_inst_pe_1_6_5_n38) );
  NOR2_X1 npu_inst_pe_1_6_5_U16 ( .A1(npu_inst_pe_1_6_5_n44), .A2(
        npu_inst_pe_1_6_5_n2), .ZN(npu_inst_pe_1_6_5_n42) );
  BUF_X1 npu_inst_pe_1_6_5_U15 ( .A(npu_inst_n76), .Z(npu_inst_pe_1_6_5_n7) );
  INV_X1 npu_inst_pe_1_6_5_U14 ( .A(npu_inst_n104), .ZN(npu_inst_pe_1_6_5_n11)
         );
  INV_X1 npu_inst_pe_1_6_5_U13 ( .A(npu_inst_pe_1_6_5_n38), .ZN(
        npu_inst_pe_1_6_5_n113) );
  INV_X1 npu_inst_pe_1_6_5_U12 ( .A(npu_inst_pe_1_6_5_n58), .ZN(
        npu_inst_pe_1_6_5_n118) );
  INV_X1 npu_inst_pe_1_6_5_U11 ( .A(npu_inst_pe_1_6_5_n54), .ZN(
        npu_inst_pe_1_6_5_n117) );
  INV_X1 npu_inst_pe_1_6_5_U10 ( .A(npu_inst_pe_1_6_5_n50), .ZN(
        npu_inst_pe_1_6_5_n116) );
  INV_X1 npu_inst_pe_1_6_5_U9 ( .A(npu_inst_pe_1_6_5_n46), .ZN(
        npu_inst_pe_1_6_5_n115) );
  INV_X1 npu_inst_pe_1_6_5_U8 ( .A(npu_inst_pe_1_6_5_n42), .ZN(
        npu_inst_pe_1_6_5_n114) );
  BUF_X1 npu_inst_pe_1_6_5_U7 ( .A(npu_inst_pe_1_6_5_n11), .Z(
        npu_inst_pe_1_6_5_n10) );
  BUF_X1 npu_inst_pe_1_6_5_U6 ( .A(npu_inst_pe_1_6_5_n11), .Z(
        npu_inst_pe_1_6_5_n9) );
  BUF_X1 npu_inst_pe_1_6_5_U5 ( .A(npu_inst_pe_1_6_5_n11), .Z(
        npu_inst_pe_1_6_5_n8) );
  NOR2_X1 npu_inst_pe_1_6_5_U4 ( .A1(npu_inst_pe_1_6_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_5_n1), .ZN(npu_inst_pe_1_6_5_n76) );
  NOR2_X1 npu_inst_pe_1_6_5_U3 ( .A1(npu_inst_pe_1_6_5_n27), .A2(
        npu_inst_pe_1_6_5_n1), .ZN(npu_inst_pe_1_6_5_n77) );
  FA_X1 npu_inst_pe_1_6_5_sub_77_U2_1 ( .A(npu_inst_int_data_res_6__5__1_), 
        .B(npu_inst_pe_1_6_5_n13), .CI(npu_inst_pe_1_6_5_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_6_5_sub_77_carry_2_), .S(npu_inst_pe_1_6_5_N66) );
  FA_X1 npu_inst_pe_1_6_5_add_79_U1_1 ( .A(npu_inst_int_data_res_6__5__1_), 
        .B(npu_inst_pe_1_6_5_int_data_1_), .CI(
        npu_inst_pe_1_6_5_add_79_carry_1_), .CO(
        npu_inst_pe_1_6_5_add_79_carry_2_), .S(npu_inst_pe_1_6_5_N74) );
  NAND3_X1 npu_inst_pe_1_6_5_U101 ( .A1(npu_inst_pe_1_6_5_n4), .A2(
        npu_inst_pe_1_6_5_n6), .A3(npu_inst_pe_1_6_5_n7), .ZN(
        npu_inst_pe_1_6_5_n44) );
  NAND3_X1 npu_inst_pe_1_6_5_U100 ( .A1(npu_inst_pe_1_6_5_n3), .A2(
        npu_inst_pe_1_6_5_n6), .A3(npu_inst_pe_1_6_5_n7), .ZN(
        npu_inst_pe_1_6_5_n40) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_5_n33), .CK(
        npu_inst_pe_1_6_5_net3259), .RN(npu_inst_pe_1_6_5_n8), .Q(
        npu_inst_int_data_res_6__5__6_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_5_n34), .CK(
        npu_inst_pe_1_6_5_net3259), .RN(npu_inst_pe_1_6_5_n8), .Q(
        npu_inst_int_data_res_6__5__5_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_5_n35), .CK(
        npu_inst_pe_1_6_5_net3259), .RN(npu_inst_pe_1_6_5_n8), .Q(
        npu_inst_int_data_res_6__5__4_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_5_n36), .CK(
        npu_inst_pe_1_6_5_net3259), .RN(npu_inst_pe_1_6_5_n8), .Q(
        npu_inst_int_data_res_6__5__3_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_5_n98), .CK(
        npu_inst_pe_1_6_5_net3259), .RN(npu_inst_pe_1_6_5_n8), .Q(
        npu_inst_int_data_res_6__5__2_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_5_n99), .CK(
        npu_inst_pe_1_6_5_net3259), .RN(npu_inst_pe_1_6_5_n8), .Q(
        npu_inst_int_data_res_6__5__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_5_n32), .CK(
        npu_inst_pe_1_6_5_net3259), .RN(npu_inst_pe_1_6_5_n8), .Q(
        npu_inst_int_data_res_6__5__7_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_5_n100), 
        .CK(npu_inst_pe_1_6_5_net3259), .RN(npu_inst_pe_1_6_5_n8), .Q(
        npu_inst_int_data_res_6__5__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_weight_reg_0_ ( .D(npu_inst_n90), .CK(
        npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n8), .Q(
        npu_inst_pe_1_6_5_int_q_weight_0_), .QN(npu_inst_pe_1_6_5_n27) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_weight_reg_1_ ( .D(npu_inst_n96), .CK(
        npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n8), .Q(
        npu_inst_pe_1_6_5_int_q_weight_1_), .QN(npu_inst_pe_1_6_5_n26) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_5_n112), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n8), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_5_n106), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n8), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_5_n111), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_5_n105), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_5_n110), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_5_n104), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_5_n109), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_5_n103), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_5_n108), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_5_n102), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_5_n107), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_5_n101), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_5_n86), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_5_n87), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n9), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_5_n88), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_5_n89), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_5_n90), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_5_n91), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_5_n92), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_5_n93), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_5_n94), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_5_n95), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_5_n96), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_5_n97), 
        .CK(npu_inst_pe_1_6_5_net3265), .RN(npu_inst_pe_1_6_5_n10), .Q(
        npu_inst_pe_1_6_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_5_net3259) );
  CLKGATETST_X1 npu_inst_pe_1_6_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n43), .SE(1'b0), .GCK(npu_inst_pe_1_6_5_net3265) );
  MUX2_X1 npu_inst_pe_1_6_6_U153 ( .A(npu_inst_pe_1_6_6_n31), .B(
        npu_inst_pe_1_6_6_n28), .S(npu_inst_pe_1_6_6_n7), .Z(
        npu_inst_pe_1_6_6_N93) );
  MUX2_X1 npu_inst_pe_1_6_6_U152 ( .A(npu_inst_pe_1_6_6_n30), .B(
        npu_inst_pe_1_6_6_n29), .S(npu_inst_pe_1_6_6_n5), .Z(
        npu_inst_pe_1_6_6_n31) );
  MUX2_X1 npu_inst_pe_1_6_6_U151 ( .A(npu_inst_pe_1_6_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_6_n3), .Z(
        npu_inst_pe_1_6_6_n30) );
  MUX2_X1 npu_inst_pe_1_6_6_U150 ( .A(npu_inst_pe_1_6_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_6_n3), .Z(
        npu_inst_pe_1_6_6_n29) );
  MUX2_X1 npu_inst_pe_1_6_6_U149 ( .A(npu_inst_pe_1_6_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_6_n3), .Z(
        npu_inst_pe_1_6_6_n28) );
  MUX2_X1 npu_inst_pe_1_6_6_U148 ( .A(npu_inst_pe_1_6_6_n25), .B(
        npu_inst_pe_1_6_6_n22), .S(npu_inst_pe_1_6_6_n7), .Z(
        npu_inst_pe_1_6_6_N94) );
  MUX2_X1 npu_inst_pe_1_6_6_U147 ( .A(npu_inst_pe_1_6_6_n24), .B(
        npu_inst_pe_1_6_6_n23), .S(npu_inst_pe_1_6_6_n5), .Z(
        npu_inst_pe_1_6_6_n25) );
  MUX2_X1 npu_inst_pe_1_6_6_U146 ( .A(npu_inst_pe_1_6_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_6_n3), .Z(
        npu_inst_pe_1_6_6_n24) );
  MUX2_X1 npu_inst_pe_1_6_6_U145 ( .A(npu_inst_pe_1_6_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_6_n3), .Z(
        npu_inst_pe_1_6_6_n23) );
  MUX2_X1 npu_inst_pe_1_6_6_U144 ( .A(npu_inst_pe_1_6_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_6_n3), .Z(
        npu_inst_pe_1_6_6_n22) );
  MUX2_X1 npu_inst_pe_1_6_6_U143 ( .A(npu_inst_pe_1_6_6_n21), .B(
        npu_inst_pe_1_6_6_n18), .S(npu_inst_pe_1_6_6_n7), .Z(
        npu_inst_int_data_x_6__6__1_) );
  MUX2_X1 npu_inst_pe_1_6_6_U142 ( .A(npu_inst_pe_1_6_6_n20), .B(
        npu_inst_pe_1_6_6_n19), .S(npu_inst_pe_1_6_6_n5), .Z(
        npu_inst_pe_1_6_6_n21) );
  MUX2_X1 npu_inst_pe_1_6_6_U141 ( .A(npu_inst_pe_1_6_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_6_n3), .Z(
        npu_inst_pe_1_6_6_n20) );
  MUX2_X1 npu_inst_pe_1_6_6_U140 ( .A(npu_inst_pe_1_6_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_6_n3), .Z(
        npu_inst_pe_1_6_6_n19) );
  MUX2_X1 npu_inst_pe_1_6_6_U139 ( .A(npu_inst_pe_1_6_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_6_n3), .Z(
        npu_inst_pe_1_6_6_n18) );
  MUX2_X1 npu_inst_pe_1_6_6_U138 ( .A(npu_inst_pe_1_6_6_n17), .B(
        npu_inst_pe_1_6_6_n14), .S(npu_inst_pe_1_6_6_n7), .Z(
        npu_inst_int_data_x_6__6__0_) );
  MUX2_X1 npu_inst_pe_1_6_6_U137 ( .A(npu_inst_pe_1_6_6_n16), .B(
        npu_inst_pe_1_6_6_n15), .S(npu_inst_pe_1_6_6_n5), .Z(
        npu_inst_pe_1_6_6_n17) );
  MUX2_X1 npu_inst_pe_1_6_6_U136 ( .A(npu_inst_pe_1_6_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_6_n3), .Z(
        npu_inst_pe_1_6_6_n16) );
  MUX2_X1 npu_inst_pe_1_6_6_U135 ( .A(npu_inst_pe_1_6_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_6_n3), .Z(
        npu_inst_pe_1_6_6_n15) );
  MUX2_X1 npu_inst_pe_1_6_6_U134 ( .A(npu_inst_pe_1_6_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_6_n3), .Z(
        npu_inst_pe_1_6_6_n14) );
  XOR2_X1 npu_inst_pe_1_6_6_U133 ( .A(npu_inst_pe_1_6_6_int_data_0_), .B(
        npu_inst_int_data_res_6__6__0_), .Z(npu_inst_pe_1_6_6_N73) );
  AND2_X1 npu_inst_pe_1_6_6_U132 ( .A1(npu_inst_int_data_res_6__6__0_), .A2(
        npu_inst_pe_1_6_6_int_data_0_), .ZN(npu_inst_pe_1_6_6_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_6_U131 ( .A(npu_inst_int_data_res_6__6__0_), .B(
        npu_inst_pe_1_6_6_n12), .ZN(npu_inst_pe_1_6_6_N65) );
  OR2_X1 npu_inst_pe_1_6_6_U130 ( .A1(npu_inst_pe_1_6_6_n12), .A2(
        npu_inst_int_data_res_6__6__0_), .ZN(npu_inst_pe_1_6_6_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_6_U129 ( .A(npu_inst_int_data_res_6__6__2_), .B(
        npu_inst_pe_1_6_6_add_79_carry_2_), .Z(npu_inst_pe_1_6_6_N75) );
  AND2_X1 npu_inst_pe_1_6_6_U128 ( .A1(npu_inst_pe_1_6_6_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_6__6__2_), .ZN(
        npu_inst_pe_1_6_6_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_6_U127 ( .A(npu_inst_int_data_res_6__6__3_), .B(
        npu_inst_pe_1_6_6_add_79_carry_3_), .Z(npu_inst_pe_1_6_6_N76) );
  AND2_X1 npu_inst_pe_1_6_6_U126 ( .A1(npu_inst_pe_1_6_6_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_6__6__3_), .ZN(
        npu_inst_pe_1_6_6_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_6_U125 ( .A(npu_inst_int_data_res_6__6__4_), .B(
        npu_inst_pe_1_6_6_add_79_carry_4_), .Z(npu_inst_pe_1_6_6_N77) );
  AND2_X1 npu_inst_pe_1_6_6_U124 ( .A1(npu_inst_pe_1_6_6_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_6__6__4_), .ZN(
        npu_inst_pe_1_6_6_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_6_U123 ( .A(npu_inst_int_data_res_6__6__5_), .B(
        npu_inst_pe_1_6_6_add_79_carry_5_), .Z(npu_inst_pe_1_6_6_N78) );
  AND2_X1 npu_inst_pe_1_6_6_U122 ( .A1(npu_inst_pe_1_6_6_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_6__6__5_), .ZN(
        npu_inst_pe_1_6_6_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_6_U121 ( .A(npu_inst_int_data_res_6__6__6_), .B(
        npu_inst_pe_1_6_6_add_79_carry_6_), .Z(npu_inst_pe_1_6_6_N79) );
  AND2_X1 npu_inst_pe_1_6_6_U120 ( .A1(npu_inst_pe_1_6_6_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_6__6__6_), .ZN(
        npu_inst_pe_1_6_6_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_6_U119 ( .A(npu_inst_int_data_res_6__6__7_), .B(
        npu_inst_pe_1_6_6_add_79_carry_7_), .Z(npu_inst_pe_1_6_6_N80) );
  XNOR2_X1 npu_inst_pe_1_6_6_U118 ( .A(npu_inst_pe_1_6_6_sub_77_carry_2_), .B(
        npu_inst_int_data_res_6__6__2_), .ZN(npu_inst_pe_1_6_6_N67) );
  OR2_X1 npu_inst_pe_1_6_6_U117 ( .A1(npu_inst_int_data_res_6__6__2_), .A2(
        npu_inst_pe_1_6_6_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_6_6_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_6_U116 ( .A(npu_inst_pe_1_6_6_sub_77_carry_3_), .B(
        npu_inst_int_data_res_6__6__3_), .ZN(npu_inst_pe_1_6_6_N68) );
  OR2_X1 npu_inst_pe_1_6_6_U115 ( .A1(npu_inst_int_data_res_6__6__3_), .A2(
        npu_inst_pe_1_6_6_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_6_6_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_6_U114 ( .A(npu_inst_pe_1_6_6_sub_77_carry_4_), .B(
        npu_inst_int_data_res_6__6__4_), .ZN(npu_inst_pe_1_6_6_N69) );
  OR2_X1 npu_inst_pe_1_6_6_U113 ( .A1(npu_inst_int_data_res_6__6__4_), .A2(
        npu_inst_pe_1_6_6_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_6_6_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_6_U112 ( .A(npu_inst_pe_1_6_6_sub_77_carry_5_), .B(
        npu_inst_int_data_res_6__6__5_), .ZN(npu_inst_pe_1_6_6_N70) );
  OR2_X1 npu_inst_pe_1_6_6_U111 ( .A1(npu_inst_int_data_res_6__6__5_), .A2(
        npu_inst_pe_1_6_6_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_6_6_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_6_U110 ( .A(npu_inst_pe_1_6_6_sub_77_carry_6_), .B(
        npu_inst_int_data_res_6__6__6_), .ZN(npu_inst_pe_1_6_6_N71) );
  OR2_X1 npu_inst_pe_1_6_6_U109 ( .A1(npu_inst_int_data_res_6__6__6_), .A2(
        npu_inst_pe_1_6_6_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_6_6_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_6_U108 ( .A(npu_inst_int_data_res_6__6__7_), .B(
        npu_inst_pe_1_6_6_sub_77_carry_7_), .ZN(npu_inst_pe_1_6_6_N72) );
  INV_X1 npu_inst_pe_1_6_6_U107 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_6_6_n6)
         );
  INV_X1 npu_inst_pe_1_6_6_U106 ( .A(npu_inst_pe_1_6_6_n6), .ZN(
        npu_inst_pe_1_6_6_n5) );
  INV_X1 npu_inst_pe_1_6_6_U105 ( .A(npu_inst_n35), .ZN(npu_inst_pe_1_6_6_n2)
         );
  AOI22_X1 npu_inst_pe_1_6_6_U104 ( .A1(npu_inst_int_data_y_7__6__0_), .A2(
        npu_inst_pe_1_6_6_n58), .B1(npu_inst_pe_1_6_6_n118), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_6_n57) );
  INV_X1 npu_inst_pe_1_6_6_U103 ( .A(npu_inst_pe_1_6_6_n57), .ZN(
        npu_inst_pe_1_6_6_n107) );
  AOI22_X1 npu_inst_pe_1_6_6_U102 ( .A1(npu_inst_int_data_y_7__6__0_), .A2(
        npu_inst_pe_1_6_6_n54), .B1(npu_inst_pe_1_6_6_n117), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_6_n53) );
  INV_X1 npu_inst_pe_1_6_6_U99 ( .A(npu_inst_pe_1_6_6_n53), .ZN(
        npu_inst_pe_1_6_6_n108) );
  AOI22_X1 npu_inst_pe_1_6_6_U98 ( .A1(npu_inst_int_data_y_7__6__0_), .A2(
        npu_inst_pe_1_6_6_n50), .B1(npu_inst_pe_1_6_6_n116), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_6_n49) );
  INV_X1 npu_inst_pe_1_6_6_U97 ( .A(npu_inst_pe_1_6_6_n49), .ZN(
        npu_inst_pe_1_6_6_n109) );
  AOI22_X1 npu_inst_pe_1_6_6_U96 ( .A1(npu_inst_int_data_y_7__6__0_), .A2(
        npu_inst_pe_1_6_6_n46), .B1(npu_inst_pe_1_6_6_n115), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_6_n45) );
  INV_X1 npu_inst_pe_1_6_6_U95 ( .A(npu_inst_pe_1_6_6_n45), .ZN(
        npu_inst_pe_1_6_6_n110) );
  AOI22_X1 npu_inst_pe_1_6_6_U94 ( .A1(npu_inst_int_data_y_7__6__0_), .A2(
        npu_inst_pe_1_6_6_n42), .B1(npu_inst_pe_1_6_6_n114), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_6_n41) );
  INV_X1 npu_inst_pe_1_6_6_U93 ( .A(npu_inst_pe_1_6_6_n41), .ZN(
        npu_inst_pe_1_6_6_n111) );
  AOI22_X1 npu_inst_pe_1_6_6_U92 ( .A1(npu_inst_int_data_y_7__6__1_), .A2(
        npu_inst_pe_1_6_6_n58), .B1(npu_inst_pe_1_6_6_n118), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_6_n59) );
  INV_X1 npu_inst_pe_1_6_6_U91 ( .A(npu_inst_pe_1_6_6_n59), .ZN(
        npu_inst_pe_1_6_6_n101) );
  AOI22_X1 npu_inst_pe_1_6_6_U90 ( .A1(npu_inst_int_data_y_7__6__1_), .A2(
        npu_inst_pe_1_6_6_n54), .B1(npu_inst_pe_1_6_6_n117), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_6_n55) );
  INV_X1 npu_inst_pe_1_6_6_U89 ( .A(npu_inst_pe_1_6_6_n55), .ZN(
        npu_inst_pe_1_6_6_n102) );
  AOI22_X1 npu_inst_pe_1_6_6_U88 ( .A1(npu_inst_int_data_y_7__6__1_), .A2(
        npu_inst_pe_1_6_6_n50), .B1(npu_inst_pe_1_6_6_n116), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_6_n51) );
  INV_X1 npu_inst_pe_1_6_6_U87 ( .A(npu_inst_pe_1_6_6_n51), .ZN(
        npu_inst_pe_1_6_6_n103) );
  AOI22_X1 npu_inst_pe_1_6_6_U86 ( .A1(npu_inst_int_data_y_7__6__1_), .A2(
        npu_inst_pe_1_6_6_n46), .B1(npu_inst_pe_1_6_6_n115), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_6_n47) );
  INV_X1 npu_inst_pe_1_6_6_U85 ( .A(npu_inst_pe_1_6_6_n47), .ZN(
        npu_inst_pe_1_6_6_n104) );
  AOI22_X1 npu_inst_pe_1_6_6_U84 ( .A1(npu_inst_int_data_y_7__6__1_), .A2(
        npu_inst_pe_1_6_6_n42), .B1(npu_inst_pe_1_6_6_n114), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_6_n43) );
  INV_X1 npu_inst_pe_1_6_6_U83 ( .A(npu_inst_pe_1_6_6_n43), .ZN(
        npu_inst_pe_1_6_6_n105) );
  AOI22_X1 npu_inst_pe_1_6_6_U82 ( .A1(npu_inst_pe_1_6_6_n38), .A2(
        npu_inst_int_data_y_7__6__1_), .B1(npu_inst_pe_1_6_6_n113), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_6_n39) );
  INV_X1 npu_inst_pe_1_6_6_U81 ( .A(npu_inst_pe_1_6_6_n39), .ZN(
        npu_inst_pe_1_6_6_n106) );
  AND2_X1 npu_inst_pe_1_6_6_U80 ( .A1(npu_inst_pe_1_6_6_N93), .A2(npu_inst_n35), .ZN(npu_inst_int_data_y_6__6__0_) );
  NAND2_X1 npu_inst_pe_1_6_6_U79 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_6_n60), .ZN(npu_inst_pe_1_6_6_n74) );
  OAI21_X1 npu_inst_pe_1_6_6_U78 ( .B1(npu_inst_pe_1_6_6_n63), .B2(
        npu_inst_pe_1_6_6_n60), .A(npu_inst_pe_1_6_6_n74), .ZN(
        npu_inst_pe_1_6_6_n97) );
  NAND2_X1 npu_inst_pe_1_6_6_U77 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_6_n60), .ZN(npu_inst_pe_1_6_6_n73) );
  OAI21_X1 npu_inst_pe_1_6_6_U76 ( .B1(npu_inst_pe_1_6_6_n61), .B2(
        npu_inst_pe_1_6_6_n60), .A(npu_inst_pe_1_6_6_n73), .ZN(
        npu_inst_pe_1_6_6_n96) );
  NAND2_X1 npu_inst_pe_1_6_6_U75 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_6_n56), .ZN(npu_inst_pe_1_6_6_n72) );
  OAI21_X1 npu_inst_pe_1_6_6_U74 ( .B1(npu_inst_pe_1_6_6_n63), .B2(
        npu_inst_pe_1_6_6_n56), .A(npu_inst_pe_1_6_6_n72), .ZN(
        npu_inst_pe_1_6_6_n95) );
  NAND2_X1 npu_inst_pe_1_6_6_U73 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_6_n56), .ZN(npu_inst_pe_1_6_6_n71) );
  OAI21_X1 npu_inst_pe_1_6_6_U72 ( .B1(npu_inst_pe_1_6_6_n61), .B2(
        npu_inst_pe_1_6_6_n56), .A(npu_inst_pe_1_6_6_n71), .ZN(
        npu_inst_pe_1_6_6_n94) );
  NAND2_X1 npu_inst_pe_1_6_6_U71 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_6_n52), .ZN(npu_inst_pe_1_6_6_n70) );
  OAI21_X1 npu_inst_pe_1_6_6_U70 ( .B1(npu_inst_pe_1_6_6_n63), .B2(
        npu_inst_pe_1_6_6_n52), .A(npu_inst_pe_1_6_6_n70), .ZN(
        npu_inst_pe_1_6_6_n93) );
  NAND2_X1 npu_inst_pe_1_6_6_U69 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_6_n52), .ZN(npu_inst_pe_1_6_6_n69) );
  OAI21_X1 npu_inst_pe_1_6_6_U68 ( .B1(npu_inst_pe_1_6_6_n61), .B2(
        npu_inst_pe_1_6_6_n52), .A(npu_inst_pe_1_6_6_n69), .ZN(
        npu_inst_pe_1_6_6_n92) );
  NAND2_X1 npu_inst_pe_1_6_6_U67 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_6_n48), .ZN(npu_inst_pe_1_6_6_n68) );
  OAI21_X1 npu_inst_pe_1_6_6_U66 ( .B1(npu_inst_pe_1_6_6_n63), .B2(
        npu_inst_pe_1_6_6_n48), .A(npu_inst_pe_1_6_6_n68), .ZN(
        npu_inst_pe_1_6_6_n91) );
  NAND2_X1 npu_inst_pe_1_6_6_U65 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_6_n48), .ZN(npu_inst_pe_1_6_6_n67) );
  OAI21_X1 npu_inst_pe_1_6_6_U64 ( .B1(npu_inst_pe_1_6_6_n61), .B2(
        npu_inst_pe_1_6_6_n48), .A(npu_inst_pe_1_6_6_n67), .ZN(
        npu_inst_pe_1_6_6_n90) );
  NAND2_X1 npu_inst_pe_1_6_6_U63 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_6_n44), .ZN(npu_inst_pe_1_6_6_n66) );
  OAI21_X1 npu_inst_pe_1_6_6_U62 ( .B1(npu_inst_pe_1_6_6_n63), .B2(
        npu_inst_pe_1_6_6_n44), .A(npu_inst_pe_1_6_6_n66), .ZN(
        npu_inst_pe_1_6_6_n89) );
  NAND2_X1 npu_inst_pe_1_6_6_U61 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_6_n44), .ZN(npu_inst_pe_1_6_6_n65) );
  OAI21_X1 npu_inst_pe_1_6_6_U60 ( .B1(npu_inst_pe_1_6_6_n61), .B2(
        npu_inst_pe_1_6_6_n44), .A(npu_inst_pe_1_6_6_n65), .ZN(
        npu_inst_pe_1_6_6_n88) );
  NAND2_X1 npu_inst_pe_1_6_6_U59 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_6_n40), .ZN(npu_inst_pe_1_6_6_n64) );
  OAI21_X1 npu_inst_pe_1_6_6_U58 ( .B1(npu_inst_pe_1_6_6_n63), .B2(
        npu_inst_pe_1_6_6_n40), .A(npu_inst_pe_1_6_6_n64), .ZN(
        npu_inst_pe_1_6_6_n87) );
  NAND2_X1 npu_inst_pe_1_6_6_U57 ( .A1(npu_inst_pe_1_6_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_6_n40), .ZN(npu_inst_pe_1_6_6_n62) );
  OAI21_X1 npu_inst_pe_1_6_6_U56 ( .B1(npu_inst_pe_1_6_6_n61), .B2(
        npu_inst_pe_1_6_6_n40), .A(npu_inst_pe_1_6_6_n62), .ZN(
        npu_inst_pe_1_6_6_n86) );
  AOI22_X1 npu_inst_pe_1_6_6_U55 ( .A1(npu_inst_pe_1_6_6_n38), .A2(
        npu_inst_int_data_y_7__6__0_), .B1(npu_inst_pe_1_6_6_n113), .B2(
        npu_inst_pe_1_6_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_6_n37) );
  INV_X1 npu_inst_pe_1_6_6_U54 ( .A(npu_inst_pe_1_6_6_n37), .ZN(
        npu_inst_pe_1_6_6_n112) );
  AND2_X1 npu_inst_pe_1_6_6_U53 ( .A1(npu_inst_n35), .A2(npu_inst_pe_1_6_6_N94), .ZN(npu_inst_int_data_y_6__6__1_) );
  AOI222_X1 npu_inst_pe_1_6_6_U52 ( .A1(npu_inst_int_data_res_7__6__0_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N73), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N65), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n84) );
  INV_X1 npu_inst_pe_1_6_6_U51 ( .A(npu_inst_pe_1_6_6_n84), .ZN(
        npu_inst_pe_1_6_6_n100) );
  AOI222_X1 npu_inst_pe_1_6_6_U50 ( .A1(npu_inst_pe_1_6_6_n1), .A2(
        npu_inst_int_data_res_7__6__7_), .B1(npu_inst_pe_1_6_6_N80), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N72), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n75) );
  INV_X1 npu_inst_pe_1_6_6_U49 ( .A(npu_inst_pe_1_6_6_n75), .ZN(
        npu_inst_pe_1_6_6_n32) );
  AOI222_X1 npu_inst_pe_1_6_6_U48 ( .A1(npu_inst_int_data_res_7__6__1_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N74), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N66), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n83) );
  INV_X1 npu_inst_pe_1_6_6_U47 ( .A(npu_inst_pe_1_6_6_n83), .ZN(
        npu_inst_pe_1_6_6_n99) );
  AOI222_X1 npu_inst_pe_1_6_6_U46 ( .A1(npu_inst_int_data_res_7__6__3_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N76), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N68), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n81) );
  INV_X1 npu_inst_pe_1_6_6_U45 ( .A(npu_inst_pe_1_6_6_n81), .ZN(
        npu_inst_pe_1_6_6_n36) );
  AOI222_X1 npu_inst_pe_1_6_6_U44 ( .A1(npu_inst_int_data_res_7__6__4_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N77), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N69), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n80) );
  INV_X1 npu_inst_pe_1_6_6_U43 ( .A(npu_inst_pe_1_6_6_n80), .ZN(
        npu_inst_pe_1_6_6_n35) );
  AOI222_X1 npu_inst_pe_1_6_6_U42 ( .A1(npu_inst_int_data_res_7__6__5_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N78), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N70), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n79) );
  INV_X1 npu_inst_pe_1_6_6_U41 ( .A(npu_inst_pe_1_6_6_n79), .ZN(
        npu_inst_pe_1_6_6_n34) );
  AOI222_X1 npu_inst_pe_1_6_6_U40 ( .A1(npu_inst_int_data_res_7__6__6_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N79), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N71), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n78) );
  INV_X1 npu_inst_pe_1_6_6_U39 ( .A(npu_inst_pe_1_6_6_n78), .ZN(
        npu_inst_pe_1_6_6_n33) );
  AND2_X1 npu_inst_pe_1_6_6_U38 ( .A1(npu_inst_int_data_x_6__6__1_), .A2(
        npu_inst_pe_1_6_6_int_q_weight_1_), .ZN(npu_inst_pe_1_6_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_6_U37 ( .A1(npu_inst_int_data_x_6__6__0_), .A2(
        npu_inst_pe_1_6_6_int_q_weight_1_), .ZN(npu_inst_pe_1_6_6_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_6_6_U36 ( .A(npu_inst_pe_1_6_6_int_data_1_), .ZN(
        npu_inst_pe_1_6_6_n13) );
  NOR3_X1 npu_inst_pe_1_6_6_U35 ( .A1(npu_inst_pe_1_6_6_n26), .A2(npu_inst_n35), .A3(npu_inst_int_ckg[9]), .ZN(npu_inst_pe_1_6_6_n85) );
  OR2_X1 npu_inst_pe_1_6_6_U34 ( .A1(npu_inst_pe_1_6_6_n85), .A2(
        npu_inst_pe_1_6_6_n1), .ZN(npu_inst_pe_1_6_6_N84) );
  AOI222_X1 npu_inst_pe_1_6_6_U33 ( .A1(npu_inst_int_data_res_7__6__2_), .A2(
        npu_inst_pe_1_6_6_n1), .B1(npu_inst_pe_1_6_6_N75), .B2(
        npu_inst_pe_1_6_6_n76), .C1(npu_inst_pe_1_6_6_N67), .C2(
        npu_inst_pe_1_6_6_n77), .ZN(npu_inst_pe_1_6_6_n82) );
  INV_X1 npu_inst_pe_1_6_6_U32 ( .A(npu_inst_pe_1_6_6_n82), .ZN(
        npu_inst_pe_1_6_6_n98) );
  AOI22_X1 npu_inst_pe_1_6_6_U31 ( .A1(npu_inst_n35), .A2(
        npu_inst_int_data_y_7__6__1_), .B1(npu_inst_pe_1_6_6_n2), .B2(
        npu_inst_int_data_x_6__7__1_), .ZN(npu_inst_pe_1_6_6_n63) );
  AOI22_X1 npu_inst_pe_1_6_6_U30 ( .A1(npu_inst_n35), .A2(
        npu_inst_int_data_y_7__6__0_), .B1(npu_inst_pe_1_6_6_n2), .B2(
        npu_inst_int_data_x_6__7__0_), .ZN(npu_inst_pe_1_6_6_n61) );
  INV_X1 npu_inst_pe_1_6_6_U29 ( .A(npu_inst_pe_1_6_6_int_data_0_), .ZN(
        npu_inst_pe_1_6_6_n12) );
  INV_X1 npu_inst_pe_1_6_6_U28 ( .A(npu_inst_n49), .ZN(npu_inst_pe_1_6_6_n4)
         );
  OR3_X1 npu_inst_pe_1_6_6_U27 ( .A1(npu_inst_pe_1_6_6_n5), .A2(
        npu_inst_pe_1_6_6_n7), .A3(npu_inst_pe_1_6_6_n4), .ZN(
        npu_inst_pe_1_6_6_n56) );
  OR3_X1 npu_inst_pe_1_6_6_U26 ( .A1(npu_inst_pe_1_6_6_n4), .A2(
        npu_inst_pe_1_6_6_n7), .A3(npu_inst_pe_1_6_6_n6), .ZN(
        npu_inst_pe_1_6_6_n48) );
  INV_X1 npu_inst_pe_1_6_6_U25 ( .A(npu_inst_pe_1_6_6_n4), .ZN(
        npu_inst_pe_1_6_6_n3) );
  OR3_X1 npu_inst_pe_1_6_6_U24 ( .A1(npu_inst_pe_1_6_6_n3), .A2(
        npu_inst_pe_1_6_6_n7), .A3(npu_inst_pe_1_6_6_n6), .ZN(
        npu_inst_pe_1_6_6_n52) );
  OR3_X1 npu_inst_pe_1_6_6_U23 ( .A1(npu_inst_pe_1_6_6_n5), .A2(
        npu_inst_pe_1_6_6_n7), .A3(npu_inst_pe_1_6_6_n3), .ZN(
        npu_inst_pe_1_6_6_n60) );
  BUF_X1 npu_inst_pe_1_6_6_U22 ( .A(npu_inst_n14), .Z(npu_inst_pe_1_6_6_n1) );
  NOR2_X1 npu_inst_pe_1_6_6_U21 ( .A1(npu_inst_pe_1_6_6_n60), .A2(
        npu_inst_pe_1_6_6_n2), .ZN(npu_inst_pe_1_6_6_n58) );
  NOR2_X1 npu_inst_pe_1_6_6_U20 ( .A1(npu_inst_pe_1_6_6_n56), .A2(
        npu_inst_pe_1_6_6_n2), .ZN(npu_inst_pe_1_6_6_n54) );
  NOR2_X1 npu_inst_pe_1_6_6_U19 ( .A1(npu_inst_pe_1_6_6_n52), .A2(
        npu_inst_pe_1_6_6_n2), .ZN(npu_inst_pe_1_6_6_n50) );
  NOR2_X1 npu_inst_pe_1_6_6_U18 ( .A1(npu_inst_pe_1_6_6_n48), .A2(
        npu_inst_pe_1_6_6_n2), .ZN(npu_inst_pe_1_6_6_n46) );
  NOR2_X1 npu_inst_pe_1_6_6_U17 ( .A1(npu_inst_pe_1_6_6_n40), .A2(
        npu_inst_pe_1_6_6_n2), .ZN(npu_inst_pe_1_6_6_n38) );
  NOR2_X1 npu_inst_pe_1_6_6_U16 ( .A1(npu_inst_pe_1_6_6_n44), .A2(
        npu_inst_pe_1_6_6_n2), .ZN(npu_inst_pe_1_6_6_n42) );
  BUF_X1 npu_inst_pe_1_6_6_U15 ( .A(npu_inst_n76), .Z(npu_inst_pe_1_6_6_n7) );
  INV_X1 npu_inst_pe_1_6_6_U14 ( .A(npu_inst_n104), .ZN(npu_inst_pe_1_6_6_n11)
         );
  INV_X1 npu_inst_pe_1_6_6_U13 ( .A(npu_inst_pe_1_6_6_n38), .ZN(
        npu_inst_pe_1_6_6_n113) );
  INV_X1 npu_inst_pe_1_6_6_U12 ( .A(npu_inst_pe_1_6_6_n58), .ZN(
        npu_inst_pe_1_6_6_n118) );
  INV_X1 npu_inst_pe_1_6_6_U11 ( .A(npu_inst_pe_1_6_6_n54), .ZN(
        npu_inst_pe_1_6_6_n117) );
  INV_X1 npu_inst_pe_1_6_6_U10 ( .A(npu_inst_pe_1_6_6_n50), .ZN(
        npu_inst_pe_1_6_6_n116) );
  INV_X1 npu_inst_pe_1_6_6_U9 ( .A(npu_inst_pe_1_6_6_n46), .ZN(
        npu_inst_pe_1_6_6_n115) );
  INV_X1 npu_inst_pe_1_6_6_U8 ( .A(npu_inst_pe_1_6_6_n42), .ZN(
        npu_inst_pe_1_6_6_n114) );
  BUF_X1 npu_inst_pe_1_6_6_U7 ( .A(npu_inst_pe_1_6_6_n11), .Z(
        npu_inst_pe_1_6_6_n10) );
  BUF_X1 npu_inst_pe_1_6_6_U6 ( .A(npu_inst_pe_1_6_6_n11), .Z(
        npu_inst_pe_1_6_6_n9) );
  BUF_X1 npu_inst_pe_1_6_6_U5 ( .A(npu_inst_pe_1_6_6_n11), .Z(
        npu_inst_pe_1_6_6_n8) );
  NOR2_X1 npu_inst_pe_1_6_6_U4 ( .A1(npu_inst_pe_1_6_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_6_n1), .ZN(npu_inst_pe_1_6_6_n76) );
  NOR2_X1 npu_inst_pe_1_6_6_U3 ( .A1(npu_inst_pe_1_6_6_n27), .A2(
        npu_inst_pe_1_6_6_n1), .ZN(npu_inst_pe_1_6_6_n77) );
  FA_X1 npu_inst_pe_1_6_6_sub_77_U2_1 ( .A(npu_inst_int_data_res_6__6__1_), 
        .B(npu_inst_pe_1_6_6_n13), .CI(npu_inst_pe_1_6_6_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_6_6_sub_77_carry_2_), .S(npu_inst_pe_1_6_6_N66) );
  FA_X1 npu_inst_pe_1_6_6_add_79_U1_1 ( .A(npu_inst_int_data_res_6__6__1_), 
        .B(npu_inst_pe_1_6_6_int_data_1_), .CI(
        npu_inst_pe_1_6_6_add_79_carry_1_), .CO(
        npu_inst_pe_1_6_6_add_79_carry_2_), .S(npu_inst_pe_1_6_6_N74) );
  NAND3_X1 npu_inst_pe_1_6_6_U101 ( .A1(npu_inst_pe_1_6_6_n4), .A2(
        npu_inst_pe_1_6_6_n6), .A3(npu_inst_pe_1_6_6_n7), .ZN(
        npu_inst_pe_1_6_6_n44) );
  NAND3_X1 npu_inst_pe_1_6_6_U100 ( .A1(npu_inst_pe_1_6_6_n3), .A2(
        npu_inst_pe_1_6_6_n6), .A3(npu_inst_pe_1_6_6_n7), .ZN(
        npu_inst_pe_1_6_6_n40) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_6_n33), .CK(
        npu_inst_pe_1_6_6_net3236), .RN(npu_inst_pe_1_6_6_n8), .Q(
        npu_inst_int_data_res_6__6__6_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_6_n34), .CK(
        npu_inst_pe_1_6_6_net3236), .RN(npu_inst_pe_1_6_6_n8), .Q(
        npu_inst_int_data_res_6__6__5_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_6_n35), .CK(
        npu_inst_pe_1_6_6_net3236), .RN(npu_inst_pe_1_6_6_n8), .Q(
        npu_inst_int_data_res_6__6__4_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_6_n36), .CK(
        npu_inst_pe_1_6_6_net3236), .RN(npu_inst_pe_1_6_6_n8), .Q(
        npu_inst_int_data_res_6__6__3_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_6_n98), .CK(
        npu_inst_pe_1_6_6_net3236), .RN(npu_inst_pe_1_6_6_n8), .Q(
        npu_inst_int_data_res_6__6__2_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_6_n99), .CK(
        npu_inst_pe_1_6_6_net3236), .RN(npu_inst_pe_1_6_6_n8), .Q(
        npu_inst_int_data_res_6__6__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_6_n32), .CK(
        npu_inst_pe_1_6_6_net3236), .RN(npu_inst_pe_1_6_6_n8), .Q(
        npu_inst_int_data_res_6__6__7_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_6_n100), 
        .CK(npu_inst_pe_1_6_6_net3236), .RN(npu_inst_pe_1_6_6_n8), .Q(
        npu_inst_int_data_res_6__6__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_weight_reg_0_ ( .D(npu_inst_n90), .CK(
        npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n8), .Q(
        npu_inst_pe_1_6_6_int_q_weight_0_), .QN(npu_inst_pe_1_6_6_n27) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_weight_reg_1_ ( .D(npu_inst_n96), .CK(
        npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n8), .Q(
        npu_inst_pe_1_6_6_int_q_weight_1_), .QN(npu_inst_pe_1_6_6_n26) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_6_n112), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n8), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_6_n106), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n8), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_6_n111), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_6_n105), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_6_n110), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_6_n104), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_6_n109), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_6_n103), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_6_n108), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_6_n102), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_6_n107), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_6_n101), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_6_n86), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_6_n87), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n9), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_6_n88), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_6_n89), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_6_n90), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_6_n91), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_6_n92), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_6_n93), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_6_n94), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_6_n95), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_6_n96), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_6_n97), 
        .CK(npu_inst_pe_1_6_6_net3242), .RN(npu_inst_pe_1_6_6_n10), .Q(
        npu_inst_pe_1_6_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_6_net3236) );
  CLKGATETST_X1 npu_inst_pe_1_6_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n43), .SE(1'b0), .GCK(npu_inst_pe_1_6_6_net3242) );
  MUX2_X1 npu_inst_pe_1_6_7_U153 ( .A(npu_inst_pe_1_6_7_n31), .B(
        npu_inst_pe_1_6_7_n28), .S(npu_inst_pe_1_6_7_n7), .Z(
        npu_inst_pe_1_6_7_N93) );
  MUX2_X1 npu_inst_pe_1_6_7_U152 ( .A(npu_inst_pe_1_6_7_n30), .B(
        npu_inst_pe_1_6_7_n29), .S(npu_inst_pe_1_6_7_n5), .Z(
        npu_inst_pe_1_6_7_n31) );
  MUX2_X1 npu_inst_pe_1_6_7_U151 ( .A(npu_inst_pe_1_6_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_6_7_n3), .Z(
        npu_inst_pe_1_6_7_n30) );
  MUX2_X1 npu_inst_pe_1_6_7_U150 ( .A(npu_inst_pe_1_6_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_6_7_n3), .Z(
        npu_inst_pe_1_6_7_n29) );
  MUX2_X1 npu_inst_pe_1_6_7_U149 ( .A(npu_inst_pe_1_6_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_6_7_n3), .Z(
        npu_inst_pe_1_6_7_n28) );
  MUX2_X1 npu_inst_pe_1_6_7_U148 ( .A(npu_inst_pe_1_6_7_n25), .B(
        npu_inst_pe_1_6_7_n22), .S(npu_inst_pe_1_6_7_n7), .Z(
        npu_inst_pe_1_6_7_N94) );
  MUX2_X1 npu_inst_pe_1_6_7_U147 ( .A(npu_inst_pe_1_6_7_n24), .B(
        npu_inst_pe_1_6_7_n23), .S(npu_inst_pe_1_6_7_n5), .Z(
        npu_inst_pe_1_6_7_n25) );
  MUX2_X1 npu_inst_pe_1_6_7_U146 ( .A(npu_inst_pe_1_6_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_6_7_n3), .Z(
        npu_inst_pe_1_6_7_n24) );
  MUX2_X1 npu_inst_pe_1_6_7_U145 ( .A(npu_inst_pe_1_6_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_6_7_n3), .Z(
        npu_inst_pe_1_6_7_n23) );
  MUX2_X1 npu_inst_pe_1_6_7_U144 ( .A(npu_inst_pe_1_6_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_6_7_n3), .Z(
        npu_inst_pe_1_6_7_n22) );
  MUX2_X1 npu_inst_pe_1_6_7_U143 ( .A(npu_inst_pe_1_6_7_n21), .B(
        npu_inst_pe_1_6_7_n18), .S(npu_inst_pe_1_6_7_n7), .Z(
        npu_inst_int_data_x_6__7__1_) );
  MUX2_X1 npu_inst_pe_1_6_7_U142 ( .A(npu_inst_pe_1_6_7_n20), .B(
        npu_inst_pe_1_6_7_n19), .S(npu_inst_pe_1_6_7_n5), .Z(
        npu_inst_pe_1_6_7_n21) );
  MUX2_X1 npu_inst_pe_1_6_7_U141 ( .A(npu_inst_pe_1_6_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_6_7_n3), .Z(
        npu_inst_pe_1_6_7_n20) );
  MUX2_X1 npu_inst_pe_1_6_7_U140 ( .A(npu_inst_pe_1_6_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_6_7_n3), .Z(
        npu_inst_pe_1_6_7_n19) );
  MUX2_X1 npu_inst_pe_1_6_7_U139 ( .A(npu_inst_pe_1_6_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_6_7_n3), .Z(
        npu_inst_pe_1_6_7_n18) );
  MUX2_X1 npu_inst_pe_1_6_7_U138 ( .A(npu_inst_pe_1_6_7_n17), .B(
        npu_inst_pe_1_6_7_n14), .S(npu_inst_pe_1_6_7_n7), .Z(
        npu_inst_int_data_x_6__7__0_) );
  MUX2_X1 npu_inst_pe_1_6_7_U137 ( .A(npu_inst_pe_1_6_7_n16), .B(
        npu_inst_pe_1_6_7_n15), .S(npu_inst_pe_1_6_7_n5), .Z(
        npu_inst_pe_1_6_7_n17) );
  MUX2_X1 npu_inst_pe_1_6_7_U136 ( .A(npu_inst_pe_1_6_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_6_7_n3), .Z(
        npu_inst_pe_1_6_7_n16) );
  MUX2_X1 npu_inst_pe_1_6_7_U135 ( .A(npu_inst_pe_1_6_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_6_7_n3), .Z(
        npu_inst_pe_1_6_7_n15) );
  MUX2_X1 npu_inst_pe_1_6_7_U134 ( .A(npu_inst_pe_1_6_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_6_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_6_7_n3), .Z(
        npu_inst_pe_1_6_7_n14) );
  XOR2_X1 npu_inst_pe_1_6_7_U133 ( .A(npu_inst_pe_1_6_7_int_data_0_), .B(
        npu_inst_int_data_res_6__7__0_), .Z(npu_inst_pe_1_6_7_N73) );
  AND2_X1 npu_inst_pe_1_6_7_U132 ( .A1(npu_inst_int_data_res_6__7__0_), .A2(
        npu_inst_pe_1_6_7_int_data_0_), .ZN(npu_inst_pe_1_6_7_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_6_7_U131 ( .A(npu_inst_int_data_res_6__7__0_), .B(
        npu_inst_pe_1_6_7_n12), .ZN(npu_inst_pe_1_6_7_N65) );
  OR2_X1 npu_inst_pe_1_6_7_U130 ( .A1(npu_inst_pe_1_6_7_n12), .A2(
        npu_inst_int_data_res_6__7__0_), .ZN(npu_inst_pe_1_6_7_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_6_7_U129 ( .A(npu_inst_int_data_res_6__7__2_), .B(
        npu_inst_pe_1_6_7_add_79_carry_2_), .Z(npu_inst_pe_1_6_7_N75) );
  AND2_X1 npu_inst_pe_1_6_7_U128 ( .A1(npu_inst_pe_1_6_7_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_6__7__2_), .ZN(
        npu_inst_pe_1_6_7_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_6_7_U127 ( .A(npu_inst_int_data_res_6__7__3_), .B(
        npu_inst_pe_1_6_7_add_79_carry_3_), .Z(npu_inst_pe_1_6_7_N76) );
  AND2_X1 npu_inst_pe_1_6_7_U126 ( .A1(npu_inst_pe_1_6_7_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_6__7__3_), .ZN(
        npu_inst_pe_1_6_7_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_6_7_U125 ( .A(npu_inst_int_data_res_6__7__4_), .B(
        npu_inst_pe_1_6_7_add_79_carry_4_), .Z(npu_inst_pe_1_6_7_N77) );
  AND2_X1 npu_inst_pe_1_6_7_U124 ( .A1(npu_inst_pe_1_6_7_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_6__7__4_), .ZN(
        npu_inst_pe_1_6_7_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_6_7_U123 ( .A(npu_inst_int_data_res_6__7__5_), .B(
        npu_inst_pe_1_6_7_add_79_carry_5_), .Z(npu_inst_pe_1_6_7_N78) );
  AND2_X1 npu_inst_pe_1_6_7_U122 ( .A1(npu_inst_pe_1_6_7_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_6__7__5_), .ZN(
        npu_inst_pe_1_6_7_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_6_7_U121 ( .A(npu_inst_int_data_res_6__7__6_), .B(
        npu_inst_pe_1_6_7_add_79_carry_6_), .Z(npu_inst_pe_1_6_7_N79) );
  AND2_X1 npu_inst_pe_1_6_7_U120 ( .A1(npu_inst_pe_1_6_7_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_6__7__6_), .ZN(
        npu_inst_pe_1_6_7_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_6_7_U119 ( .A(npu_inst_int_data_res_6__7__7_), .B(
        npu_inst_pe_1_6_7_add_79_carry_7_), .Z(npu_inst_pe_1_6_7_N80) );
  XNOR2_X1 npu_inst_pe_1_6_7_U118 ( .A(npu_inst_pe_1_6_7_sub_77_carry_2_), .B(
        npu_inst_int_data_res_6__7__2_), .ZN(npu_inst_pe_1_6_7_N67) );
  OR2_X1 npu_inst_pe_1_6_7_U117 ( .A1(npu_inst_int_data_res_6__7__2_), .A2(
        npu_inst_pe_1_6_7_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_6_7_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_6_7_U116 ( .A(npu_inst_pe_1_6_7_sub_77_carry_3_), .B(
        npu_inst_int_data_res_6__7__3_), .ZN(npu_inst_pe_1_6_7_N68) );
  OR2_X1 npu_inst_pe_1_6_7_U115 ( .A1(npu_inst_int_data_res_6__7__3_), .A2(
        npu_inst_pe_1_6_7_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_6_7_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_6_7_U114 ( .A(npu_inst_pe_1_6_7_sub_77_carry_4_), .B(
        npu_inst_int_data_res_6__7__4_), .ZN(npu_inst_pe_1_6_7_N69) );
  OR2_X1 npu_inst_pe_1_6_7_U113 ( .A1(npu_inst_int_data_res_6__7__4_), .A2(
        npu_inst_pe_1_6_7_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_6_7_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_6_7_U112 ( .A(npu_inst_pe_1_6_7_sub_77_carry_5_), .B(
        npu_inst_int_data_res_6__7__5_), .ZN(npu_inst_pe_1_6_7_N70) );
  OR2_X1 npu_inst_pe_1_6_7_U111 ( .A1(npu_inst_int_data_res_6__7__5_), .A2(
        npu_inst_pe_1_6_7_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_6_7_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_6_7_U110 ( .A(npu_inst_pe_1_6_7_sub_77_carry_6_), .B(
        npu_inst_int_data_res_6__7__6_), .ZN(npu_inst_pe_1_6_7_N71) );
  OR2_X1 npu_inst_pe_1_6_7_U109 ( .A1(npu_inst_int_data_res_6__7__6_), .A2(
        npu_inst_pe_1_6_7_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_6_7_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_6_7_U108 ( .A(npu_inst_int_data_res_6__7__7_), .B(
        npu_inst_pe_1_6_7_sub_77_carry_7_), .ZN(npu_inst_pe_1_6_7_N72) );
  INV_X1 npu_inst_pe_1_6_7_U107 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_6_7_n6)
         );
  INV_X1 npu_inst_pe_1_6_7_U106 ( .A(npu_inst_pe_1_6_7_n6), .ZN(
        npu_inst_pe_1_6_7_n5) );
  INV_X1 npu_inst_pe_1_6_7_U105 ( .A(npu_inst_n35), .ZN(npu_inst_pe_1_6_7_n2)
         );
  AOI22_X1 npu_inst_pe_1_6_7_U104 ( .A1(npu_inst_int_data_y_7__7__0_), .A2(
        npu_inst_pe_1_6_7_n58), .B1(npu_inst_pe_1_6_7_n118), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_6_7_n57) );
  INV_X1 npu_inst_pe_1_6_7_U103 ( .A(npu_inst_pe_1_6_7_n57), .ZN(
        npu_inst_pe_1_6_7_n107) );
  AOI22_X1 npu_inst_pe_1_6_7_U102 ( .A1(npu_inst_int_data_y_7__7__0_), .A2(
        npu_inst_pe_1_6_7_n54), .B1(npu_inst_pe_1_6_7_n117), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_6_7_n53) );
  INV_X1 npu_inst_pe_1_6_7_U99 ( .A(npu_inst_pe_1_6_7_n53), .ZN(
        npu_inst_pe_1_6_7_n108) );
  AOI22_X1 npu_inst_pe_1_6_7_U98 ( .A1(npu_inst_int_data_y_7__7__0_), .A2(
        npu_inst_pe_1_6_7_n50), .B1(npu_inst_pe_1_6_7_n116), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_6_7_n49) );
  INV_X1 npu_inst_pe_1_6_7_U97 ( .A(npu_inst_pe_1_6_7_n49), .ZN(
        npu_inst_pe_1_6_7_n109) );
  AOI22_X1 npu_inst_pe_1_6_7_U96 ( .A1(npu_inst_int_data_y_7__7__0_), .A2(
        npu_inst_pe_1_6_7_n46), .B1(npu_inst_pe_1_6_7_n115), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_6_7_n45) );
  INV_X1 npu_inst_pe_1_6_7_U95 ( .A(npu_inst_pe_1_6_7_n45), .ZN(
        npu_inst_pe_1_6_7_n110) );
  AOI22_X1 npu_inst_pe_1_6_7_U94 ( .A1(npu_inst_int_data_y_7__7__0_), .A2(
        npu_inst_pe_1_6_7_n42), .B1(npu_inst_pe_1_6_7_n114), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_6_7_n41) );
  INV_X1 npu_inst_pe_1_6_7_U93 ( .A(npu_inst_pe_1_6_7_n41), .ZN(
        npu_inst_pe_1_6_7_n111) );
  AOI22_X1 npu_inst_pe_1_6_7_U92 ( .A1(npu_inst_int_data_y_7__7__1_), .A2(
        npu_inst_pe_1_6_7_n58), .B1(npu_inst_pe_1_6_7_n118), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_6_7_n59) );
  INV_X1 npu_inst_pe_1_6_7_U91 ( .A(npu_inst_pe_1_6_7_n59), .ZN(
        npu_inst_pe_1_6_7_n101) );
  AOI22_X1 npu_inst_pe_1_6_7_U90 ( .A1(npu_inst_int_data_y_7__7__1_), .A2(
        npu_inst_pe_1_6_7_n54), .B1(npu_inst_pe_1_6_7_n117), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_6_7_n55) );
  INV_X1 npu_inst_pe_1_6_7_U89 ( .A(npu_inst_pe_1_6_7_n55), .ZN(
        npu_inst_pe_1_6_7_n102) );
  AOI22_X1 npu_inst_pe_1_6_7_U88 ( .A1(npu_inst_int_data_y_7__7__1_), .A2(
        npu_inst_pe_1_6_7_n50), .B1(npu_inst_pe_1_6_7_n116), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_6_7_n51) );
  INV_X1 npu_inst_pe_1_6_7_U87 ( .A(npu_inst_pe_1_6_7_n51), .ZN(
        npu_inst_pe_1_6_7_n103) );
  AOI22_X1 npu_inst_pe_1_6_7_U86 ( .A1(npu_inst_int_data_y_7__7__1_), .A2(
        npu_inst_pe_1_6_7_n46), .B1(npu_inst_pe_1_6_7_n115), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_6_7_n47) );
  INV_X1 npu_inst_pe_1_6_7_U85 ( .A(npu_inst_pe_1_6_7_n47), .ZN(
        npu_inst_pe_1_6_7_n104) );
  AOI22_X1 npu_inst_pe_1_6_7_U84 ( .A1(npu_inst_int_data_y_7__7__1_), .A2(
        npu_inst_pe_1_6_7_n42), .B1(npu_inst_pe_1_6_7_n114), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_6_7_n43) );
  INV_X1 npu_inst_pe_1_6_7_U83 ( .A(npu_inst_pe_1_6_7_n43), .ZN(
        npu_inst_pe_1_6_7_n105) );
  AOI22_X1 npu_inst_pe_1_6_7_U82 ( .A1(npu_inst_pe_1_6_7_n38), .A2(
        npu_inst_int_data_y_7__7__1_), .B1(npu_inst_pe_1_6_7_n113), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_6_7_n39) );
  INV_X1 npu_inst_pe_1_6_7_U81 ( .A(npu_inst_pe_1_6_7_n39), .ZN(
        npu_inst_pe_1_6_7_n106) );
  AND2_X1 npu_inst_pe_1_6_7_U80 ( .A1(npu_inst_pe_1_6_7_N93), .A2(npu_inst_n35), .ZN(npu_inst_int_data_y_6__7__0_) );
  AOI22_X1 npu_inst_pe_1_6_7_U79 ( .A1(npu_inst_pe_1_6_7_n38), .A2(
        npu_inst_int_data_y_7__7__0_), .B1(npu_inst_pe_1_6_7_n113), .B2(
        npu_inst_pe_1_6_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_6_7_n37) );
  INV_X1 npu_inst_pe_1_6_7_U78 ( .A(npu_inst_pe_1_6_7_n37), .ZN(
        npu_inst_pe_1_6_7_n112) );
  AND2_X1 npu_inst_pe_1_6_7_U77 ( .A1(npu_inst_n35), .A2(npu_inst_pe_1_6_7_N94), .ZN(npu_inst_int_data_y_6__7__1_) );
  AOI222_X1 npu_inst_pe_1_6_7_U76 ( .A1(npu_inst_int_data_res_7__7__0_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N73), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N65), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n84) );
  INV_X1 npu_inst_pe_1_6_7_U75 ( .A(npu_inst_pe_1_6_7_n84), .ZN(
        npu_inst_pe_1_6_7_n100) );
  AOI222_X1 npu_inst_pe_1_6_7_U74 ( .A1(npu_inst_pe_1_6_7_n1), .A2(
        npu_inst_int_data_res_7__7__7_), .B1(npu_inst_pe_1_6_7_N80), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N72), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n75) );
  INV_X1 npu_inst_pe_1_6_7_U73 ( .A(npu_inst_pe_1_6_7_n75), .ZN(
        npu_inst_pe_1_6_7_n32) );
  AOI222_X1 npu_inst_pe_1_6_7_U72 ( .A1(npu_inst_int_data_res_7__7__1_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N74), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N66), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n83) );
  INV_X1 npu_inst_pe_1_6_7_U71 ( .A(npu_inst_pe_1_6_7_n83), .ZN(
        npu_inst_pe_1_6_7_n99) );
  AOI222_X1 npu_inst_pe_1_6_7_U70 ( .A1(npu_inst_int_data_res_7__7__3_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N76), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N68), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n81) );
  INV_X1 npu_inst_pe_1_6_7_U69 ( .A(npu_inst_pe_1_6_7_n81), .ZN(
        npu_inst_pe_1_6_7_n36) );
  AOI222_X1 npu_inst_pe_1_6_7_U68 ( .A1(npu_inst_int_data_res_7__7__4_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N77), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N69), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n80) );
  INV_X1 npu_inst_pe_1_6_7_U67 ( .A(npu_inst_pe_1_6_7_n80), .ZN(
        npu_inst_pe_1_6_7_n35) );
  AOI222_X1 npu_inst_pe_1_6_7_U66 ( .A1(npu_inst_int_data_res_7__7__5_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N78), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N70), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n79) );
  INV_X1 npu_inst_pe_1_6_7_U65 ( .A(npu_inst_pe_1_6_7_n79), .ZN(
        npu_inst_pe_1_6_7_n34) );
  AOI222_X1 npu_inst_pe_1_6_7_U64 ( .A1(npu_inst_int_data_res_7__7__6_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N79), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N71), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n78) );
  INV_X1 npu_inst_pe_1_6_7_U63 ( .A(npu_inst_pe_1_6_7_n78), .ZN(
        npu_inst_pe_1_6_7_n33) );
  AND2_X1 npu_inst_pe_1_6_7_U62 ( .A1(npu_inst_int_data_x_6__7__1_), .A2(
        npu_inst_pe_1_6_7_int_q_weight_1_), .ZN(npu_inst_pe_1_6_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_6_7_U61 ( .A1(npu_inst_int_data_x_6__7__0_), .A2(
        npu_inst_pe_1_6_7_int_q_weight_1_), .ZN(npu_inst_pe_1_6_7_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_6_7_U60 ( .A(npu_inst_pe_1_6_7_int_data_1_), .ZN(
        npu_inst_pe_1_6_7_n13) );
  NAND2_X1 npu_inst_pe_1_6_7_U59 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_6_7_n60), .ZN(npu_inst_pe_1_6_7_n74) );
  OAI21_X1 npu_inst_pe_1_6_7_U58 ( .B1(npu_inst_pe_1_6_7_n63), .B2(
        npu_inst_pe_1_6_7_n60), .A(npu_inst_pe_1_6_7_n74), .ZN(
        npu_inst_pe_1_6_7_n97) );
  NAND2_X1 npu_inst_pe_1_6_7_U57 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_6_7_n60), .ZN(npu_inst_pe_1_6_7_n73) );
  OAI21_X1 npu_inst_pe_1_6_7_U56 ( .B1(npu_inst_pe_1_6_7_n61), .B2(
        npu_inst_pe_1_6_7_n60), .A(npu_inst_pe_1_6_7_n73), .ZN(
        npu_inst_pe_1_6_7_n96) );
  NAND2_X1 npu_inst_pe_1_6_7_U55 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_6_7_n56), .ZN(npu_inst_pe_1_6_7_n72) );
  OAI21_X1 npu_inst_pe_1_6_7_U54 ( .B1(npu_inst_pe_1_6_7_n63), .B2(
        npu_inst_pe_1_6_7_n56), .A(npu_inst_pe_1_6_7_n72), .ZN(
        npu_inst_pe_1_6_7_n95) );
  NAND2_X1 npu_inst_pe_1_6_7_U53 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_6_7_n56), .ZN(npu_inst_pe_1_6_7_n71) );
  OAI21_X1 npu_inst_pe_1_6_7_U52 ( .B1(npu_inst_pe_1_6_7_n61), .B2(
        npu_inst_pe_1_6_7_n56), .A(npu_inst_pe_1_6_7_n71), .ZN(
        npu_inst_pe_1_6_7_n94) );
  NAND2_X1 npu_inst_pe_1_6_7_U51 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_6_7_n52), .ZN(npu_inst_pe_1_6_7_n70) );
  OAI21_X1 npu_inst_pe_1_6_7_U50 ( .B1(npu_inst_pe_1_6_7_n63), .B2(
        npu_inst_pe_1_6_7_n52), .A(npu_inst_pe_1_6_7_n70), .ZN(
        npu_inst_pe_1_6_7_n93) );
  NAND2_X1 npu_inst_pe_1_6_7_U49 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_6_7_n52), .ZN(npu_inst_pe_1_6_7_n69) );
  OAI21_X1 npu_inst_pe_1_6_7_U48 ( .B1(npu_inst_pe_1_6_7_n61), .B2(
        npu_inst_pe_1_6_7_n52), .A(npu_inst_pe_1_6_7_n69), .ZN(
        npu_inst_pe_1_6_7_n92) );
  NAND2_X1 npu_inst_pe_1_6_7_U47 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_6_7_n48), .ZN(npu_inst_pe_1_6_7_n68) );
  OAI21_X1 npu_inst_pe_1_6_7_U46 ( .B1(npu_inst_pe_1_6_7_n63), .B2(
        npu_inst_pe_1_6_7_n48), .A(npu_inst_pe_1_6_7_n68), .ZN(
        npu_inst_pe_1_6_7_n91) );
  NAND2_X1 npu_inst_pe_1_6_7_U45 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_6_7_n48), .ZN(npu_inst_pe_1_6_7_n67) );
  OAI21_X1 npu_inst_pe_1_6_7_U44 ( .B1(npu_inst_pe_1_6_7_n61), .B2(
        npu_inst_pe_1_6_7_n48), .A(npu_inst_pe_1_6_7_n67), .ZN(
        npu_inst_pe_1_6_7_n90) );
  NAND2_X1 npu_inst_pe_1_6_7_U43 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_6_7_n44), .ZN(npu_inst_pe_1_6_7_n66) );
  OAI21_X1 npu_inst_pe_1_6_7_U42 ( .B1(npu_inst_pe_1_6_7_n63), .B2(
        npu_inst_pe_1_6_7_n44), .A(npu_inst_pe_1_6_7_n66), .ZN(
        npu_inst_pe_1_6_7_n89) );
  NAND2_X1 npu_inst_pe_1_6_7_U41 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_6_7_n44), .ZN(npu_inst_pe_1_6_7_n65) );
  OAI21_X1 npu_inst_pe_1_6_7_U40 ( .B1(npu_inst_pe_1_6_7_n61), .B2(
        npu_inst_pe_1_6_7_n44), .A(npu_inst_pe_1_6_7_n65), .ZN(
        npu_inst_pe_1_6_7_n88) );
  NAND2_X1 npu_inst_pe_1_6_7_U39 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_6_7_n40), .ZN(npu_inst_pe_1_6_7_n64) );
  OAI21_X1 npu_inst_pe_1_6_7_U38 ( .B1(npu_inst_pe_1_6_7_n63), .B2(
        npu_inst_pe_1_6_7_n40), .A(npu_inst_pe_1_6_7_n64), .ZN(
        npu_inst_pe_1_6_7_n87) );
  NAND2_X1 npu_inst_pe_1_6_7_U37 ( .A1(npu_inst_pe_1_6_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_6_7_n40), .ZN(npu_inst_pe_1_6_7_n62) );
  OAI21_X1 npu_inst_pe_1_6_7_U36 ( .B1(npu_inst_pe_1_6_7_n61), .B2(
        npu_inst_pe_1_6_7_n40), .A(npu_inst_pe_1_6_7_n62), .ZN(
        npu_inst_pe_1_6_7_n86) );
  NOR3_X1 npu_inst_pe_1_6_7_U35 ( .A1(npu_inst_pe_1_6_7_n26), .A2(npu_inst_n35), .A3(npu_inst_int_ckg[8]), .ZN(npu_inst_pe_1_6_7_n85) );
  OR2_X1 npu_inst_pe_1_6_7_U34 ( .A1(npu_inst_pe_1_6_7_n85), .A2(
        npu_inst_pe_1_6_7_n1), .ZN(npu_inst_pe_1_6_7_N84) );
  AOI222_X1 npu_inst_pe_1_6_7_U33 ( .A1(npu_inst_int_data_res_7__7__2_), .A2(
        npu_inst_pe_1_6_7_n1), .B1(npu_inst_pe_1_6_7_N75), .B2(
        npu_inst_pe_1_6_7_n76), .C1(npu_inst_pe_1_6_7_N67), .C2(
        npu_inst_pe_1_6_7_n77), .ZN(npu_inst_pe_1_6_7_n82) );
  INV_X1 npu_inst_pe_1_6_7_U32 ( .A(npu_inst_pe_1_6_7_n82), .ZN(
        npu_inst_pe_1_6_7_n98) );
  INV_X1 npu_inst_pe_1_6_7_U31 ( .A(npu_inst_pe_1_6_7_int_data_0_), .ZN(
        npu_inst_pe_1_6_7_n12) );
  INV_X1 npu_inst_pe_1_6_7_U30 ( .A(npu_inst_n49), .ZN(npu_inst_pe_1_6_7_n4)
         );
  AOI22_X1 npu_inst_pe_1_6_7_U29 ( .A1(npu_inst_n35), .A2(
        npu_inst_int_data_y_7__7__1_), .B1(npu_inst_pe_1_6_7_n2), .B2(
        int_i_data_h_npu[3]), .ZN(npu_inst_pe_1_6_7_n63) );
  AOI22_X1 npu_inst_pe_1_6_7_U28 ( .A1(npu_inst_n35), .A2(
        npu_inst_int_data_y_7__7__0_), .B1(npu_inst_pe_1_6_7_n2), .B2(
        int_i_data_h_npu[2]), .ZN(npu_inst_pe_1_6_7_n61) );
  OR3_X1 npu_inst_pe_1_6_7_U27 ( .A1(npu_inst_pe_1_6_7_n5), .A2(
        npu_inst_pe_1_6_7_n7), .A3(npu_inst_pe_1_6_7_n4), .ZN(
        npu_inst_pe_1_6_7_n56) );
  OR3_X1 npu_inst_pe_1_6_7_U26 ( .A1(npu_inst_pe_1_6_7_n4), .A2(
        npu_inst_pe_1_6_7_n7), .A3(npu_inst_pe_1_6_7_n6), .ZN(
        npu_inst_pe_1_6_7_n48) );
  INV_X1 npu_inst_pe_1_6_7_U25 ( .A(npu_inst_pe_1_6_7_n4), .ZN(
        npu_inst_pe_1_6_7_n3) );
  OR3_X1 npu_inst_pe_1_6_7_U24 ( .A1(npu_inst_pe_1_6_7_n3), .A2(
        npu_inst_pe_1_6_7_n7), .A3(npu_inst_pe_1_6_7_n6), .ZN(
        npu_inst_pe_1_6_7_n52) );
  OR3_X1 npu_inst_pe_1_6_7_U23 ( .A1(npu_inst_pe_1_6_7_n5), .A2(
        npu_inst_pe_1_6_7_n7), .A3(npu_inst_pe_1_6_7_n3), .ZN(
        npu_inst_pe_1_6_7_n60) );
  BUF_X1 npu_inst_pe_1_6_7_U22 ( .A(npu_inst_n13), .Z(npu_inst_pe_1_6_7_n1) );
  NOR2_X1 npu_inst_pe_1_6_7_U21 ( .A1(npu_inst_pe_1_6_7_n60), .A2(
        npu_inst_pe_1_6_7_n2), .ZN(npu_inst_pe_1_6_7_n58) );
  NOR2_X1 npu_inst_pe_1_6_7_U20 ( .A1(npu_inst_pe_1_6_7_n56), .A2(
        npu_inst_pe_1_6_7_n2), .ZN(npu_inst_pe_1_6_7_n54) );
  NOR2_X1 npu_inst_pe_1_6_7_U19 ( .A1(npu_inst_pe_1_6_7_n52), .A2(
        npu_inst_pe_1_6_7_n2), .ZN(npu_inst_pe_1_6_7_n50) );
  NOR2_X1 npu_inst_pe_1_6_7_U18 ( .A1(npu_inst_pe_1_6_7_n48), .A2(
        npu_inst_pe_1_6_7_n2), .ZN(npu_inst_pe_1_6_7_n46) );
  NOR2_X1 npu_inst_pe_1_6_7_U17 ( .A1(npu_inst_pe_1_6_7_n40), .A2(
        npu_inst_pe_1_6_7_n2), .ZN(npu_inst_pe_1_6_7_n38) );
  NOR2_X1 npu_inst_pe_1_6_7_U16 ( .A1(npu_inst_pe_1_6_7_n44), .A2(
        npu_inst_pe_1_6_7_n2), .ZN(npu_inst_pe_1_6_7_n42) );
  BUF_X1 npu_inst_pe_1_6_7_U15 ( .A(npu_inst_n76), .Z(npu_inst_pe_1_6_7_n7) );
  INV_X1 npu_inst_pe_1_6_7_U14 ( .A(npu_inst_n104), .ZN(npu_inst_pe_1_6_7_n11)
         );
  INV_X1 npu_inst_pe_1_6_7_U13 ( .A(npu_inst_pe_1_6_7_n38), .ZN(
        npu_inst_pe_1_6_7_n113) );
  INV_X1 npu_inst_pe_1_6_7_U12 ( .A(npu_inst_pe_1_6_7_n58), .ZN(
        npu_inst_pe_1_6_7_n118) );
  INV_X1 npu_inst_pe_1_6_7_U11 ( .A(npu_inst_pe_1_6_7_n54), .ZN(
        npu_inst_pe_1_6_7_n117) );
  INV_X1 npu_inst_pe_1_6_7_U10 ( .A(npu_inst_pe_1_6_7_n50), .ZN(
        npu_inst_pe_1_6_7_n116) );
  INV_X1 npu_inst_pe_1_6_7_U9 ( .A(npu_inst_pe_1_6_7_n46), .ZN(
        npu_inst_pe_1_6_7_n115) );
  INV_X1 npu_inst_pe_1_6_7_U8 ( .A(npu_inst_pe_1_6_7_n42), .ZN(
        npu_inst_pe_1_6_7_n114) );
  BUF_X1 npu_inst_pe_1_6_7_U7 ( .A(npu_inst_pe_1_6_7_n11), .Z(
        npu_inst_pe_1_6_7_n10) );
  BUF_X1 npu_inst_pe_1_6_7_U6 ( .A(npu_inst_pe_1_6_7_n11), .Z(
        npu_inst_pe_1_6_7_n9) );
  BUF_X1 npu_inst_pe_1_6_7_U5 ( .A(npu_inst_pe_1_6_7_n11), .Z(
        npu_inst_pe_1_6_7_n8) );
  NOR2_X1 npu_inst_pe_1_6_7_U4 ( .A1(npu_inst_pe_1_6_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_6_7_n1), .ZN(npu_inst_pe_1_6_7_n76) );
  NOR2_X1 npu_inst_pe_1_6_7_U3 ( .A1(npu_inst_pe_1_6_7_n27), .A2(
        npu_inst_pe_1_6_7_n1), .ZN(npu_inst_pe_1_6_7_n77) );
  FA_X1 npu_inst_pe_1_6_7_sub_77_U2_1 ( .A(npu_inst_int_data_res_6__7__1_), 
        .B(npu_inst_pe_1_6_7_n13), .CI(npu_inst_pe_1_6_7_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_6_7_sub_77_carry_2_), .S(npu_inst_pe_1_6_7_N66) );
  FA_X1 npu_inst_pe_1_6_7_add_79_U1_1 ( .A(npu_inst_int_data_res_6__7__1_), 
        .B(npu_inst_pe_1_6_7_int_data_1_), .CI(
        npu_inst_pe_1_6_7_add_79_carry_1_), .CO(
        npu_inst_pe_1_6_7_add_79_carry_2_), .S(npu_inst_pe_1_6_7_N74) );
  NAND3_X1 npu_inst_pe_1_6_7_U101 ( .A1(npu_inst_pe_1_6_7_n4), .A2(
        npu_inst_pe_1_6_7_n6), .A3(npu_inst_pe_1_6_7_n7), .ZN(
        npu_inst_pe_1_6_7_n44) );
  NAND3_X1 npu_inst_pe_1_6_7_U100 ( .A1(npu_inst_pe_1_6_7_n3), .A2(
        npu_inst_pe_1_6_7_n6), .A3(npu_inst_pe_1_6_7_n7), .ZN(
        npu_inst_pe_1_6_7_n40) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_6_7_n33), .CK(
        npu_inst_pe_1_6_7_net3213), .RN(npu_inst_pe_1_6_7_n8), .Q(
        npu_inst_int_data_res_6__7__6_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_6_7_n34), .CK(
        npu_inst_pe_1_6_7_net3213), .RN(npu_inst_pe_1_6_7_n8), .Q(
        npu_inst_int_data_res_6__7__5_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_6_7_n35), .CK(
        npu_inst_pe_1_6_7_net3213), .RN(npu_inst_pe_1_6_7_n8), .Q(
        npu_inst_int_data_res_6__7__4_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_6_7_n36), .CK(
        npu_inst_pe_1_6_7_net3213), .RN(npu_inst_pe_1_6_7_n8), .Q(
        npu_inst_int_data_res_6__7__3_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_6_7_n98), .CK(
        npu_inst_pe_1_6_7_net3213), .RN(npu_inst_pe_1_6_7_n8), .Q(
        npu_inst_int_data_res_6__7__2_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_6_7_n99), .CK(
        npu_inst_pe_1_6_7_net3213), .RN(npu_inst_pe_1_6_7_n8), .Q(
        npu_inst_int_data_res_6__7__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_6_7_n32), .CK(
        npu_inst_pe_1_6_7_net3213), .RN(npu_inst_pe_1_6_7_n8), .Q(
        npu_inst_int_data_res_6__7__7_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_6_7_n100), 
        .CK(npu_inst_pe_1_6_7_net3213), .RN(npu_inst_pe_1_6_7_n8), .Q(
        npu_inst_int_data_res_6__7__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_weight_reg_0_ ( .D(npu_inst_n90), .CK(
        npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n8), .Q(
        npu_inst_pe_1_6_7_int_q_weight_0_), .QN(npu_inst_pe_1_6_7_n27) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_weight_reg_1_ ( .D(npu_inst_n96), .CK(
        npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n8), .Q(
        npu_inst_pe_1_6_7_int_q_weight_1_), .QN(npu_inst_pe_1_6_7_n26) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_6_7_n112), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n8), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_6_7_n106), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n8), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_6_7_n111), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_6_7_n105), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_6_7_n110), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_6_7_n104), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_6_7_n109), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_6_7_n103), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_6_7_n108), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_6_7_n102), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_6_7_n107), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_6_7_n101), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_6_7_n86), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_6_7_n87), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n9), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_6_7_n88), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_6_7_n89), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_6_7_n90), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_6_7_n91), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_6_7_n92), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_6_7_n93), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_6_7_n94), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_6_7_n95), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_6_7_n96), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_6_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_6_7_n97), 
        .CK(npu_inst_pe_1_6_7_net3219), .RN(npu_inst_pe_1_6_7_n10), .Q(
        npu_inst_pe_1_6_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_6_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_6_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_6_7_net3213) );
  CLKGATETST_X1 npu_inst_pe_1_6_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n43), .SE(1'b0), .GCK(npu_inst_pe_1_6_7_net3219) );
  MUX2_X1 npu_inst_pe_1_7_0_U153 ( .A(npu_inst_pe_1_7_0_n31), .B(
        npu_inst_pe_1_7_0_n28), .S(npu_inst_pe_1_7_0_n7), .Z(
        npu_inst_pe_1_7_0_N93) );
  MUX2_X1 npu_inst_pe_1_7_0_U152 ( .A(npu_inst_pe_1_7_0_n30), .B(
        npu_inst_pe_1_7_0_n29), .S(npu_inst_pe_1_7_0_n5), .Z(
        npu_inst_pe_1_7_0_n31) );
  MUX2_X1 npu_inst_pe_1_7_0_U151 ( .A(npu_inst_pe_1_7_0_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_0_n3), .Z(
        npu_inst_pe_1_7_0_n30) );
  MUX2_X1 npu_inst_pe_1_7_0_U150 ( .A(npu_inst_pe_1_7_0_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_0_n3), .Z(
        npu_inst_pe_1_7_0_n29) );
  MUX2_X1 npu_inst_pe_1_7_0_U149 ( .A(npu_inst_pe_1_7_0_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_0_n3), .Z(
        npu_inst_pe_1_7_0_n28) );
  MUX2_X1 npu_inst_pe_1_7_0_U148 ( .A(npu_inst_pe_1_7_0_n25), .B(
        npu_inst_pe_1_7_0_n22), .S(npu_inst_pe_1_7_0_n7), .Z(
        npu_inst_pe_1_7_0_N94) );
  MUX2_X1 npu_inst_pe_1_7_0_U147 ( .A(npu_inst_pe_1_7_0_n24), .B(
        npu_inst_pe_1_7_0_n23), .S(npu_inst_pe_1_7_0_n5), .Z(
        npu_inst_pe_1_7_0_n25) );
  MUX2_X1 npu_inst_pe_1_7_0_U146 ( .A(npu_inst_pe_1_7_0_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_0_n3), .Z(
        npu_inst_pe_1_7_0_n24) );
  MUX2_X1 npu_inst_pe_1_7_0_U145 ( .A(npu_inst_pe_1_7_0_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_0_n3), .Z(
        npu_inst_pe_1_7_0_n23) );
  MUX2_X1 npu_inst_pe_1_7_0_U144 ( .A(npu_inst_pe_1_7_0_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_0_n3), .Z(
        npu_inst_pe_1_7_0_n22) );
  MUX2_X1 npu_inst_pe_1_7_0_U143 ( .A(npu_inst_pe_1_7_0_n21), .B(
        npu_inst_pe_1_7_0_n18), .S(npu_inst_pe_1_7_0_n7), .Z(
        npu_inst_pe_1_7_0_o_data_h_1_) );
  MUX2_X1 npu_inst_pe_1_7_0_U142 ( .A(npu_inst_pe_1_7_0_n20), .B(
        npu_inst_pe_1_7_0_n19), .S(npu_inst_pe_1_7_0_n5), .Z(
        npu_inst_pe_1_7_0_n21) );
  MUX2_X1 npu_inst_pe_1_7_0_U141 ( .A(npu_inst_pe_1_7_0_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_0_n3), .Z(
        npu_inst_pe_1_7_0_n20) );
  MUX2_X1 npu_inst_pe_1_7_0_U140 ( .A(npu_inst_pe_1_7_0_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_0_n3), .Z(
        npu_inst_pe_1_7_0_n19) );
  MUX2_X1 npu_inst_pe_1_7_0_U139 ( .A(npu_inst_pe_1_7_0_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_0_n3), .Z(
        npu_inst_pe_1_7_0_n18) );
  MUX2_X1 npu_inst_pe_1_7_0_U138 ( .A(npu_inst_pe_1_7_0_n17), .B(
        npu_inst_pe_1_7_0_n14), .S(npu_inst_pe_1_7_0_n7), .Z(
        npu_inst_pe_1_7_0_o_data_h_0_) );
  MUX2_X1 npu_inst_pe_1_7_0_U137 ( .A(npu_inst_pe_1_7_0_n16), .B(
        npu_inst_pe_1_7_0_n15), .S(npu_inst_pe_1_7_0_n5), .Z(
        npu_inst_pe_1_7_0_n17) );
  MUX2_X1 npu_inst_pe_1_7_0_U136 ( .A(npu_inst_pe_1_7_0_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_0_n3), .Z(
        npu_inst_pe_1_7_0_n16) );
  MUX2_X1 npu_inst_pe_1_7_0_U135 ( .A(npu_inst_pe_1_7_0_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_0_n3), .Z(
        npu_inst_pe_1_7_0_n15) );
  MUX2_X1 npu_inst_pe_1_7_0_U134 ( .A(npu_inst_pe_1_7_0_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_0_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_0_n3), .Z(
        npu_inst_pe_1_7_0_n14) );
  XOR2_X1 npu_inst_pe_1_7_0_U133 ( .A(npu_inst_pe_1_7_0_int_data_0_), .B(
        npu_inst_int_data_res_7__0__0_), .Z(npu_inst_pe_1_7_0_N73) );
  AND2_X1 npu_inst_pe_1_7_0_U132 ( .A1(npu_inst_int_data_res_7__0__0_), .A2(
        npu_inst_pe_1_7_0_int_data_0_), .ZN(npu_inst_pe_1_7_0_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_0_U131 ( .A(npu_inst_int_data_res_7__0__0_), .B(
        npu_inst_pe_1_7_0_n12), .ZN(npu_inst_pe_1_7_0_N65) );
  OR2_X1 npu_inst_pe_1_7_0_U130 ( .A1(npu_inst_pe_1_7_0_n12), .A2(
        npu_inst_int_data_res_7__0__0_), .ZN(npu_inst_pe_1_7_0_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_0_U129 ( .A(npu_inst_int_data_res_7__0__2_), .B(
        npu_inst_pe_1_7_0_add_79_carry_2_), .Z(npu_inst_pe_1_7_0_N75) );
  AND2_X1 npu_inst_pe_1_7_0_U128 ( .A1(npu_inst_pe_1_7_0_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_7__0__2_), .ZN(
        npu_inst_pe_1_7_0_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_0_U127 ( .A(npu_inst_int_data_res_7__0__3_), .B(
        npu_inst_pe_1_7_0_add_79_carry_3_), .Z(npu_inst_pe_1_7_0_N76) );
  AND2_X1 npu_inst_pe_1_7_0_U126 ( .A1(npu_inst_pe_1_7_0_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_7__0__3_), .ZN(
        npu_inst_pe_1_7_0_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_0_U125 ( .A(npu_inst_int_data_res_7__0__4_), .B(
        npu_inst_pe_1_7_0_add_79_carry_4_), .Z(npu_inst_pe_1_7_0_N77) );
  AND2_X1 npu_inst_pe_1_7_0_U124 ( .A1(npu_inst_pe_1_7_0_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_7__0__4_), .ZN(
        npu_inst_pe_1_7_0_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_0_U123 ( .A(npu_inst_int_data_res_7__0__5_), .B(
        npu_inst_pe_1_7_0_add_79_carry_5_), .Z(npu_inst_pe_1_7_0_N78) );
  AND2_X1 npu_inst_pe_1_7_0_U122 ( .A1(npu_inst_pe_1_7_0_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_7__0__5_), .ZN(
        npu_inst_pe_1_7_0_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_0_U121 ( .A(npu_inst_int_data_res_7__0__6_), .B(
        npu_inst_pe_1_7_0_add_79_carry_6_), .Z(npu_inst_pe_1_7_0_N79) );
  AND2_X1 npu_inst_pe_1_7_0_U120 ( .A1(npu_inst_pe_1_7_0_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_7__0__6_), .ZN(
        npu_inst_pe_1_7_0_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_0_U119 ( .A(npu_inst_int_data_res_7__0__7_), .B(
        npu_inst_pe_1_7_0_add_79_carry_7_), .Z(npu_inst_pe_1_7_0_N80) );
  XNOR2_X1 npu_inst_pe_1_7_0_U118 ( .A(npu_inst_pe_1_7_0_sub_77_carry_2_), .B(
        npu_inst_int_data_res_7__0__2_), .ZN(npu_inst_pe_1_7_0_N67) );
  OR2_X1 npu_inst_pe_1_7_0_U117 ( .A1(npu_inst_int_data_res_7__0__2_), .A2(
        npu_inst_pe_1_7_0_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_7_0_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_0_U116 ( .A(npu_inst_pe_1_7_0_sub_77_carry_3_), .B(
        npu_inst_int_data_res_7__0__3_), .ZN(npu_inst_pe_1_7_0_N68) );
  OR2_X1 npu_inst_pe_1_7_0_U115 ( .A1(npu_inst_int_data_res_7__0__3_), .A2(
        npu_inst_pe_1_7_0_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_7_0_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_0_U114 ( .A(npu_inst_pe_1_7_0_sub_77_carry_4_), .B(
        npu_inst_int_data_res_7__0__4_), .ZN(npu_inst_pe_1_7_0_N69) );
  OR2_X1 npu_inst_pe_1_7_0_U113 ( .A1(npu_inst_int_data_res_7__0__4_), .A2(
        npu_inst_pe_1_7_0_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_7_0_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_0_U112 ( .A(npu_inst_pe_1_7_0_sub_77_carry_5_), .B(
        npu_inst_int_data_res_7__0__5_), .ZN(npu_inst_pe_1_7_0_N70) );
  OR2_X1 npu_inst_pe_1_7_0_U111 ( .A1(npu_inst_int_data_res_7__0__5_), .A2(
        npu_inst_pe_1_7_0_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_7_0_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_0_U110 ( .A(npu_inst_pe_1_7_0_sub_77_carry_6_), .B(
        npu_inst_int_data_res_7__0__6_), .ZN(npu_inst_pe_1_7_0_N71) );
  OR2_X1 npu_inst_pe_1_7_0_U109 ( .A1(npu_inst_int_data_res_7__0__6_), .A2(
        npu_inst_pe_1_7_0_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_7_0_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_0_U108 ( .A(npu_inst_int_data_res_7__0__7_), .B(
        npu_inst_pe_1_7_0_sub_77_carry_7_), .ZN(npu_inst_pe_1_7_0_N72) );
  INV_X1 npu_inst_pe_1_7_0_U107 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_7_0_n6)
         );
  INV_X1 npu_inst_pe_1_7_0_U106 ( .A(npu_inst_pe_1_7_0_n6), .ZN(
        npu_inst_pe_1_7_0_n5) );
  INV_X1 npu_inst_pe_1_7_0_U105 ( .A(npu_inst_n35), .ZN(npu_inst_pe_1_7_0_n2)
         );
  AOI22_X1 npu_inst_pe_1_7_0_U104 ( .A1(npu_inst_pe_1_7_0_n38), .A2(
        int_i_data_v_npu[15]), .B1(npu_inst_pe_1_7_0_n113), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_0_n39) );
  INV_X1 npu_inst_pe_1_7_0_U103 ( .A(npu_inst_pe_1_7_0_n39), .ZN(
        npu_inst_pe_1_7_0_n111) );
  AOI22_X1 npu_inst_pe_1_7_0_U102 ( .A1(npu_inst_pe_1_7_0_n38), .A2(
        int_i_data_v_npu[14]), .B1(npu_inst_pe_1_7_0_n113), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_0_n37) );
  INV_X1 npu_inst_pe_1_7_0_U99 ( .A(npu_inst_pe_1_7_0_n37), .ZN(
        npu_inst_pe_1_7_0_n112) );
  AOI22_X1 npu_inst_pe_1_7_0_U98 ( .A1(int_i_data_v_npu[15]), .A2(
        npu_inst_pe_1_7_0_n58), .B1(npu_inst_pe_1_7_0_n118), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_0_n59) );
  INV_X1 npu_inst_pe_1_7_0_U97 ( .A(npu_inst_pe_1_7_0_n59), .ZN(
        npu_inst_pe_1_7_0_n101) );
  AOI22_X1 npu_inst_pe_1_7_0_U96 ( .A1(int_i_data_v_npu[14]), .A2(
        npu_inst_pe_1_7_0_n58), .B1(npu_inst_pe_1_7_0_n118), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_0_n57) );
  INV_X1 npu_inst_pe_1_7_0_U95 ( .A(npu_inst_pe_1_7_0_n57), .ZN(
        npu_inst_pe_1_7_0_n102) );
  AOI22_X1 npu_inst_pe_1_7_0_U94 ( .A1(int_i_data_v_npu[15]), .A2(
        npu_inst_pe_1_7_0_n54), .B1(npu_inst_pe_1_7_0_n117), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_0_n55) );
  INV_X1 npu_inst_pe_1_7_0_U93 ( .A(npu_inst_pe_1_7_0_n55), .ZN(
        npu_inst_pe_1_7_0_n103) );
  AOI22_X1 npu_inst_pe_1_7_0_U92 ( .A1(int_i_data_v_npu[14]), .A2(
        npu_inst_pe_1_7_0_n54), .B1(npu_inst_pe_1_7_0_n117), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_0_n53) );
  INV_X1 npu_inst_pe_1_7_0_U91 ( .A(npu_inst_pe_1_7_0_n53), .ZN(
        npu_inst_pe_1_7_0_n104) );
  AOI22_X1 npu_inst_pe_1_7_0_U90 ( .A1(int_i_data_v_npu[15]), .A2(
        npu_inst_pe_1_7_0_n50), .B1(npu_inst_pe_1_7_0_n116), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_0_n51) );
  INV_X1 npu_inst_pe_1_7_0_U89 ( .A(npu_inst_pe_1_7_0_n51), .ZN(
        npu_inst_pe_1_7_0_n105) );
  AOI22_X1 npu_inst_pe_1_7_0_U88 ( .A1(int_i_data_v_npu[14]), .A2(
        npu_inst_pe_1_7_0_n50), .B1(npu_inst_pe_1_7_0_n116), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_0_n49) );
  INV_X1 npu_inst_pe_1_7_0_U87 ( .A(npu_inst_pe_1_7_0_n49), .ZN(
        npu_inst_pe_1_7_0_n106) );
  AOI22_X1 npu_inst_pe_1_7_0_U86 ( .A1(int_i_data_v_npu[15]), .A2(
        npu_inst_pe_1_7_0_n46), .B1(npu_inst_pe_1_7_0_n115), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_0_n47) );
  INV_X1 npu_inst_pe_1_7_0_U85 ( .A(npu_inst_pe_1_7_0_n47), .ZN(
        npu_inst_pe_1_7_0_n107) );
  AOI22_X1 npu_inst_pe_1_7_0_U84 ( .A1(int_i_data_v_npu[14]), .A2(
        npu_inst_pe_1_7_0_n46), .B1(npu_inst_pe_1_7_0_n115), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_0_n45) );
  INV_X1 npu_inst_pe_1_7_0_U83 ( .A(npu_inst_pe_1_7_0_n45), .ZN(
        npu_inst_pe_1_7_0_n108) );
  AOI22_X1 npu_inst_pe_1_7_0_U82 ( .A1(int_i_data_v_npu[15]), .A2(
        npu_inst_pe_1_7_0_n42), .B1(npu_inst_pe_1_7_0_n114), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_0_n43) );
  INV_X1 npu_inst_pe_1_7_0_U81 ( .A(npu_inst_pe_1_7_0_n43), .ZN(
        npu_inst_pe_1_7_0_n109) );
  AOI22_X1 npu_inst_pe_1_7_0_U80 ( .A1(int_i_data_v_npu[14]), .A2(
        npu_inst_pe_1_7_0_n42), .B1(npu_inst_pe_1_7_0_n114), .B2(
        npu_inst_pe_1_7_0_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_0_n41) );
  INV_X1 npu_inst_pe_1_7_0_U79 ( .A(npu_inst_pe_1_7_0_n41), .ZN(
        npu_inst_pe_1_7_0_n110) );
  AND2_X1 npu_inst_pe_1_7_0_U78 ( .A1(npu_inst_pe_1_7_0_N93), .A2(npu_inst_n35), .ZN(npu_inst_int_data_y_7__0__0_) );
  NAND2_X1 npu_inst_pe_1_7_0_U77 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_0_n60), .ZN(npu_inst_pe_1_7_0_n74) );
  OAI21_X1 npu_inst_pe_1_7_0_U76 ( .B1(npu_inst_pe_1_7_0_n63), .B2(
        npu_inst_pe_1_7_0_n60), .A(npu_inst_pe_1_7_0_n74), .ZN(
        npu_inst_pe_1_7_0_n97) );
  NAND2_X1 npu_inst_pe_1_7_0_U75 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_0_n60), .ZN(npu_inst_pe_1_7_0_n73) );
  OAI21_X1 npu_inst_pe_1_7_0_U74 ( .B1(npu_inst_pe_1_7_0_n61), .B2(
        npu_inst_pe_1_7_0_n60), .A(npu_inst_pe_1_7_0_n73), .ZN(
        npu_inst_pe_1_7_0_n96) );
  NAND2_X1 npu_inst_pe_1_7_0_U73 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_0_n56), .ZN(npu_inst_pe_1_7_0_n72) );
  OAI21_X1 npu_inst_pe_1_7_0_U72 ( .B1(npu_inst_pe_1_7_0_n63), .B2(
        npu_inst_pe_1_7_0_n56), .A(npu_inst_pe_1_7_0_n72), .ZN(
        npu_inst_pe_1_7_0_n95) );
  NAND2_X1 npu_inst_pe_1_7_0_U71 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_0_n56), .ZN(npu_inst_pe_1_7_0_n71) );
  OAI21_X1 npu_inst_pe_1_7_0_U70 ( .B1(npu_inst_pe_1_7_0_n61), .B2(
        npu_inst_pe_1_7_0_n56), .A(npu_inst_pe_1_7_0_n71), .ZN(
        npu_inst_pe_1_7_0_n94) );
  NAND2_X1 npu_inst_pe_1_7_0_U69 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_0_n52), .ZN(npu_inst_pe_1_7_0_n70) );
  OAI21_X1 npu_inst_pe_1_7_0_U68 ( .B1(npu_inst_pe_1_7_0_n63), .B2(
        npu_inst_pe_1_7_0_n52), .A(npu_inst_pe_1_7_0_n70), .ZN(
        npu_inst_pe_1_7_0_n93) );
  NAND2_X1 npu_inst_pe_1_7_0_U67 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_0_n52), .ZN(npu_inst_pe_1_7_0_n69) );
  OAI21_X1 npu_inst_pe_1_7_0_U66 ( .B1(npu_inst_pe_1_7_0_n61), .B2(
        npu_inst_pe_1_7_0_n52), .A(npu_inst_pe_1_7_0_n69), .ZN(
        npu_inst_pe_1_7_0_n92) );
  NAND2_X1 npu_inst_pe_1_7_0_U65 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_0_n48), .ZN(npu_inst_pe_1_7_0_n68) );
  OAI21_X1 npu_inst_pe_1_7_0_U64 ( .B1(npu_inst_pe_1_7_0_n63), .B2(
        npu_inst_pe_1_7_0_n48), .A(npu_inst_pe_1_7_0_n68), .ZN(
        npu_inst_pe_1_7_0_n91) );
  NAND2_X1 npu_inst_pe_1_7_0_U63 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_0_n48), .ZN(npu_inst_pe_1_7_0_n67) );
  OAI21_X1 npu_inst_pe_1_7_0_U62 ( .B1(npu_inst_pe_1_7_0_n61), .B2(
        npu_inst_pe_1_7_0_n48), .A(npu_inst_pe_1_7_0_n67), .ZN(
        npu_inst_pe_1_7_0_n90) );
  NAND2_X1 npu_inst_pe_1_7_0_U61 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_0_n44), .ZN(npu_inst_pe_1_7_0_n66) );
  OAI21_X1 npu_inst_pe_1_7_0_U60 ( .B1(npu_inst_pe_1_7_0_n63), .B2(
        npu_inst_pe_1_7_0_n44), .A(npu_inst_pe_1_7_0_n66), .ZN(
        npu_inst_pe_1_7_0_n89) );
  NAND2_X1 npu_inst_pe_1_7_0_U59 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_0_n44), .ZN(npu_inst_pe_1_7_0_n65) );
  OAI21_X1 npu_inst_pe_1_7_0_U58 ( .B1(npu_inst_pe_1_7_0_n61), .B2(
        npu_inst_pe_1_7_0_n44), .A(npu_inst_pe_1_7_0_n65), .ZN(
        npu_inst_pe_1_7_0_n88) );
  NAND2_X1 npu_inst_pe_1_7_0_U57 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_0_n40), .ZN(npu_inst_pe_1_7_0_n64) );
  OAI21_X1 npu_inst_pe_1_7_0_U56 ( .B1(npu_inst_pe_1_7_0_n63), .B2(
        npu_inst_pe_1_7_0_n40), .A(npu_inst_pe_1_7_0_n64), .ZN(
        npu_inst_pe_1_7_0_n87) );
  NAND2_X1 npu_inst_pe_1_7_0_U55 ( .A1(npu_inst_pe_1_7_0_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_0_n40), .ZN(npu_inst_pe_1_7_0_n62) );
  OAI21_X1 npu_inst_pe_1_7_0_U54 ( .B1(npu_inst_pe_1_7_0_n61), .B2(
        npu_inst_pe_1_7_0_n40), .A(npu_inst_pe_1_7_0_n62), .ZN(
        npu_inst_pe_1_7_0_n86) );
  AND2_X1 npu_inst_pe_1_7_0_U53 ( .A1(npu_inst_n35), .A2(npu_inst_pe_1_7_0_N94), .ZN(npu_inst_int_data_y_7__0__1_) );
  AOI22_X1 npu_inst_pe_1_7_0_U52 ( .A1(npu_inst_n35), .A2(int_i_data_v_npu[15]), .B1(npu_inst_pe_1_7_0_n2), .B2(npu_inst_int_data_x_7__1__1_), .ZN(
        npu_inst_pe_1_7_0_n63) );
  AOI22_X1 npu_inst_pe_1_7_0_U51 ( .A1(npu_inst_n35), .A2(int_i_data_v_npu[14]), .B1(npu_inst_pe_1_7_0_n2), .B2(npu_inst_int_data_x_7__1__0_), .ZN(
        npu_inst_pe_1_7_0_n61) );
  AOI222_X1 npu_inst_pe_1_7_0_U50 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N73), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N65), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n84) );
  INV_X1 npu_inst_pe_1_7_0_U49 ( .A(npu_inst_pe_1_7_0_n84), .ZN(
        npu_inst_pe_1_7_0_n100) );
  AOI222_X1 npu_inst_pe_1_7_0_U48 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N74), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N66), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n83) );
  INV_X1 npu_inst_pe_1_7_0_U47 ( .A(npu_inst_pe_1_7_0_n83), .ZN(
        npu_inst_pe_1_7_0_n99) );
  AOI222_X1 npu_inst_pe_1_7_0_U46 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N75), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N67), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n82) );
  INV_X1 npu_inst_pe_1_7_0_U45 ( .A(npu_inst_pe_1_7_0_n82), .ZN(
        npu_inst_pe_1_7_0_n98) );
  AOI222_X1 npu_inst_pe_1_7_0_U44 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N76), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N68), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n81) );
  INV_X1 npu_inst_pe_1_7_0_U43 ( .A(npu_inst_pe_1_7_0_n81), .ZN(
        npu_inst_pe_1_7_0_n36) );
  AOI222_X1 npu_inst_pe_1_7_0_U42 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N77), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N69), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n80) );
  INV_X1 npu_inst_pe_1_7_0_U41 ( .A(npu_inst_pe_1_7_0_n80), .ZN(
        npu_inst_pe_1_7_0_n35) );
  AOI222_X1 npu_inst_pe_1_7_0_U40 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N78), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N70), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n79) );
  INV_X1 npu_inst_pe_1_7_0_U39 ( .A(npu_inst_pe_1_7_0_n79), .ZN(
        npu_inst_pe_1_7_0_n34) );
  AOI222_X1 npu_inst_pe_1_7_0_U38 ( .A1(1'b0), .A2(npu_inst_pe_1_7_0_n1), .B1(
        npu_inst_pe_1_7_0_N79), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N71), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n78) );
  INV_X1 npu_inst_pe_1_7_0_U37 ( .A(npu_inst_pe_1_7_0_n78), .ZN(
        npu_inst_pe_1_7_0_n33) );
  AOI222_X1 npu_inst_pe_1_7_0_U36 ( .A1(npu_inst_pe_1_7_0_n1), .A2(1'b0), .B1(
        npu_inst_pe_1_7_0_N80), .B2(npu_inst_pe_1_7_0_n76), .C1(
        npu_inst_pe_1_7_0_N72), .C2(npu_inst_pe_1_7_0_n77), .ZN(
        npu_inst_pe_1_7_0_n75) );
  INV_X1 npu_inst_pe_1_7_0_U35 ( .A(npu_inst_pe_1_7_0_n75), .ZN(
        npu_inst_pe_1_7_0_n32) );
  AND2_X1 npu_inst_pe_1_7_0_U34 ( .A1(npu_inst_pe_1_7_0_o_data_h_1_), .A2(
        npu_inst_pe_1_7_0_int_q_weight_1_), .ZN(npu_inst_pe_1_7_0_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_0_U33 ( .A1(npu_inst_pe_1_7_0_o_data_h_0_), .A2(
        npu_inst_pe_1_7_0_int_q_weight_1_), .ZN(npu_inst_pe_1_7_0_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_0_U32 ( .A(npu_inst_pe_1_7_0_int_data_1_), .ZN(
        npu_inst_pe_1_7_0_n13) );
  NOR3_X1 npu_inst_pe_1_7_0_U31 ( .A1(npu_inst_pe_1_7_0_n26), .A2(npu_inst_n35), .A3(npu_inst_int_ckg[7]), .ZN(npu_inst_pe_1_7_0_n85) );
  OR2_X1 npu_inst_pe_1_7_0_U30 ( .A1(npu_inst_pe_1_7_0_n85), .A2(
        npu_inst_pe_1_7_0_n1), .ZN(npu_inst_pe_1_7_0_N84) );
  INV_X1 npu_inst_pe_1_7_0_U29 ( .A(npu_inst_pe_1_7_0_int_data_0_), .ZN(
        npu_inst_pe_1_7_0_n12) );
  INV_X1 npu_inst_pe_1_7_0_U28 ( .A(npu_inst_n49), .ZN(npu_inst_pe_1_7_0_n4)
         );
  OR3_X1 npu_inst_pe_1_7_0_U27 ( .A1(npu_inst_pe_1_7_0_n5), .A2(
        npu_inst_pe_1_7_0_n7), .A3(npu_inst_pe_1_7_0_n4), .ZN(
        npu_inst_pe_1_7_0_n56) );
  OR3_X1 npu_inst_pe_1_7_0_U26 ( .A1(npu_inst_pe_1_7_0_n4), .A2(
        npu_inst_pe_1_7_0_n7), .A3(npu_inst_pe_1_7_0_n6), .ZN(
        npu_inst_pe_1_7_0_n48) );
  INV_X1 npu_inst_pe_1_7_0_U25 ( .A(npu_inst_pe_1_7_0_n4), .ZN(
        npu_inst_pe_1_7_0_n3) );
  OR3_X1 npu_inst_pe_1_7_0_U24 ( .A1(npu_inst_pe_1_7_0_n3), .A2(
        npu_inst_pe_1_7_0_n7), .A3(npu_inst_pe_1_7_0_n6), .ZN(
        npu_inst_pe_1_7_0_n52) );
  OR3_X1 npu_inst_pe_1_7_0_U23 ( .A1(npu_inst_pe_1_7_0_n5), .A2(
        npu_inst_pe_1_7_0_n7), .A3(npu_inst_pe_1_7_0_n3), .ZN(
        npu_inst_pe_1_7_0_n60) );
  BUF_X1 npu_inst_pe_1_7_0_U22 ( .A(npu_inst_n13), .Z(npu_inst_pe_1_7_0_n1) );
  NOR2_X1 npu_inst_pe_1_7_0_U21 ( .A1(npu_inst_pe_1_7_0_n60), .A2(
        npu_inst_pe_1_7_0_n2), .ZN(npu_inst_pe_1_7_0_n58) );
  NOR2_X1 npu_inst_pe_1_7_0_U20 ( .A1(npu_inst_pe_1_7_0_n56), .A2(
        npu_inst_pe_1_7_0_n2), .ZN(npu_inst_pe_1_7_0_n54) );
  NOR2_X1 npu_inst_pe_1_7_0_U19 ( .A1(npu_inst_pe_1_7_0_n52), .A2(
        npu_inst_pe_1_7_0_n2), .ZN(npu_inst_pe_1_7_0_n50) );
  NOR2_X1 npu_inst_pe_1_7_0_U18 ( .A1(npu_inst_pe_1_7_0_n48), .A2(
        npu_inst_pe_1_7_0_n2), .ZN(npu_inst_pe_1_7_0_n46) );
  NOR2_X1 npu_inst_pe_1_7_0_U17 ( .A1(npu_inst_pe_1_7_0_n40), .A2(
        npu_inst_pe_1_7_0_n2), .ZN(npu_inst_pe_1_7_0_n38) );
  NOR2_X1 npu_inst_pe_1_7_0_U16 ( .A1(npu_inst_pe_1_7_0_n44), .A2(
        npu_inst_pe_1_7_0_n2), .ZN(npu_inst_pe_1_7_0_n42) );
  BUF_X1 npu_inst_pe_1_7_0_U15 ( .A(npu_inst_n75), .Z(npu_inst_pe_1_7_0_n7) );
  INV_X1 npu_inst_pe_1_7_0_U14 ( .A(npu_inst_n104), .ZN(npu_inst_pe_1_7_0_n11)
         );
  INV_X1 npu_inst_pe_1_7_0_U13 ( .A(npu_inst_pe_1_7_0_n38), .ZN(
        npu_inst_pe_1_7_0_n113) );
  INV_X1 npu_inst_pe_1_7_0_U12 ( .A(npu_inst_pe_1_7_0_n58), .ZN(
        npu_inst_pe_1_7_0_n118) );
  INV_X1 npu_inst_pe_1_7_0_U11 ( .A(npu_inst_pe_1_7_0_n54), .ZN(
        npu_inst_pe_1_7_0_n117) );
  INV_X1 npu_inst_pe_1_7_0_U10 ( .A(npu_inst_pe_1_7_0_n50), .ZN(
        npu_inst_pe_1_7_0_n116) );
  INV_X1 npu_inst_pe_1_7_0_U9 ( .A(npu_inst_pe_1_7_0_n46), .ZN(
        npu_inst_pe_1_7_0_n115) );
  INV_X1 npu_inst_pe_1_7_0_U8 ( .A(npu_inst_pe_1_7_0_n42), .ZN(
        npu_inst_pe_1_7_0_n114) );
  BUF_X1 npu_inst_pe_1_7_0_U7 ( .A(npu_inst_pe_1_7_0_n11), .Z(
        npu_inst_pe_1_7_0_n10) );
  BUF_X1 npu_inst_pe_1_7_0_U6 ( .A(npu_inst_pe_1_7_0_n11), .Z(
        npu_inst_pe_1_7_0_n9) );
  BUF_X1 npu_inst_pe_1_7_0_U5 ( .A(npu_inst_pe_1_7_0_n11), .Z(
        npu_inst_pe_1_7_0_n8) );
  NOR2_X1 npu_inst_pe_1_7_0_U4 ( .A1(npu_inst_pe_1_7_0_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_0_n1), .ZN(npu_inst_pe_1_7_0_n76) );
  NOR2_X1 npu_inst_pe_1_7_0_U3 ( .A1(npu_inst_pe_1_7_0_n27), .A2(
        npu_inst_pe_1_7_0_n1), .ZN(npu_inst_pe_1_7_0_n77) );
  FA_X1 npu_inst_pe_1_7_0_sub_77_U2_1 ( .A(npu_inst_int_data_res_7__0__1_), 
        .B(npu_inst_pe_1_7_0_n13), .CI(npu_inst_pe_1_7_0_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_7_0_sub_77_carry_2_), .S(npu_inst_pe_1_7_0_N66) );
  FA_X1 npu_inst_pe_1_7_0_add_79_U1_1 ( .A(npu_inst_int_data_res_7__0__1_), 
        .B(npu_inst_pe_1_7_0_int_data_1_), .CI(
        npu_inst_pe_1_7_0_add_79_carry_1_), .CO(
        npu_inst_pe_1_7_0_add_79_carry_2_), .S(npu_inst_pe_1_7_0_N74) );
  NAND3_X1 npu_inst_pe_1_7_0_U101 ( .A1(npu_inst_pe_1_7_0_n4), .A2(
        npu_inst_pe_1_7_0_n6), .A3(npu_inst_pe_1_7_0_n7), .ZN(
        npu_inst_pe_1_7_0_n44) );
  NAND3_X1 npu_inst_pe_1_7_0_U100 ( .A1(npu_inst_pe_1_7_0_n3), .A2(
        npu_inst_pe_1_7_0_n6), .A3(npu_inst_pe_1_7_0_n7), .ZN(
        npu_inst_pe_1_7_0_n40) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_0_n33), .CK(
        npu_inst_pe_1_7_0_net3190), .RN(npu_inst_pe_1_7_0_n8), .Q(
        npu_inst_int_data_res_7__0__6_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_0_n34), .CK(
        npu_inst_pe_1_7_0_net3190), .RN(npu_inst_pe_1_7_0_n8), .Q(
        npu_inst_int_data_res_7__0__5_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_0_n35), .CK(
        npu_inst_pe_1_7_0_net3190), .RN(npu_inst_pe_1_7_0_n8), .Q(
        npu_inst_int_data_res_7__0__4_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_0_n36), .CK(
        npu_inst_pe_1_7_0_net3190), .RN(npu_inst_pe_1_7_0_n8), .Q(
        npu_inst_int_data_res_7__0__3_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_0_n98), .CK(
        npu_inst_pe_1_7_0_net3190), .RN(npu_inst_pe_1_7_0_n8), .Q(
        npu_inst_int_data_res_7__0__2_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_0_n99), .CK(
        npu_inst_pe_1_7_0_net3190), .RN(npu_inst_pe_1_7_0_n8), .Q(
        npu_inst_int_data_res_7__0__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_0_n32), .CK(
        npu_inst_pe_1_7_0_net3190), .RN(npu_inst_pe_1_7_0_n8), .Q(
        npu_inst_int_data_res_7__0__7_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_0_n100), 
        .CK(npu_inst_pe_1_7_0_net3190), .RN(npu_inst_pe_1_7_0_n8), .Q(
        npu_inst_int_data_res_7__0__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_weight_reg_0_ ( .D(npu_inst_n90), .CK(
        npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n8), .Q(
        npu_inst_pe_1_7_0_int_q_weight_0_), .QN(npu_inst_pe_1_7_0_n27) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_weight_reg_1_ ( .D(npu_inst_n96), .CK(
        npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n8), .Q(
        npu_inst_pe_1_7_0_int_q_weight_1_), .QN(npu_inst_pe_1_7_0_n26) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_0_n112), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n8), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_0_n111), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n8), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_0_n110), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_0_n109), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_0_n108), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_0_n107), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_0_n106), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_0_n105), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_0_n104), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_0_n103), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_0_n102), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_0_n101), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_0_n86), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_0_n87), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n9), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_0_n88), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_0_n89), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_0_n90), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_0_n91), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_0_n92), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_0_n93), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_0_n94), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_0_n95), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_0_n96), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_0_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_0_n97), 
        .CK(npu_inst_pe_1_7_0_net3196), .RN(npu_inst_pe_1_7_0_n10), .Q(
        npu_inst_pe_1_7_0_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_0_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_0_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_0_net3190) );
  CLKGATETST_X1 npu_inst_pe_1_7_0_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n43), .SE(1'b0), .GCK(npu_inst_pe_1_7_0_net3196) );
  MUX2_X1 npu_inst_pe_1_7_1_U153 ( .A(npu_inst_pe_1_7_1_n31), .B(
        npu_inst_pe_1_7_1_n28), .S(npu_inst_pe_1_7_1_n7), .Z(
        npu_inst_pe_1_7_1_N93) );
  MUX2_X1 npu_inst_pe_1_7_1_U152 ( .A(npu_inst_pe_1_7_1_n30), .B(
        npu_inst_pe_1_7_1_n29), .S(npu_inst_pe_1_7_1_n5), .Z(
        npu_inst_pe_1_7_1_n31) );
  MUX2_X1 npu_inst_pe_1_7_1_U151 ( .A(npu_inst_pe_1_7_1_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_1_n3), .Z(
        npu_inst_pe_1_7_1_n30) );
  MUX2_X1 npu_inst_pe_1_7_1_U150 ( .A(npu_inst_pe_1_7_1_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_1_n3), .Z(
        npu_inst_pe_1_7_1_n29) );
  MUX2_X1 npu_inst_pe_1_7_1_U149 ( .A(npu_inst_pe_1_7_1_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_1_n3), .Z(
        npu_inst_pe_1_7_1_n28) );
  MUX2_X1 npu_inst_pe_1_7_1_U148 ( .A(npu_inst_pe_1_7_1_n25), .B(
        npu_inst_pe_1_7_1_n22), .S(npu_inst_pe_1_7_1_n7), .Z(
        npu_inst_pe_1_7_1_N94) );
  MUX2_X1 npu_inst_pe_1_7_1_U147 ( .A(npu_inst_pe_1_7_1_n24), .B(
        npu_inst_pe_1_7_1_n23), .S(npu_inst_pe_1_7_1_n5), .Z(
        npu_inst_pe_1_7_1_n25) );
  MUX2_X1 npu_inst_pe_1_7_1_U146 ( .A(npu_inst_pe_1_7_1_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_1_n3), .Z(
        npu_inst_pe_1_7_1_n24) );
  MUX2_X1 npu_inst_pe_1_7_1_U145 ( .A(npu_inst_pe_1_7_1_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_1_n3), .Z(
        npu_inst_pe_1_7_1_n23) );
  MUX2_X1 npu_inst_pe_1_7_1_U144 ( .A(npu_inst_pe_1_7_1_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_1_n3), .Z(
        npu_inst_pe_1_7_1_n22) );
  MUX2_X1 npu_inst_pe_1_7_1_U143 ( .A(npu_inst_pe_1_7_1_n21), .B(
        npu_inst_pe_1_7_1_n18), .S(npu_inst_pe_1_7_1_n7), .Z(
        npu_inst_int_data_x_7__1__1_) );
  MUX2_X1 npu_inst_pe_1_7_1_U142 ( .A(npu_inst_pe_1_7_1_n20), .B(
        npu_inst_pe_1_7_1_n19), .S(npu_inst_pe_1_7_1_n5), .Z(
        npu_inst_pe_1_7_1_n21) );
  MUX2_X1 npu_inst_pe_1_7_1_U141 ( .A(npu_inst_pe_1_7_1_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_1_n3), .Z(
        npu_inst_pe_1_7_1_n20) );
  MUX2_X1 npu_inst_pe_1_7_1_U140 ( .A(npu_inst_pe_1_7_1_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_1_n3), .Z(
        npu_inst_pe_1_7_1_n19) );
  MUX2_X1 npu_inst_pe_1_7_1_U139 ( .A(npu_inst_pe_1_7_1_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_1_n3), .Z(
        npu_inst_pe_1_7_1_n18) );
  MUX2_X1 npu_inst_pe_1_7_1_U138 ( .A(npu_inst_pe_1_7_1_n17), .B(
        npu_inst_pe_1_7_1_n14), .S(npu_inst_pe_1_7_1_n7), .Z(
        npu_inst_int_data_x_7__1__0_) );
  MUX2_X1 npu_inst_pe_1_7_1_U137 ( .A(npu_inst_pe_1_7_1_n16), .B(
        npu_inst_pe_1_7_1_n15), .S(npu_inst_pe_1_7_1_n5), .Z(
        npu_inst_pe_1_7_1_n17) );
  MUX2_X1 npu_inst_pe_1_7_1_U136 ( .A(npu_inst_pe_1_7_1_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_1_n3), .Z(
        npu_inst_pe_1_7_1_n16) );
  MUX2_X1 npu_inst_pe_1_7_1_U135 ( .A(npu_inst_pe_1_7_1_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_1_n3), .Z(
        npu_inst_pe_1_7_1_n15) );
  MUX2_X1 npu_inst_pe_1_7_1_U134 ( .A(npu_inst_pe_1_7_1_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_1_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_1_n3), .Z(
        npu_inst_pe_1_7_1_n14) );
  XOR2_X1 npu_inst_pe_1_7_1_U133 ( .A(npu_inst_pe_1_7_1_int_data_0_), .B(
        npu_inst_int_data_res_7__1__0_), .Z(npu_inst_pe_1_7_1_N73) );
  AND2_X1 npu_inst_pe_1_7_1_U132 ( .A1(npu_inst_int_data_res_7__1__0_), .A2(
        npu_inst_pe_1_7_1_int_data_0_), .ZN(npu_inst_pe_1_7_1_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_1_U131 ( .A(npu_inst_int_data_res_7__1__0_), .B(
        npu_inst_pe_1_7_1_n12), .ZN(npu_inst_pe_1_7_1_N65) );
  OR2_X1 npu_inst_pe_1_7_1_U130 ( .A1(npu_inst_pe_1_7_1_n12), .A2(
        npu_inst_int_data_res_7__1__0_), .ZN(npu_inst_pe_1_7_1_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_1_U129 ( .A(npu_inst_int_data_res_7__1__2_), .B(
        npu_inst_pe_1_7_1_add_79_carry_2_), .Z(npu_inst_pe_1_7_1_N75) );
  AND2_X1 npu_inst_pe_1_7_1_U128 ( .A1(npu_inst_pe_1_7_1_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_7__1__2_), .ZN(
        npu_inst_pe_1_7_1_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_1_U127 ( .A(npu_inst_int_data_res_7__1__3_), .B(
        npu_inst_pe_1_7_1_add_79_carry_3_), .Z(npu_inst_pe_1_7_1_N76) );
  AND2_X1 npu_inst_pe_1_7_1_U126 ( .A1(npu_inst_pe_1_7_1_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_7__1__3_), .ZN(
        npu_inst_pe_1_7_1_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_1_U125 ( .A(npu_inst_int_data_res_7__1__4_), .B(
        npu_inst_pe_1_7_1_add_79_carry_4_), .Z(npu_inst_pe_1_7_1_N77) );
  AND2_X1 npu_inst_pe_1_7_1_U124 ( .A1(npu_inst_pe_1_7_1_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_7__1__4_), .ZN(
        npu_inst_pe_1_7_1_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_1_U123 ( .A(npu_inst_int_data_res_7__1__5_), .B(
        npu_inst_pe_1_7_1_add_79_carry_5_), .Z(npu_inst_pe_1_7_1_N78) );
  AND2_X1 npu_inst_pe_1_7_1_U122 ( .A1(npu_inst_pe_1_7_1_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_7__1__5_), .ZN(
        npu_inst_pe_1_7_1_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_1_U121 ( .A(npu_inst_int_data_res_7__1__6_), .B(
        npu_inst_pe_1_7_1_add_79_carry_6_), .Z(npu_inst_pe_1_7_1_N79) );
  AND2_X1 npu_inst_pe_1_7_1_U120 ( .A1(npu_inst_pe_1_7_1_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_7__1__6_), .ZN(
        npu_inst_pe_1_7_1_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_1_U119 ( .A(npu_inst_int_data_res_7__1__7_), .B(
        npu_inst_pe_1_7_1_add_79_carry_7_), .Z(npu_inst_pe_1_7_1_N80) );
  XNOR2_X1 npu_inst_pe_1_7_1_U118 ( .A(npu_inst_pe_1_7_1_sub_77_carry_2_), .B(
        npu_inst_int_data_res_7__1__2_), .ZN(npu_inst_pe_1_7_1_N67) );
  OR2_X1 npu_inst_pe_1_7_1_U117 ( .A1(npu_inst_int_data_res_7__1__2_), .A2(
        npu_inst_pe_1_7_1_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_7_1_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_1_U116 ( .A(npu_inst_pe_1_7_1_sub_77_carry_3_), .B(
        npu_inst_int_data_res_7__1__3_), .ZN(npu_inst_pe_1_7_1_N68) );
  OR2_X1 npu_inst_pe_1_7_1_U115 ( .A1(npu_inst_int_data_res_7__1__3_), .A2(
        npu_inst_pe_1_7_1_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_7_1_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_1_U114 ( .A(npu_inst_pe_1_7_1_sub_77_carry_4_), .B(
        npu_inst_int_data_res_7__1__4_), .ZN(npu_inst_pe_1_7_1_N69) );
  OR2_X1 npu_inst_pe_1_7_1_U113 ( .A1(npu_inst_int_data_res_7__1__4_), .A2(
        npu_inst_pe_1_7_1_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_7_1_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_1_U112 ( .A(npu_inst_pe_1_7_1_sub_77_carry_5_), .B(
        npu_inst_int_data_res_7__1__5_), .ZN(npu_inst_pe_1_7_1_N70) );
  OR2_X1 npu_inst_pe_1_7_1_U111 ( .A1(npu_inst_int_data_res_7__1__5_), .A2(
        npu_inst_pe_1_7_1_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_7_1_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_1_U110 ( .A(npu_inst_pe_1_7_1_sub_77_carry_6_), .B(
        npu_inst_int_data_res_7__1__6_), .ZN(npu_inst_pe_1_7_1_N71) );
  OR2_X1 npu_inst_pe_1_7_1_U109 ( .A1(npu_inst_int_data_res_7__1__6_), .A2(
        npu_inst_pe_1_7_1_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_7_1_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_1_U108 ( .A(npu_inst_int_data_res_7__1__7_), .B(
        npu_inst_pe_1_7_1_sub_77_carry_7_), .ZN(npu_inst_pe_1_7_1_N72) );
  INV_X1 npu_inst_pe_1_7_1_U107 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_7_1_n6)
         );
  INV_X1 npu_inst_pe_1_7_1_U106 ( .A(npu_inst_pe_1_7_1_n6), .ZN(
        npu_inst_pe_1_7_1_n5) );
  INV_X1 npu_inst_pe_1_7_1_U105 ( .A(npu_inst_n34), .ZN(npu_inst_pe_1_7_1_n2)
         );
  AOI22_X1 npu_inst_pe_1_7_1_U104 ( .A1(npu_inst_pe_1_7_1_n38), .A2(
        int_i_data_v_npu[13]), .B1(npu_inst_pe_1_7_1_n113), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_1_n39) );
  INV_X1 npu_inst_pe_1_7_1_U103 ( .A(npu_inst_pe_1_7_1_n39), .ZN(
        npu_inst_pe_1_7_1_n111) );
  AOI22_X1 npu_inst_pe_1_7_1_U102 ( .A1(npu_inst_pe_1_7_1_n38), .A2(
        int_i_data_v_npu[12]), .B1(npu_inst_pe_1_7_1_n113), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_1_n37) );
  INV_X1 npu_inst_pe_1_7_1_U99 ( .A(npu_inst_pe_1_7_1_n37), .ZN(
        npu_inst_pe_1_7_1_n112) );
  AOI22_X1 npu_inst_pe_1_7_1_U98 ( .A1(int_i_data_v_npu[13]), .A2(
        npu_inst_pe_1_7_1_n58), .B1(npu_inst_pe_1_7_1_n118), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_1_n59) );
  INV_X1 npu_inst_pe_1_7_1_U97 ( .A(npu_inst_pe_1_7_1_n59), .ZN(
        npu_inst_pe_1_7_1_n101) );
  AOI22_X1 npu_inst_pe_1_7_1_U96 ( .A1(int_i_data_v_npu[12]), .A2(
        npu_inst_pe_1_7_1_n58), .B1(npu_inst_pe_1_7_1_n118), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_1_n57) );
  INV_X1 npu_inst_pe_1_7_1_U95 ( .A(npu_inst_pe_1_7_1_n57), .ZN(
        npu_inst_pe_1_7_1_n102) );
  AOI22_X1 npu_inst_pe_1_7_1_U94 ( .A1(int_i_data_v_npu[13]), .A2(
        npu_inst_pe_1_7_1_n54), .B1(npu_inst_pe_1_7_1_n117), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_1_n55) );
  INV_X1 npu_inst_pe_1_7_1_U93 ( .A(npu_inst_pe_1_7_1_n55), .ZN(
        npu_inst_pe_1_7_1_n103) );
  AOI22_X1 npu_inst_pe_1_7_1_U92 ( .A1(int_i_data_v_npu[12]), .A2(
        npu_inst_pe_1_7_1_n54), .B1(npu_inst_pe_1_7_1_n117), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_1_n53) );
  INV_X1 npu_inst_pe_1_7_1_U91 ( .A(npu_inst_pe_1_7_1_n53), .ZN(
        npu_inst_pe_1_7_1_n104) );
  AOI22_X1 npu_inst_pe_1_7_1_U90 ( .A1(int_i_data_v_npu[13]), .A2(
        npu_inst_pe_1_7_1_n50), .B1(npu_inst_pe_1_7_1_n116), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_1_n51) );
  INV_X1 npu_inst_pe_1_7_1_U89 ( .A(npu_inst_pe_1_7_1_n51), .ZN(
        npu_inst_pe_1_7_1_n105) );
  AOI22_X1 npu_inst_pe_1_7_1_U88 ( .A1(int_i_data_v_npu[12]), .A2(
        npu_inst_pe_1_7_1_n50), .B1(npu_inst_pe_1_7_1_n116), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_1_n49) );
  INV_X1 npu_inst_pe_1_7_1_U87 ( .A(npu_inst_pe_1_7_1_n49), .ZN(
        npu_inst_pe_1_7_1_n106) );
  AOI22_X1 npu_inst_pe_1_7_1_U86 ( .A1(int_i_data_v_npu[13]), .A2(
        npu_inst_pe_1_7_1_n46), .B1(npu_inst_pe_1_7_1_n115), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_1_n47) );
  INV_X1 npu_inst_pe_1_7_1_U85 ( .A(npu_inst_pe_1_7_1_n47), .ZN(
        npu_inst_pe_1_7_1_n107) );
  AOI22_X1 npu_inst_pe_1_7_1_U84 ( .A1(int_i_data_v_npu[12]), .A2(
        npu_inst_pe_1_7_1_n46), .B1(npu_inst_pe_1_7_1_n115), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_1_n45) );
  INV_X1 npu_inst_pe_1_7_1_U83 ( .A(npu_inst_pe_1_7_1_n45), .ZN(
        npu_inst_pe_1_7_1_n108) );
  AOI22_X1 npu_inst_pe_1_7_1_U82 ( .A1(int_i_data_v_npu[13]), .A2(
        npu_inst_pe_1_7_1_n42), .B1(npu_inst_pe_1_7_1_n114), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_1_n43) );
  INV_X1 npu_inst_pe_1_7_1_U81 ( .A(npu_inst_pe_1_7_1_n43), .ZN(
        npu_inst_pe_1_7_1_n109) );
  AOI22_X1 npu_inst_pe_1_7_1_U80 ( .A1(int_i_data_v_npu[12]), .A2(
        npu_inst_pe_1_7_1_n42), .B1(npu_inst_pe_1_7_1_n114), .B2(
        npu_inst_pe_1_7_1_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_1_n41) );
  INV_X1 npu_inst_pe_1_7_1_U79 ( .A(npu_inst_pe_1_7_1_n41), .ZN(
        npu_inst_pe_1_7_1_n110) );
  AND2_X1 npu_inst_pe_1_7_1_U78 ( .A1(npu_inst_pe_1_7_1_N93), .A2(npu_inst_n34), .ZN(npu_inst_int_data_y_7__1__0_) );
  NAND2_X1 npu_inst_pe_1_7_1_U77 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_1_n60), .ZN(npu_inst_pe_1_7_1_n74) );
  OAI21_X1 npu_inst_pe_1_7_1_U76 ( .B1(npu_inst_pe_1_7_1_n63), .B2(
        npu_inst_pe_1_7_1_n60), .A(npu_inst_pe_1_7_1_n74), .ZN(
        npu_inst_pe_1_7_1_n97) );
  NAND2_X1 npu_inst_pe_1_7_1_U75 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_1_n60), .ZN(npu_inst_pe_1_7_1_n73) );
  OAI21_X1 npu_inst_pe_1_7_1_U74 ( .B1(npu_inst_pe_1_7_1_n61), .B2(
        npu_inst_pe_1_7_1_n60), .A(npu_inst_pe_1_7_1_n73), .ZN(
        npu_inst_pe_1_7_1_n96) );
  NAND2_X1 npu_inst_pe_1_7_1_U73 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_1_n56), .ZN(npu_inst_pe_1_7_1_n72) );
  OAI21_X1 npu_inst_pe_1_7_1_U72 ( .B1(npu_inst_pe_1_7_1_n63), .B2(
        npu_inst_pe_1_7_1_n56), .A(npu_inst_pe_1_7_1_n72), .ZN(
        npu_inst_pe_1_7_1_n95) );
  NAND2_X1 npu_inst_pe_1_7_1_U71 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_1_n56), .ZN(npu_inst_pe_1_7_1_n71) );
  OAI21_X1 npu_inst_pe_1_7_1_U70 ( .B1(npu_inst_pe_1_7_1_n61), .B2(
        npu_inst_pe_1_7_1_n56), .A(npu_inst_pe_1_7_1_n71), .ZN(
        npu_inst_pe_1_7_1_n94) );
  NAND2_X1 npu_inst_pe_1_7_1_U69 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_1_n52), .ZN(npu_inst_pe_1_7_1_n70) );
  OAI21_X1 npu_inst_pe_1_7_1_U68 ( .B1(npu_inst_pe_1_7_1_n63), .B2(
        npu_inst_pe_1_7_1_n52), .A(npu_inst_pe_1_7_1_n70), .ZN(
        npu_inst_pe_1_7_1_n93) );
  NAND2_X1 npu_inst_pe_1_7_1_U67 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_1_n52), .ZN(npu_inst_pe_1_7_1_n69) );
  OAI21_X1 npu_inst_pe_1_7_1_U66 ( .B1(npu_inst_pe_1_7_1_n61), .B2(
        npu_inst_pe_1_7_1_n52), .A(npu_inst_pe_1_7_1_n69), .ZN(
        npu_inst_pe_1_7_1_n92) );
  NAND2_X1 npu_inst_pe_1_7_1_U65 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_1_n48), .ZN(npu_inst_pe_1_7_1_n68) );
  OAI21_X1 npu_inst_pe_1_7_1_U64 ( .B1(npu_inst_pe_1_7_1_n63), .B2(
        npu_inst_pe_1_7_1_n48), .A(npu_inst_pe_1_7_1_n68), .ZN(
        npu_inst_pe_1_7_1_n91) );
  NAND2_X1 npu_inst_pe_1_7_1_U63 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_1_n48), .ZN(npu_inst_pe_1_7_1_n67) );
  OAI21_X1 npu_inst_pe_1_7_1_U62 ( .B1(npu_inst_pe_1_7_1_n61), .B2(
        npu_inst_pe_1_7_1_n48), .A(npu_inst_pe_1_7_1_n67), .ZN(
        npu_inst_pe_1_7_1_n90) );
  NAND2_X1 npu_inst_pe_1_7_1_U61 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_1_n44), .ZN(npu_inst_pe_1_7_1_n66) );
  OAI21_X1 npu_inst_pe_1_7_1_U60 ( .B1(npu_inst_pe_1_7_1_n63), .B2(
        npu_inst_pe_1_7_1_n44), .A(npu_inst_pe_1_7_1_n66), .ZN(
        npu_inst_pe_1_7_1_n89) );
  NAND2_X1 npu_inst_pe_1_7_1_U59 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_1_n44), .ZN(npu_inst_pe_1_7_1_n65) );
  OAI21_X1 npu_inst_pe_1_7_1_U58 ( .B1(npu_inst_pe_1_7_1_n61), .B2(
        npu_inst_pe_1_7_1_n44), .A(npu_inst_pe_1_7_1_n65), .ZN(
        npu_inst_pe_1_7_1_n88) );
  NAND2_X1 npu_inst_pe_1_7_1_U57 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_1_n40), .ZN(npu_inst_pe_1_7_1_n64) );
  OAI21_X1 npu_inst_pe_1_7_1_U56 ( .B1(npu_inst_pe_1_7_1_n63), .B2(
        npu_inst_pe_1_7_1_n40), .A(npu_inst_pe_1_7_1_n64), .ZN(
        npu_inst_pe_1_7_1_n87) );
  NAND2_X1 npu_inst_pe_1_7_1_U55 ( .A1(npu_inst_pe_1_7_1_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_1_n40), .ZN(npu_inst_pe_1_7_1_n62) );
  OAI21_X1 npu_inst_pe_1_7_1_U54 ( .B1(npu_inst_pe_1_7_1_n61), .B2(
        npu_inst_pe_1_7_1_n40), .A(npu_inst_pe_1_7_1_n62), .ZN(
        npu_inst_pe_1_7_1_n86) );
  AND2_X1 npu_inst_pe_1_7_1_U53 ( .A1(npu_inst_n34), .A2(npu_inst_pe_1_7_1_N94), .ZN(npu_inst_int_data_y_7__1__1_) );
  AOI22_X1 npu_inst_pe_1_7_1_U52 ( .A1(npu_inst_n34), .A2(int_i_data_v_npu[13]), .B1(npu_inst_pe_1_7_1_n2), .B2(npu_inst_int_data_x_7__2__1_), .ZN(
        npu_inst_pe_1_7_1_n63) );
  AOI22_X1 npu_inst_pe_1_7_1_U51 ( .A1(npu_inst_n34), .A2(int_i_data_v_npu[12]), .B1(npu_inst_pe_1_7_1_n2), .B2(npu_inst_int_data_x_7__2__0_), .ZN(
        npu_inst_pe_1_7_1_n61) );
  AOI222_X1 npu_inst_pe_1_7_1_U50 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N73), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N65), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n84) );
  INV_X1 npu_inst_pe_1_7_1_U49 ( .A(npu_inst_pe_1_7_1_n84), .ZN(
        npu_inst_pe_1_7_1_n100) );
  AOI222_X1 npu_inst_pe_1_7_1_U48 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N74), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N66), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n83) );
  INV_X1 npu_inst_pe_1_7_1_U47 ( .A(npu_inst_pe_1_7_1_n83), .ZN(
        npu_inst_pe_1_7_1_n99) );
  AOI222_X1 npu_inst_pe_1_7_1_U46 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N75), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N67), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n82) );
  INV_X1 npu_inst_pe_1_7_1_U45 ( .A(npu_inst_pe_1_7_1_n82), .ZN(
        npu_inst_pe_1_7_1_n98) );
  AOI222_X1 npu_inst_pe_1_7_1_U44 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N76), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N68), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n81) );
  INV_X1 npu_inst_pe_1_7_1_U43 ( .A(npu_inst_pe_1_7_1_n81), .ZN(
        npu_inst_pe_1_7_1_n36) );
  AOI222_X1 npu_inst_pe_1_7_1_U42 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N77), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N69), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n80) );
  INV_X1 npu_inst_pe_1_7_1_U41 ( .A(npu_inst_pe_1_7_1_n80), .ZN(
        npu_inst_pe_1_7_1_n35) );
  AOI222_X1 npu_inst_pe_1_7_1_U40 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N78), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N70), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n79) );
  INV_X1 npu_inst_pe_1_7_1_U39 ( .A(npu_inst_pe_1_7_1_n79), .ZN(
        npu_inst_pe_1_7_1_n34) );
  AOI222_X1 npu_inst_pe_1_7_1_U38 ( .A1(1'b0), .A2(npu_inst_pe_1_7_1_n1), .B1(
        npu_inst_pe_1_7_1_N79), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N71), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n78) );
  INV_X1 npu_inst_pe_1_7_1_U37 ( .A(npu_inst_pe_1_7_1_n78), .ZN(
        npu_inst_pe_1_7_1_n33) );
  AOI222_X1 npu_inst_pe_1_7_1_U36 ( .A1(npu_inst_pe_1_7_1_n1), .A2(1'b0), .B1(
        npu_inst_pe_1_7_1_N80), .B2(npu_inst_pe_1_7_1_n76), .C1(
        npu_inst_pe_1_7_1_N72), .C2(npu_inst_pe_1_7_1_n77), .ZN(
        npu_inst_pe_1_7_1_n75) );
  INV_X1 npu_inst_pe_1_7_1_U35 ( .A(npu_inst_pe_1_7_1_n75), .ZN(
        npu_inst_pe_1_7_1_n32) );
  AND2_X1 npu_inst_pe_1_7_1_U34 ( .A1(npu_inst_int_data_x_7__1__1_), .A2(
        npu_inst_pe_1_7_1_int_q_weight_1_), .ZN(npu_inst_pe_1_7_1_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_1_U33 ( .A1(npu_inst_int_data_x_7__1__0_), .A2(
        npu_inst_pe_1_7_1_int_q_weight_1_), .ZN(npu_inst_pe_1_7_1_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_1_U32 ( .A(npu_inst_pe_1_7_1_int_data_1_), .ZN(
        npu_inst_pe_1_7_1_n13) );
  NOR3_X1 npu_inst_pe_1_7_1_U31 ( .A1(npu_inst_pe_1_7_1_n26), .A2(npu_inst_n34), .A3(npu_inst_int_ckg[6]), .ZN(npu_inst_pe_1_7_1_n85) );
  OR2_X1 npu_inst_pe_1_7_1_U30 ( .A1(npu_inst_pe_1_7_1_n85), .A2(
        npu_inst_pe_1_7_1_n1), .ZN(npu_inst_pe_1_7_1_N84) );
  INV_X1 npu_inst_pe_1_7_1_U29 ( .A(npu_inst_pe_1_7_1_int_data_0_), .ZN(
        npu_inst_pe_1_7_1_n12) );
  INV_X1 npu_inst_pe_1_7_1_U28 ( .A(npu_inst_n49), .ZN(npu_inst_pe_1_7_1_n4)
         );
  OR3_X1 npu_inst_pe_1_7_1_U27 ( .A1(npu_inst_pe_1_7_1_n5), .A2(
        npu_inst_pe_1_7_1_n7), .A3(npu_inst_pe_1_7_1_n4), .ZN(
        npu_inst_pe_1_7_1_n56) );
  OR3_X1 npu_inst_pe_1_7_1_U26 ( .A1(npu_inst_pe_1_7_1_n4), .A2(
        npu_inst_pe_1_7_1_n7), .A3(npu_inst_pe_1_7_1_n6), .ZN(
        npu_inst_pe_1_7_1_n48) );
  INV_X1 npu_inst_pe_1_7_1_U25 ( .A(npu_inst_pe_1_7_1_n4), .ZN(
        npu_inst_pe_1_7_1_n3) );
  OR3_X1 npu_inst_pe_1_7_1_U24 ( .A1(npu_inst_pe_1_7_1_n3), .A2(
        npu_inst_pe_1_7_1_n7), .A3(npu_inst_pe_1_7_1_n6), .ZN(
        npu_inst_pe_1_7_1_n52) );
  OR3_X1 npu_inst_pe_1_7_1_U23 ( .A1(npu_inst_pe_1_7_1_n5), .A2(
        npu_inst_pe_1_7_1_n7), .A3(npu_inst_pe_1_7_1_n3), .ZN(
        npu_inst_pe_1_7_1_n60) );
  BUF_X1 npu_inst_pe_1_7_1_U22 ( .A(npu_inst_n13), .Z(npu_inst_pe_1_7_1_n1) );
  NOR2_X1 npu_inst_pe_1_7_1_U21 ( .A1(npu_inst_pe_1_7_1_n60), .A2(
        npu_inst_pe_1_7_1_n2), .ZN(npu_inst_pe_1_7_1_n58) );
  NOR2_X1 npu_inst_pe_1_7_1_U20 ( .A1(npu_inst_pe_1_7_1_n56), .A2(
        npu_inst_pe_1_7_1_n2), .ZN(npu_inst_pe_1_7_1_n54) );
  NOR2_X1 npu_inst_pe_1_7_1_U19 ( .A1(npu_inst_pe_1_7_1_n52), .A2(
        npu_inst_pe_1_7_1_n2), .ZN(npu_inst_pe_1_7_1_n50) );
  NOR2_X1 npu_inst_pe_1_7_1_U18 ( .A1(npu_inst_pe_1_7_1_n48), .A2(
        npu_inst_pe_1_7_1_n2), .ZN(npu_inst_pe_1_7_1_n46) );
  NOR2_X1 npu_inst_pe_1_7_1_U17 ( .A1(npu_inst_pe_1_7_1_n40), .A2(
        npu_inst_pe_1_7_1_n2), .ZN(npu_inst_pe_1_7_1_n38) );
  NOR2_X1 npu_inst_pe_1_7_1_U16 ( .A1(npu_inst_pe_1_7_1_n44), .A2(
        npu_inst_pe_1_7_1_n2), .ZN(npu_inst_pe_1_7_1_n42) );
  BUF_X1 npu_inst_pe_1_7_1_U15 ( .A(npu_inst_n75), .Z(npu_inst_pe_1_7_1_n7) );
  INV_X1 npu_inst_pe_1_7_1_U14 ( .A(npu_inst_n104), .ZN(npu_inst_pe_1_7_1_n11)
         );
  INV_X1 npu_inst_pe_1_7_1_U13 ( .A(npu_inst_pe_1_7_1_n38), .ZN(
        npu_inst_pe_1_7_1_n113) );
  INV_X1 npu_inst_pe_1_7_1_U12 ( .A(npu_inst_pe_1_7_1_n58), .ZN(
        npu_inst_pe_1_7_1_n118) );
  INV_X1 npu_inst_pe_1_7_1_U11 ( .A(npu_inst_pe_1_7_1_n54), .ZN(
        npu_inst_pe_1_7_1_n117) );
  INV_X1 npu_inst_pe_1_7_1_U10 ( .A(npu_inst_pe_1_7_1_n50), .ZN(
        npu_inst_pe_1_7_1_n116) );
  INV_X1 npu_inst_pe_1_7_1_U9 ( .A(npu_inst_pe_1_7_1_n46), .ZN(
        npu_inst_pe_1_7_1_n115) );
  INV_X1 npu_inst_pe_1_7_1_U8 ( .A(npu_inst_pe_1_7_1_n42), .ZN(
        npu_inst_pe_1_7_1_n114) );
  BUF_X1 npu_inst_pe_1_7_1_U7 ( .A(npu_inst_pe_1_7_1_n11), .Z(
        npu_inst_pe_1_7_1_n10) );
  BUF_X1 npu_inst_pe_1_7_1_U6 ( .A(npu_inst_pe_1_7_1_n11), .Z(
        npu_inst_pe_1_7_1_n9) );
  BUF_X1 npu_inst_pe_1_7_1_U5 ( .A(npu_inst_pe_1_7_1_n11), .Z(
        npu_inst_pe_1_7_1_n8) );
  NOR2_X1 npu_inst_pe_1_7_1_U4 ( .A1(npu_inst_pe_1_7_1_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_1_n1), .ZN(npu_inst_pe_1_7_1_n76) );
  NOR2_X1 npu_inst_pe_1_7_1_U3 ( .A1(npu_inst_pe_1_7_1_n27), .A2(
        npu_inst_pe_1_7_1_n1), .ZN(npu_inst_pe_1_7_1_n77) );
  FA_X1 npu_inst_pe_1_7_1_sub_77_U2_1 ( .A(npu_inst_int_data_res_7__1__1_), 
        .B(npu_inst_pe_1_7_1_n13), .CI(npu_inst_pe_1_7_1_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_7_1_sub_77_carry_2_), .S(npu_inst_pe_1_7_1_N66) );
  FA_X1 npu_inst_pe_1_7_1_add_79_U1_1 ( .A(npu_inst_int_data_res_7__1__1_), 
        .B(npu_inst_pe_1_7_1_int_data_1_), .CI(
        npu_inst_pe_1_7_1_add_79_carry_1_), .CO(
        npu_inst_pe_1_7_1_add_79_carry_2_), .S(npu_inst_pe_1_7_1_N74) );
  NAND3_X1 npu_inst_pe_1_7_1_U101 ( .A1(npu_inst_pe_1_7_1_n4), .A2(
        npu_inst_pe_1_7_1_n6), .A3(npu_inst_pe_1_7_1_n7), .ZN(
        npu_inst_pe_1_7_1_n44) );
  NAND3_X1 npu_inst_pe_1_7_1_U100 ( .A1(npu_inst_pe_1_7_1_n3), .A2(
        npu_inst_pe_1_7_1_n6), .A3(npu_inst_pe_1_7_1_n7), .ZN(
        npu_inst_pe_1_7_1_n40) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_1_n33), .CK(
        npu_inst_pe_1_7_1_net3167), .RN(npu_inst_pe_1_7_1_n8), .Q(
        npu_inst_int_data_res_7__1__6_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_1_n34), .CK(
        npu_inst_pe_1_7_1_net3167), .RN(npu_inst_pe_1_7_1_n8), .Q(
        npu_inst_int_data_res_7__1__5_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_1_n35), .CK(
        npu_inst_pe_1_7_1_net3167), .RN(npu_inst_pe_1_7_1_n8), .Q(
        npu_inst_int_data_res_7__1__4_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_1_n36), .CK(
        npu_inst_pe_1_7_1_net3167), .RN(npu_inst_pe_1_7_1_n8), .Q(
        npu_inst_int_data_res_7__1__3_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_1_n98), .CK(
        npu_inst_pe_1_7_1_net3167), .RN(npu_inst_pe_1_7_1_n8), .Q(
        npu_inst_int_data_res_7__1__2_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_1_n99), .CK(
        npu_inst_pe_1_7_1_net3167), .RN(npu_inst_pe_1_7_1_n8), .Q(
        npu_inst_int_data_res_7__1__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_1_n32), .CK(
        npu_inst_pe_1_7_1_net3167), .RN(npu_inst_pe_1_7_1_n8), .Q(
        npu_inst_int_data_res_7__1__7_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_1_n100), 
        .CK(npu_inst_pe_1_7_1_net3167), .RN(npu_inst_pe_1_7_1_n8), .Q(
        npu_inst_int_data_res_7__1__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_weight_reg_0_ ( .D(npu_inst_n90), .CK(
        npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n8), .Q(
        npu_inst_pe_1_7_1_int_q_weight_0_), .QN(npu_inst_pe_1_7_1_n27) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_weight_reg_1_ ( .D(npu_inst_n96), .CK(
        npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n8), .Q(
        npu_inst_pe_1_7_1_int_q_weight_1_), .QN(npu_inst_pe_1_7_1_n26) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_1_n112), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n8), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_1_n111), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n8), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_1_n110), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_1_n109), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_1_n108), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_1_n107), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_1_n106), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_1_n105), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_1_n104), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_1_n103), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_1_n102), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_1_n101), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_1_n86), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_1_n87), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n9), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_1_n88), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_1_n89), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_1_n90), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_1_n91), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_1_n92), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_1_n93), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_1_n94), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_1_n95), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_1_n96), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_1_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_1_n97), 
        .CK(npu_inst_pe_1_7_1_net3173), .RN(npu_inst_pe_1_7_1_n10), .Q(
        npu_inst_pe_1_7_1_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_1_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_1_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_1_net3167) );
  CLKGATETST_X1 npu_inst_pe_1_7_1_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n43), .SE(1'b0), .GCK(npu_inst_pe_1_7_1_net3173) );
  MUX2_X1 npu_inst_pe_1_7_2_U153 ( .A(npu_inst_pe_1_7_2_n31), .B(
        npu_inst_pe_1_7_2_n28), .S(npu_inst_pe_1_7_2_n7), .Z(
        npu_inst_pe_1_7_2_N93) );
  MUX2_X1 npu_inst_pe_1_7_2_U152 ( .A(npu_inst_pe_1_7_2_n30), .B(
        npu_inst_pe_1_7_2_n29), .S(npu_inst_pe_1_7_2_n5), .Z(
        npu_inst_pe_1_7_2_n31) );
  MUX2_X1 npu_inst_pe_1_7_2_U151 ( .A(npu_inst_pe_1_7_2_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_2_n3), .Z(
        npu_inst_pe_1_7_2_n30) );
  MUX2_X1 npu_inst_pe_1_7_2_U150 ( .A(npu_inst_pe_1_7_2_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_2_n3), .Z(
        npu_inst_pe_1_7_2_n29) );
  MUX2_X1 npu_inst_pe_1_7_2_U149 ( .A(npu_inst_pe_1_7_2_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_2_n3), .Z(
        npu_inst_pe_1_7_2_n28) );
  MUX2_X1 npu_inst_pe_1_7_2_U148 ( .A(npu_inst_pe_1_7_2_n25), .B(
        npu_inst_pe_1_7_2_n22), .S(npu_inst_pe_1_7_2_n7), .Z(
        npu_inst_pe_1_7_2_N94) );
  MUX2_X1 npu_inst_pe_1_7_2_U147 ( .A(npu_inst_pe_1_7_2_n24), .B(
        npu_inst_pe_1_7_2_n23), .S(npu_inst_pe_1_7_2_n5), .Z(
        npu_inst_pe_1_7_2_n25) );
  MUX2_X1 npu_inst_pe_1_7_2_U146 ( .A(npu_inst_pe_1_7_2_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_2_n3), .Z(
        npu_inst_pe_1_7_2_n24) );
  MUX2_X1 npu_inst_pe_1_7_2_U145 ( .A(npu_inst_pe_1_7_2_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_2_n3), .Z(
        npu_inst_pe_1_7_2_n23) );
  MUX2_X1 npu_inst_pe_1_7_2_U144 ( .A(npu_inst_pe_1_7_2_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_2_n3), .Z(
        npu_inst_pe_1_7_2_n22) );
  MUX2_X1 npu_inst_pe_1_7_2_U143 ( .A(npu_inst_pe_1_7_2_n21), .B(
        npu_inst_pe_1_7_2_n18), .S(npu_inst_pe_1_7_2_n7), .Z(
        npu_inst_int_data_x_7__2__1_) );
  MUX2_X1 npu_inst_pe_1_7_2_U142 ( .A(npu_inst_pe_1_7_2_n20), .B(
        npu_inst_pe_1_7_2_n19), .S(npu_inst_pe_1_7_2_n5), .Z(
        npu_inst_pe_1_7_2_n21) );
  MUX2_X1 npu_inst_pe_1_7_2_U141 ( .A(npu_inst_pe_1_7_2_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_2_n3), .Z(
        npu_inst_pe_1_7_2_n20) );
  MUX2_X1 npu_inst_pe_1_7_2_U140 ( .A(npu_inst_pe_1_7_2_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_2_n3), .Z(
        npu_inst_pe_1_7_2_n19) );
  MUX2_X1 npu_inst_pe_1_7_2_U139 ( .A(npu_inst_pe_1_7_2_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_2_n3), .Z(
        npu_inst_pe_1_7_2_n18) );
  MUX2_X1 npu_inst_pe_1_7_2_U138 ( .A(npu_inst_pe_1_7_2_n17), .B(
        npu_inst_pe_1_7_2_n14), .S(npu_inst_pe_1_7_2_n7), .Z(
        npu_inst_int_data_x_7__2__0_) );
  MUX2_X1 npu_inst_pe_1_7_2_U137 ( .A(npu_inst_pe_1_7_2_n16), .B(
        npu_inst_pe_1_7_2_n15), .S(npu_inst_pe_1_7_2_n5), .Z(
        npu_inst_pe_1_7_2_n17) );
  MUX2_X1 npu_inst_pe_1_7_2_U136 ( .A(npu_inst_pe_1_7_2_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_2_n3), .Z(
        npu_inst_pe_1_7_2_n16) );
  MUX2_X1 npu_inst_pe_1_7_2_U135 ( .A(npu_inst_pe_1_7_2_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_2_n3), .Z(
        npu_inst_pe_1_7_2_n15) );
  MUX2_X1 npu_inst_pe_1_7_2_U134 ( .A(npu_inst_pe_1_7_2_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_2_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_2_n3), .Z(
        npu_inst_pe_1_7_2_n14) );
  XOR2_X1 npu_inst_pe_1_7_2_U133 ( .A(npu_inst_pe_1_7_2_int_data_0_), .B(
        npu_inst_int_data_res_7__2__0_), .Z(npu_inst_pe_1_7_2_N73) );
  AND2_X1 npu_inst_pe_1_7_2_U132 ( .A1(npu_inst_int_data_res_7__2__0_), .A2(
        npu_inst_pe_1_7_2_int_data_0_), .ZN(npu_inst_pe_1_7_2_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_2_U131 ( .A(npu_inst_int_data_res_7__2__0_), .B(
        npu_inst_pe_1_7_2_n12), .ZN(npu_inst_pe_1_7_2_N65) );
  OR2_X1 npu_inst_pe_1_7_2_U130 ( .A1(npu_inst_pe_1_7_2_n12), .A2(
        npu_inst_int_data_res_7__2__0_), .ZN(npu_inst_pe_1_7_2_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_2_U129 ( .A(npu_inst_int_data_res_7__2__2_), .B(
        npu_inst_pe_1_7_2_add_79_carry_2_), .Z(npu_inst_pe_1_7_2_N75) );
  AND2_X1 npu_inst_pe_1_7_2_U128 ( .A1(npu_inst_pe_1_7_2_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_7__2__2_), .ZN(
        npu_inst_pe_1_7_2_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_2_U127 ( .A(npu_inst_int_data_res_7__2__3_), .B(
        npu_inst_pe_1_7_2_add_79_carry_3_), .Z(npu_inst_pe_1_7_2_N76) );
  AND2_X1 npu_inst_pe_1_7_2_U126 ( .A1(npu_inst_pe_1_7_2_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_7__2__3_), .ZN(
        npu_inst_pe_1_7_2_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_2_U125 ( .A(npu_inst_int_data_res_7__2__4_), .B(
        npu_inst_pe_1_7_2_add_79_carry_4_), .Z(npu_inst_pe_1_7_2_N77) );
  AND2_X1 npu_inst_pe_1_7_2_U124 ( .A1(npu_inst_pe_1_7_2_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_7__2__4_), .ZN(
        npu_inst_pe_1_7_2_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_2_U123 ( .A(npu_inst_int_data_res_7__2__5_), .B(
        npu_inst_pe_1_7_2_add_79_carry_5_), .Z(npu_inst_pe_1_7_2_N78) );
  AND2_X1 npu_inst_pe_1_7_2_U122 ( .A1(npu_inst_pe_1_7_2_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_7__2__5_), .ZN(
        npu_inst_pe_1_7_2_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_2_U121 ( .A(npu_inst_int_data_res_7__2__6_), .B(
        npu_inst_pe_1_7_2_add_79_carry_6_), .Z(npu_inst_pe_1_7_2_N79) );
  AND2_X1 npu_inst_pe_1_7_2_U120 ( .A1(npu_inst_pe_1_7_2_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_7__2__6_), .ZN(
        npu_inst_pe_1_7_2_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_2_U119 ( .A(npu_inst_int_data_res_7__2__7_), .B(
        npu_inst_pe_1_7_2_add_79_carry_7_), .Z(npu_inst_pe_1_7_2_N80) );
  XNOR2_X1 npu_inst_pe_1_7_2_U118 ( .A(npu_inst_pe_1_7_2_sub_77_carry_2_), .B(
        npu_inst_int_data_res_7__2__2_), .ZN(npu_inst_pe_1_7_2_N67) );
  OR2_X1 npu_inst_pe_1_7_2_U117 ( .A1(npu_inst_int_data_res_7__2__2_), .A2(
        npu_inst_pe_1_7_2_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_7_2_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_2_U116 ( .A(npu_inst_pe_1_7_2_sub_77_carry_3_), .B(
        npu_inst_int_data_res_7__2__3_), .ZN(npu_inst_pe_1_7_2_N68) );
  OR2_X1 npu_inst_pe_1_7_2_U115 ( .A1(npu_inst_int_data_res_7__2__3_), .A2(
        npu_inst_pe_1_7_2_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_7_2_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_2_U114 ( .A(npu_inst_pe_1_7_2_sub_77_carry_4_), .B(
        npu_inst_int_data_res_7__2__4_), .ZN(npu_inst_pe_1_7_2_N69) );
  OR2_X1 npu_inst_pe_1_7_2_U113 ( .A1(npu_inst_int_data_res_7__2__4_), .A2(
        npu_inst_pe_1_7_2_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_7_2_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_2_U112 ( .A(npu_inst_pe_1_7_2_sub_77_carry_5_), .B(
        npu_inst_int_data_res_7__2__5_), .ZN(npu_inst_pe_1_7_2_N70) );
  OR2_X1 npu_inst_pe_1_7_2_U111 ( .A1(npu_inst_int_data_res_7__2__5_), .A2(
        npu_inst_pe_1_7_2_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_7_2_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_2_U110 ( .A(npu_inst_pe_1_7_2_sub_77_carry_6_), .B(
        npu_inst_int_data_res_7__2__6_), .ZN(npu_inst_pe_1_7_2_N71) );
  OR2_X1 npu_inst_pe_1_7_2_U109 ( .A1(npu_inst_int_data_res_7__2__6_), .A2(
        npu_inst_pe_1_7_2_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_7_2_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_2_U108 ( .A(npu_inst_int_data_res_7__2__7_), .B(
        npu_inst_pe_1_7_2_sub_77_carry_7_), .ZN(npu_inst_pe_1_7_2_N72) );
  INV_X1 npu_inst_pe_1_7_2_U107 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_7_2_n6)
         );
  INV_X1 npu_inst_pe_1_7_2_U106 ( .A(npu_inst_pe_1_7_2_n6), .ZN(
        npu_inst_pe_1_7_2_n5) );
  INV_X1 npu_inst_pe_1_7_2_U105 ( .A(npu_inst_n34), .ZN(npu_inst_pe_1_7_2_n2)
         );
  AOI22_X1 npu_inst_pe_1_7_2_U104 ( .A1(npu_inst_pe_1_7_2_n38), .A2(
        int_i_data_v_npu[11]), .B1(npu_inst_pe_1_7_2_n113), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_2_n39) );
  INV_X1 npu_inst_pe_1_7_2_U103 ( .A(npu_inst_pe_1_7_2_n39), .ZN(
        npu_inst_pe_1_7_2_n111) );
  AOI22_X1 npu_inst_pe_1_7_2_U102 ( .A1(npu_inst_pe_1_7_2_n38), .A2(
        int_i_data_v_npu[10]), .B1(npu_inst_pe_1_7_2_n113), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_2_n37) );
  INV_X1 npu_inst_pe_1_7_2_U99 ( .A(npu_inst_pe_1_7_2_n37), .ZN(
        npu_inst_pe_1_7_2_n112) );
  AOI22_X1 npu_inst_pe_1_7_2_U98 ( .A1(int_i_data_v_npu[11]), .A2(
        npu_inst_pe_1_7_2_n58), .B1(npu_inst_pe_1_7_2_n118), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_2_n59) );
  INV_X1 npu_inst_pe_1_7_2_U97 ( .A(npu_inst_pe_1_7_2_n59), .ZN(
        npu_inst_pe_1_7_2_n101) );
  AOI22_X1 npu_inst_pe_1_7_2_U96 ( .A1(int_i_data_v_npu[10]), .A2(
        npu_inst_pe_1_7_2_n58), .B1(npu_inst_pe_1_7_2_n118), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_2_n57) );
  INV_X1 npu_inst_pe_1_7_2_U95 ( .A(npu_inst_pe_1_7_2_n57), .ZN(
        npu_inst_pe_1_7_2_n102) );
  AOI22_X1 npu_inst_pe_1_7_2_U94 ( .A1(int_i_data_v_npu[11]), .A2(
        npu_inst_pe_1_7_2_n54), .B1(npu_inst_pe_1_7_2_n117), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_2_n55) );
  INV_X1 npu_inst_pe_1_7_2_U93 ( .A(npu_inst_pe_1_7_2_n55), .ZN(
        npu_inst_pe_1_7_2_n103) );
  AOI22_X1 npu_inst_pe_1_7_2_U92 ( .A1(int_i_data_v_npu[10]), .A2(
        npu_inst_pe_1_7_2_n54), .B1(npu_inst_pe_1_7_2_n117), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_2_n53) );
  INV_X1 npu_inst_pe_1_7_2_U91 ( .A(npu_inst_pe_1_7_2_n53), .ZN(
        npu_inst_pe_1_7_2_n104) );
  AOI22_X1 npu_inst_pe_1_7_2_U90 ( .A1(int_i_data_v_npu[11]), .A2(
        npu_inst_pe_1_7_2_n50), .B1(npu_inst_pe_1_7_2_n116), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_2_n51) );
  INV_X1 npu_inst_pe_1_7_2_U89 ( .A(npu_inst_pe_1_7_2_n51), .ZN(
        npu_inst_pe_1_7_2_n105) );
  AOI22_X1 npu_inst_pe_1_7_2_U88 ( .A1(int_i_data_v_npu[10]), .A2(
        npu_inst_pe_1_7_2_n50), .B1(npu_inst_pe_1_7_2_n116), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_2_n49) );
  INV_X1 npu_inst_pe_1_7_2_U87 ( .A(npu_inst_pe_1_7_2_n49), .ZN(
        npu_inst_pe_1_7_2_n106) );
  AOI22_X1 npu_inst_pe_1_7_2_U86 ( .A1(int_i_data_v_npu[11]), .A2(
        npu_inst_pe_1_7_2_n46), .B1(npu_inst_pe_1_7_2_n115), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_2_n47) );
  INV_X1 npu_inst_pe_1_7_2_U85 ( .A(npu_inst_pe_1_7_2_n47), .ZN(
        npu_inst_pe_1_7_2_n107) );
  AOI22_X1 npu_inst_pe_1_7_2_U84 ( .A1(int_i_data_v_npu[10]), .A2(
        npu_inst_pe_1_7_2_n46), .B1(npu_inst_pe_1_7_2_n115), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_2_n45) );
  INV_X1 npu_inst_pe_1_7_2_U83 ( .A(npu_inst_pe_1_7_2_n45), .ZN(
        npu_inst_pe_1_7_2_n108) );
  AOI22_X1 npu_inst_pe_1_7_2_U82 ( .A1(int_i_data_v_npu[11]), .A2(
        npu_inst_pe_1_7_2_n42), .B1(npu_inst_pe_1_7_2_n114), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_2_n43) );
  INV_X1 npu_inst_pe_1_7_2_U81 ( .A(npu_inst_pe_1_7_2_n43), .ZN(
        npu_inst_pe_1_7_2_n109) );
  AOI22_X1 npu_inst_pe_1_7_2_U80 ( .A1(int_i_data_v_npu[10]), .A2(
        npu_inst_pe_1_7_2_n42), .B1(npu_inst_pe_1_7_2_n114), .B2(
        npu_inst_pe_1_7_2_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_2_n41) );
  INV_X1 npu_inst_pe_1_7_2_U79 ( .A(npu_inst_pe_1_7_2_n41), .ZN(
        npu_inst_pe_1_7_2_n110) );
  AND2_X1 npu_inst_pe_1_7_2_U78 ( .A1(npu_inst_pe_1_7_2_N93), .A2(npu_inst_n34), .ZN(npu_inst_int_data_y_7__2__0_) );
  NAND2_X1 npu_inst_pe_1_7_2_U77 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_2_n60), .ZN(npu_inst_pe_1_7_2_n74) );
  OAI21_X1 npu_inst_pe_1_7_2_U76 ( .B1(npu_inst_pe_1_7_2_n63), .B2(
        npu_inst_pe_1_7_2_n60), .A(npu_inst_pe_1_7_2_n74), .ZN(
        npu_inst_pe_1_7_2_n97) );
  NAND2_X1 npu_inst_pe_1_7_2_U75 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_2_n60), .ZN(npu_inst_pe_1_7_2_n73) );
  OAI21_X1 npu_inst_pe_1_7_2_U74 ( .B1(npu_inst_pe_1_7_2_n61), .B2(
        npu_inst_pe_1_7_2_n60), .A(npu_inst_pe_1_7_2_n73), .ZN(
        npu_inst_pe_1_7_2_n96) );
  NAND2_X1 npu_inst_pe_1_7_2_U73 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_2_n56), .ZN(npu_inst_pe_1_7_2_n72) );
  OAI21_X1 npu_inst_pe_1_7_2_U72 ( .B1(npu_inst_pe_1_7_2_n63), .B2(
        npu_inst_pe_1_7_2_n56), .A(npu_inst_pe_1_7_2_n72), .ZN(
        npu_inst_pe_1_7_2_n95) );
  NAND2_X1 npu_inst_pe_1_7_2_U71 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_2_n56), .ZN(npu_inst_pe_1_7_2_n71) );
  OAI21_X1 npu_inst_pe_1_7_2_U70 ( .B1(npu_inst_pe_1_7_2_n61), .B2(
        npu_inst_pe_1_7_2_n56), .A(npu_inst_pe_1_7_2_n71), .ZN(
        npu_inst_pe_1_7_2_n94) );
  NAND2_X1 npu_inst_pe_1_7_2_U69 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_2_n52), .ZN(npu_inst_pe_1_7_2_n70) );
  OAI21_X1 npu_inst_pe_1_7_2_U68 ( .B1(npu_inst_pe_1_7_2_n63), .B2(
        npu_inst_pe_1_7_2_n52), .A(npu_inst_pe_1_7_2_n70), .ZN(
        npu_inst_pe_1_7_2_n93) );
  NAND2_X1 npu_inst_pe_1_7_2_U67 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_2_n52), .ZN(npu_inst_pe_1_7_2_n69) );
  OAI21_X1 npu_inst_pe_1_7_2_U66 ( .B1(npu_inst_pe_1_7_2_n61), .B2(
        npu_inst_pe_1_7_2_n52), .A(npu_inst_pe_1_7_2_n69), .ZN(
        npu_inst_pe_1_7_2_n92) );
  NAND2_X1 npu_inst_pe_1_7_2_U65 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_2_n48), .ZN(npu_inst_pe_1_7_2_n68) );
  OAI21_X1 npu_inst_pe_1_7_2_U64 ( .B1(npu_inst_pe_1_7_2_n63), .B2(
        npu_inst_pe_1_7_2_n48), .A(npu_inst_pe_1_7_2_n68), .ZN(
        npu_inst_pe_1_7_2_n91) );
  NAND2_X1 npu_inst_pe_1_7_2_U63 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_2_n48), .ZN(npu_inst_pe_1_7_2_n67) );
  OAI21_X1 npu_inst_pe_1_7_2_U62 ( .B1(npu_inst_pe_1_7_2_n61), .B2(
        npu_inst_pe_1_7_2_n48), .A(npu_inst_pe_1_7_2_n67), .ZN(
        npu_inst_pe_1_7_2_n90) );
  NAND2_X1 npu_inst_pe_1_7_2_U61 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_2_n44), .ZN(npu_inst_pe_1_7_2_n66) );
  OAI21_X1 npu_inst_pe_1_7_2_U60 ( .B1(npu_inst_pe_1_7_2_n63), .B2(
        npu_inst_pe_1_7_2_n44), .A(npu_inst_pe_1_7_2_n66), .ZN(
        npu_inst_pe_1_7_2_n89) );
  NAND2_X1 npu_inst_pe_1_7_2_U59 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_2_n44), .ZN(npu_inst_pe_1_7_2_n65) );
  OAI21_X1 npu_inst_pe_1_7_2_U58 ( .B1(npu_inst_pe_1_7_2_n61), .B2(
        npu_inst_pe_1_7_2_n44), .A(npu_inst_pe_1_7_2_n65), .ZN(
        npu_inst_pe_1_7_2_n88) );
  NAND2_X1 npu_inst_pe_1_7_2_U57 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_2_n40), .ZN(npu_inst_pe_1_7_2_n64) );
  OAI21_X1 npu_inst_pe_1_7_2_U56 ( .B1(npu_inst_pe_1_7_2_n63), .B2(
        npu_inst_pe_1_7_2_n40), .A(npu_inst_pe_1_7_2_n64), .ZN(
        npu_inst_pe_1_7_2_n87) );
  NAND2_X1 npu_inst_pe_1_7_2_U55 ( .A1(npu_inst_pe_1_7_2_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_2_n40), .ZN(npu_inst_pe_1_7_2_n62) );
  OAI21_X1 npu_inst_pe_1_7_2_U54 ( .B1(npu_inst_pe_1_7_2_n61), .B2(
        npu_inst_pe_1_7_2_n40), .A(npu_inst_pe_1_7_2_n62), .ZN(
        npu_inst_pe_1_7_2_n86) );
  AND2_X1 npu_inst_pe_1_7_2_U53 ( .A1(npu_inst_n34), .A2(npu_inst_pe_1_7_2_N94), .ZN(npu_inst_int_data_y_7__2__1_) );
  AOI22_X1 npu_inst_pe_1_7_2_U52 ( .A1(npu_inst_n34), .A2(int_i_data_v_npu[11]), .B1(npu_inst_pe_1_7_2_n2), .B2(npu_inst_int_data_x_7__3__1_), .ZN(
        npu_inst_pe_1_7_2_n63) );
  AOI22_X1 npu_inst_pe_1_7_2_U51 ( .A1(npu_inst_n34), .A2(int_i_data_v_npu[10]), .B1(npu_inst_pe_1_7_2_n2), .B2(npu_inst_int_data_x_7__3__0_), .ZN(
        npu_inst_pe_1_7_2_n61) );
  AOI222_X1 npu_inst_pe_1_7_2_U50 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N73), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N65), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n84) );
  INV_X1 npu_inst_pe_1_7_2_U49 ( .A(npu_inst_pe_1_7_2_n84), .ZN(
        npu_inst_pe_1_7_2_n100) );
  AOI222_X1 npu_inst_pe_1_7_2_U48 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N74), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N66), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n83) );
  INV_X1 npu_inst_pe_1_7_2_U47 ( .A(npu_inst_pe_1_7_2_n83), .ZN(
        npu_inst_pe_1_7_2_n99) );
  AOI222_X1 npu_inst_pe_1_7_2_U46 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N75), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N67), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n82) );
  INV_X1 npu_inst_pe_1_7_2_U45 ( .A(npu_inst_pe_1_7_2_n82), .ZN(
        npu_inst_pe_1_7_2_n98) );
  AOI222_X1 npu_inst_pe_1_7_2_U44 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N76), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N68), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n81) );
  INV_X1 npu_inst_pe_1_7_2_U43 ( .A(npu_inst_pe_1_7_2_n81), .ZN(
        npu_inst_pe_1_7_2_n36) );
  AOI222_X1 npu_inst_pe_1_7_2_U42 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N77), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N69), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n80) );
  INV_X1 npu_inst_pe_1_7_2_U41 ( .A(npu_inst_pe_1_7_2_n80), .ZN(
        npu_inst_pe_1_7_2_n35) );
  AOI222_X1 npu_inst_pe_1_7_2_U40 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N78), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N70), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n79) );
  INV_X1 npu_inst_pe_1_7_2_U39 ( .A(npu_inst_pe_1_7_2_n79), .ZN(
        npu_inst_pe_1_7_2_n34) );
  AOI222_X1 npu_inst_pe_1_7_2_U38 ( .A1(1'b0), .A2(npu_inst_pe_1_7_2_n1), .B1(
        npu_inst_pe_1_7_2_N79), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N71), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n78) );
  INV_X1 npu_inst_pe_1_7_2_U37 ( .A(npu_inst_pe_1_7_2_n78), .ZN(
        npu_inst_pe_1_7_2_n33) );
  AOI222_X1 npu_inst_pe_1_7_2_U36 ( .A1(npu_inst_pe_1_7_2_n1), .A2(1'b0), .B1(
        npu_inst_pe_1_7_2_N80), .B2(npu_inst_pe_1_7_2_n76), .C1(
        npu_inst_pe_1_7_2_N72), .C2(npu_inst_pe_1_7_2_n77), .ZN(
        npu_inst_pe_1_7_2_n75) );
  INV_X1 npu_inst_pe_1_7_2_U35 ( .A(npu_inst_pe_1_7_2_n75), .ZN(
        npu_inst_pe_1_7_2_n32) );
  AND2_X1 npu_inst_pe_1_7_2_U34 ( .A1(npu_inst_int_data_x_7__2__1_), .A2(
        npu_inst_pe_1_7_2_int_q_weight_1_), .ZN(npu_inst_pe_1_7_2_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_2_U33 ( .A1(npu_inst_int_data_x_7__2__0_), .A2(
        npu_inst_pe_1_7_2_int_q_weight_1_), .ZN(npu_inst_pe_1_7_2_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_2_U32 ( .A(npu_inst_pe_1_7_2_int_data_1_), .ZN(
        npu_inst_pe_1_7_2_n13) );
  NOR3_X1 npu_inst_pe_1_7_2_U31 ( .A1(npu_inst_pe_1_7_2_n26), .A2(npu_inst_n34), .A3(npu_inst_int_ckg[5]), .ZN(npu_inst_pe_1_7_2_n85) );
  OR2_X1 npu_inst_pe_1_7_2_U30 ( .A1(npu_inst_pe_1_7_2_n85), .A2(
        npu_inst_pe_1_7_2_n1), .ZN(npu_inst_pe_1_7_2_N84) );
  INV_X1 npu_inst_pe_1_7_2_U29 ( .A(npu_inst_pe_1_7_2_int_data_0_), .ZN(
        npu_inst_pe_1_7_2_n12) );
  INV_X1 npu_inst_pe_1_7_2_U28 ( .A(npu_inst_n49), .ZN(npu_inst_pe_1_7_2_n4)
         );
  OR3_X1 npu_inst_pe_1_7_2_U27 ( .A1(npu_inst_pe_1_7_2_n5), .A2(
        npu_inst_pe_1_7_2_n7), .A3(npu_inst_pe_1_7_2_n4), .ZN(
        npu_inst_pe_1_7_2_n56) );
  OR3_X1 npu_inst_pe_1_7_2_U26 ( .A1(npu_inst_pe_1_7_2_n4), .A2(
        npu_inst_pe_1_7_2_n7), .A3(npu_inst_pe_1_7_2_n6), .ZN(
        npu_inst_pe_1_7_2_n48) );
  INV_X1 npu_inst_pe_1_7_2_U25 ( .A(npu_inst_pe_1_7_2_n4), .ZN(
        npu_inst_pe_1_7_2_n3) );
  OR3_X1 npu_inst_pe_1_7_2_U24 ( .A1(npu_inst_pe_1_7_2_n3), .A2(
        npu_inst_pe_1_7_2_n7), .A3(npu_inst_pe_1_7_2_n6), .ZN(
        npu_inst_pe_1_7_2_n52) );
  OR3_X1 npu_inst_pe_1_7_2_U23 ( .A1(npu_inst_pe_1_7_2_n5), .A2(
        npu_inst_pe_1_7_2_n7), .A3(npu_inst_pe_1_7_2_n3), .ZN(
        npu_inst_pe_1_7_2_n60) );
  BUF_X1 npu_inst_pe_1_7_2_U22 ( .A(npu_inst_n12), .Z(npu_inst_pe_1_7_2_n1) );
  NOR2_X1 npu_inst_pe_1_7_2_U21 ( .A1(npu_inst_pe_1_7_2_n60), .A2(
        npu_inst_pe_1_7_2_n2), .ZN(npu_inst_pe_1_7_2_n58) );
  NOR2_X1 npu_inst_pe_1_7_2_U20 ( .A1(npu_inst_pe_1_7_2_n56), .A2(
        npu_inst_pe_1_7_2_n2), .ZN(npu_inst_pe_1_7_2_n54) );
  NOR2_X1 npu_inst_pe_1_7_2_U19 ( .A1(npu_inst_pe_1_7_2_n52), .A2(
        npu_inst_pe_1_7_2_n2), .ZN(npu_inst_pe_1_7_2_n50) );
  NOR2_X1 npu_inst_pe_1_7_2_U18 ( .A1(npu_inst_pe_1_7_2_n48), .A2(
        npu_inst_pe_1_7_2_n2), .ZN(npu_inst_pe_1_7_2_n46) );
  NOR2_X1 npu_inst_pe_1_7_2_U17 ( .A1(npu_inst_pe_1_7_2_n40), .A2(
        npu_inst_pe_1_7_2_n2), .ZN(npu_inst_pe_1_7_2_n38) );
  NOR2_X1 npu_inst_pe_1_7_2_U16 ( .A1(npu_inst_pe_1_7_2_n44), .A2(
        npu_inst_pe_1_7_2_n2), .ZN(npu_inst_pe_1_7_2_n42) );
  BUF_X1 npu_inst_pe_1_7_2_U15 ( .A(npu_inst_n75), .Z(npu_inst_pe_1_7_2_n7) );
  INV_X1 npu_inst_pe_1_7_2_U14 ( .A(npu_inst_n104), .ZN(npu_inst_pe_1_7_2_n11)
         );
  INV_X1 npu_inst_pe_1_7_2_U13 ( .A(npu_inst_pe_1_7_2_n38), .ZN(
        npu_inst_pe_1_7_2_n113) );
  INV_X1 npu_inst_pe_1_7_2_U12 ( .A(npu_inst_pe_1_7_2_n58), .ZN(
        npu_inst_pe_1_7_2_n118) );
  INV_X1 npu_inst_pe_1_7_2_U11 ( .A(npu_inst_pe_1_7_2_n54), .ZN(
        npu_inst_pe_1_7_2_n117) );
  INV_X1 npu_inst_pe_1_7_2_U10 ( .A(npu_inst_pe_1_7_2_n50), .ZN(
        npu_inst_pe_1_7_2_n116) );
  INV_X1 npu_inst_pe_1_7_2_U9 ( .A(npu_inst_pe_1_7_2_n46), .ZN(
        npu_inst_pe_1_7_2_n115) );
  INV_X1 npu_inst_pe_1_7_2_U8 ( .A(npu_inst_pe_1_7_2_n42), .ZN(
        npu_inst_pe_1_7_2_n114) );
  BUF_X1 npu_inst_pe_1_7_2_U7 ( .A(npu_inst_pe_1_7_2_n11), .Z(
        npu_inst_pe_1_7_2_n10) );
  BUF_X1 npu_inst_pe_1_7_2_U6 ( .A(npu_inst_pe_1_7_2_n11), .Z(
        npu_inst_pe_1_7_2_n9) );
  BUF_X1 npu_inst_pe_1_7_2_U5 ( .A(npu_inst_pe_1_7_2_n11), .Z(
        npu_inst_pe_1_7_2_n8) );
  NOR2_X1 npu_inst_pe_1_7_2_U4 ( .A1(npu_inst_pe_1_7_2_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_2_n1), .ZN(npu_inst_pe_1_7_2_n76) );
  NOR2_X1 npu_inst_pe_1_7_2_U3 ( .A1(npu_inst_pe_1_7_2_n27), .A2(
        npu_inst_pe_1_7_2_n1), .ZN(npu_inst_pe_1_7_2_n77) );
  FA_X1 npu_inst_pe_1_7_2_sub_77_U2_1 ( .A(npu_inst_int_data_res_7__2__1_), 
        .B(npu_inst_pe_1_7_2_n13), .CI(npu_inst_pe_1_7_2_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_7_2_sub_77_carry_2_), .S(npu_inst_pe_1_7_2_N66) );
  FA_X1 npu_inst_pe_1_7_2_add_79_U1_1 ( .A(npu_inst_int_data_res_7__2__1_), 
        .B(npu_inst_pe_1_7_2_int_data_1_), .CI(
        npu_inst_pe_1_7_2_add_79_carry_1_), .CO(
        npu_inst_pe_1_7_2_add_79_carry_2_), .S(npu_inst_pe_1_7_2_N74) );
  NAND3_X1 npu_inst_pe_1_7_2_U101 ( .A1(npu_inst_pe_1_7_2_n4), .A2(
        npu_inst_pe_1_7_2_n6), .A3(npu_inst_pe_1_7_2_n7), .ZN(
        npu_inst_pe_1_7_2_n44) );
  NAND3_X1 npu_inst_pe_1_7_2_U100 ( .A1(npu_inst_pe_1_7_2_n3), .A2(
        npu_inst_pe_1_7_2_n6), .A3(npu_inst_pe_1_7_2_n7), .ZN(
        npu_inst_pe_1_7_2_n40) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_2_n33), .CK(
        npu_inst_pe_1_7_2_net3144), .RN(npu_inst_pe_1_7_2_n8), .Q(
        npu_inst_int_data_res_7__2__6_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_2_n34), .CK(
        npu_inst_pe_1_7_2_net3144), .RN(npu_inst_pe_1_7_2_n8), .Q(
        npu_inst_int_data_res_7__2__5_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_2_n35), .CK(
        npu_inst_pe_1_7_2_net3144), .RN(npu_inst_pe_1_7_2_n8), .Q(
        npu_inst_int_data_res_7__2__4_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_2_n36), .CK(
        npu_inst_pe_1_7_2_net3144), .RN(npu_inst_pe_1_7_2_n8), .Q(
        npu_inst_int_data_res_7__2__3_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_2_n98), .CK(
        npu_inst_pe_1_7_2_net3144), .RN(npu_inst_pe_1_7_2_n8), .Q(
        npu_inst_int_data_res_7__2__2_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_2_n99), .CK(
        npu_inst_pe_1_7_2_net3144), .RN(npu_inst_pe_1_7_2_n8), .Q(
        npu_inst_int_data_res_7__2__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_2_n32), .CK(
        npu_inst_pe_1_7_2_net3144), .RN(npu_inst_pe_1_7_2_n8), .Q(
        npu_inst_int_data_res_7__2__7_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_2_n100), 
        .CK(npu_inst_pe_1_7_2_net3144), .RN(npu_inst_pe_1_7_2_n8), .Q(
        npu_inst_int_data_res_7__2__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_weight_reg_0_ ( .D(npu_inst_n90), .CK(
        npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n8), .Q(
        npu_inst_pe_1_7_2_int_q_weight_0_), .QN(npu_inst_pe_1_7_2_n27) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_weight_reg_1_ ( .D(npu_inst_n96), .CK(
        npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n8), .Q(
        npu_inst_pe_1_7_2_int_q_weight_1_), .QN(npu_inst_pe_1_7_2_n26) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_2_n112), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n8), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_2_n111), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n8), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_2_n110), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_2_n109), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_2_n108), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_2_n107), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_2_n106), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_2_n105), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_2_n104), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_2_n103), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_2_n102), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_2_n101), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_2_n86), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_2_n87), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n9), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_2_n88), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_2_n89), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_2_n90), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_2_n91), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_2_n92), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_2_n93), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_2_n94), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_2_n95), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_2_n96), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_2_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_2_n97), 
        .CK(npu_inst_pe_1_7_2_net3150), .RN(npu_inst_pe_1_7_2_n10), .Q(
        npu_inst_pe_1_7_2_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_2_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_2_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_2_net3144) );
  CLKGATETST_X1 npu_inst_pe_1_7_2_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n43), .SE(1'b0), .GCK(npu_inst_pe_1_7_2_net3150) );
  MUX2_X1 npu_inst_pe_1_7_3_U153 ( .A(npu_inst_pe_1_7_3_n31), .B(
        npu_inst_pe_1_7_3_n28), .S(npu_inst_pe_1_7_3_n7), .Z(
        npu_inst_pe_1_7_3_N93) );
  MUX2_X1 npu_inst_pe_1_7_3_U152 ( .A(npu_inst_pe_1_7_3_n30), .B(
        npu_inst_pe_1_7_3_n29), .S(npu_inst_pe_1_7_3_n5), .Z(
        npu_inst_pe_1_7_3_n31) );
  MUX2_X1 npu_inst_pe_1_7_3_U151 ( .A(npu_inst_pe_1_7_3_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_3_n3), .Z(
        npu_inst_pe_1_7_3_n30) );
  MUX2_X1 npu_inst_pe_1_7_3_U150 ( .A(npu_inst_pe_1_7_3_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_3_n3), .Z(
        npu_inst_pe_1_7_3_n29) );
  MUX2_X1 npu_inst_pe_1_7_3_U149 ( .A(npu_inst_pe_1_7_3_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_3_n3), .Z(
        npu_inst_pe_1_7_3_n28) );
  MUX2_X1 npu_inst_pe_1_7_3_U148 ( .A(npu_inst_pe_1_7_3_n25), .B(
        npu_inst_pe_1_7_3_n22), .S(npu_inst_pe_1_7_3_n7), .Z(
        npu_inst_pe_1_7_3_N94) );
  MUX2_X1 npu_inst_pe_1_7_3_U147 ( .A(npu_inst_pe_1_7_3_n24), .B(
        npu_inst_pe_1_7_3_n23), .S(npu_inst_pe_1_7_3_n5), .Z(
        npu_inst_pe_1_7_3_n25) );
  MUX2_X1 npu_inst_pe_1_7_3_U146 ( .A(npu_inst_pe_1_7_3_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_3_n3), .Z(
        npu_inst_pe_1_7_3_n24) );
  MUX2_X1 npu_inst_pe_1_7_3_U145 ( .A(npu_inst_pe_1_7_3_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_3_n3), .Z(
        npu_inst_pe_1_7_3_n23) );
  MUX2_X1 npu_inst_pe_1_7_3_U144 ( .A(npu_inst_pe_1_7_3_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_3_n3), .Z(
        npu_inst_pe_1_7_3_n22) );
  MUX2_X1 npu_inst_pe_1_7_3_U143 ( .A(npu_inst_pe_1_7_3_n21), .B(
        npu_inst_pe_1_7_3_n18), .S(npu_inst_pe_1_7_3_n7), .Z(
        npu_inst_int_data_x_7__3__1_) );
  MUX2_X1 npu_inst_pe_1_7_3_U142 ( .A(npu_inst_pe_1_7_3_n20), .B(
        npu_inst_pe_1_7_3_n19), .S(npu_inst_pe_1_7_3_n5), .Z(
        npu_inst_pe_1_7_3_n21) );
  MUX2_X1 npu_inst_pe_1_7_3_U141 ( .A(npu_inst_pe_1_7_3_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_3_n3), .Z(
        npu_inst_pe_1_7_3_n20) );
  MUX2_X1 npu_inst_pe_1_7_3_U140 ( .A(npu_inst_pe_1_7_3_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_3_n3), .Z(
        npu_inst_pe_1_7_3_n19) );
  MUX2_X1 npu_inst_pe_1_7_3_U139 ( .A(npu_inst_pe_1_7_3_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_3_n3), .Z(
        npu_inst_pe_1_7_3_n18) );
  MUX2_X1 npu_inst_pe_1_7_3_U138 ( .A(npu_inst_pe_1_7_3_n17), .B(
        npu_inst_pe_1_7_3_n14), .S(npu_inst_pe_1_7_3_n7), .Z(
        npu_inst_int_data_x_7__3__0_) );
  MUX2_X1 npu_inst_pe_1_7_3_U137 ( .A(npu_inst_pe_1_7_3_n16), .B(
        npu_inst_pe_1_7_3_n15), .S(npu_inst_pe_1_7_3_n5), .Z(
        npu_inst_pe_1_7_3_n17) );
  MUX2_X1 npu_inst_pe_1_7_3_U136 ( .A(npu_inst_pe_1_7_3_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_3_n3), .Z(
        npu_inst_pe_1_7_3_n16) );
  MUX2_X1 npu_inst_pe_1_7_3_U135 ( .A(npu_inst_pe_1_7_3_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_3_n3), .Z(
        npu_inst_pe_1_7_3_n15) );
  MUX2_X1 npu_inst_pe_1_7_3_U134 ( .A(npu_inst_pe_1_7_3_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_3_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_3_n3), .Z(
        npu_inst_pe_1_7_3_n14) );
  XOR2_X1 npu_inst_pe_1_7_3_U133 ( .A(npu_inst_pe_1_7_3_int_data_0_), .B(
        npu_inst_int_data_res_7__3__0_), .Z(npu_inst_pe_1_7_3_N73) );
  AND2_X1 npu_inst_pe_1_7_3_U132 ( .A1(npu_inst_int_data_res_7__3__0_), .A2(
        npu_inst_pe_1_7_3_int_data_0_), .ZN(npu_inst_pe_1_7_3_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_3_U131 ( .A(npu_inst_int_data_res_7__3__0_), .B(
        npu_inst_pe_1_7_3_n12), .ZN(npu_inst_pe_1_7_3_N65) );
  OR2_X1 npu_inst_pe_1_7_3_U130 ( .A1(npu_inst_pe_1_7_3_n12), .A2(
        npu_inst_int_data_res_7__3__0_), .ZN(npu_inst_pe_1_7_3_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_3_U129 ( .A(npu_inst_int_data_res_7__3__2_), .B(
        npu_inst_pe_1_7_3_add_79_carry_2_), .Z(npu_inst_pe_1_7_3_N75) );
  AND2_X1 npu_inst_pe_1_7_3_U128 ( .A1(npu_inst_pe_1_7_3_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_7__3__2_), .ZN(
        npu_inst_pe_1_7_3_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_3_U127 ( .A(npu_inst_int_data_res_7__3__3_), .B(
        npu_inst_pe_1_7_3_add_79_carry_3_), .Z(npu_inst_pe_1_7_3_N76) );
  AND2_X1 npu_inst_pe_1_7_3_U126 ( .A1(npu_inst_pe_1_7_3_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_7__3__3_), .ZN(
        npu_inst_pe_1_7_3_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_3_U125 ( .A(npu_inst_int_data_res_7__3__4_), .B(
        npu_inst_pe_1_7_3_add_79_carry_4_), .Z(npu_inst_pe_1_7_3_N77) );
  AND2_X1 npu_inst_pe_1_7_3_U124 ( .A1(npu_inst_pe_1_7_3_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_7__3__4_), .ZN(
        npu_inst_pe_1_7_3_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_3_U123 ( .A(npu_inst_int_data_res_7__3__5_), .B(
        npu_inst_pe_1_7_3_add_79_carry_5_), .Z(npu_inst_pe_1_7_3_N78) );
  AND2_X1 npu_inst_pe_1_7_3_U122 ( .A1(npu_inst_pe_1_7_3_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_7__3__5_), .ZN(
        npu_inst_pe_1_7_3_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_3_U121 ( .A(npu_inst_int_data_res_7__3__6_), .B(
        npu_inst_pe_1_7_3_add_79_carry_6_), .Z(npu_inst_pe_1_7_3_N79) );
  AND2_X1 npu_inst_pe_1_7_3_U120 ( .A1(npu_inst_pe_1_7_3_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_7__3__6_), .ZN(
        npu_inst_pe_1_7_3_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_3_U119 ( .A(npu_inst_int_data_res_7__3__7_), .B(
        npu_inst_pe_1_7_3_add_79_carry_7_), .Z(npu_inst_pe_1_7_3_N80) );
  XNOR2_X1 npu_inst_pe_1_7_3_U118 ( .A(npu_inst_pe_1_7_3_sub_77_carry_2_), .B(
        npu_inst_int_data_res_7__3__2_), .ZN(npu_inst_pe_1_7_3_N67) );
  OR2_X1 npu_inst_pe_1_7_3_U117 ( .A1(npu_inst_int_data_res_7__3__2_), .A2(
        npu_inst_pe_1_7_3_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_7_3_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_3_U116 ( .A(npu_inst_pe_1_7_3_sub_77_carry_3_), .B(
        npu_inst_int_data_res_7__3__3_), .ZN(npu_inst_pe_1_7_3_N68) );
  OR2_X1 npu_inst_pe_1_7_3_U115 ( .A1(npu_inst_int_data_res_7__3__3_), .A2(
        npu_inst_pe_1_7_3_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_7_3_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_3_U114 ( .A(npu_inst_pe_1_7_3_sub_77_carry_4_), .B(
        npu_inst_int_data_res_7__3__4_), .ZN(npu_inst_pe_1_7_3_N69) );
  OR2_X1 npu_inst_pe_1_7_3_U113 ( .A1(npu_inst_int_data_res_7__3__4_), .A2(
        npu_inst_pe_1_7_3_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_7_3_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_3_U112 ( .A(npu_inst_pe_1_7_3_sub_77_carry_5_), .B(
        npu_inst_int_data_res_7__3__5_), .ZN(npu_inst_pe_1_7_3_N70) );
  OR2_X1 npu_inst_pe_1_7_3_U111 ( .A1(npu_inst_int_data_res_7__3__5_), .A2(
        npu_inst_pe_1_7_3_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_7_3_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_3_U110 ( .A(npu_inst_pe_1_7_3_sub_77_carry_6_), .B(
        npu_inst_int_data_res_7__3__6_), .ZN(npu_inst_pe_1_7_3_N71) );
  OR2_X1 npu_inst_pe_1_7_3_U109 ( .A1(npu_inst_int_data_res_7__3__6_), .A2(
        npu_inst_pe_1_7_3_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_7_3_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_3_U108 ( .A(npu_inst_int_data_res_7__3__7_), .B(
        npu_inst_pe_1_7_3_sub_77_carry_7_), .ZN(npu_inst_pe_1_7_3_N72) );
  INV_X1 npu_inst_pe_1_7_3_U107 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_7_3_n6)
         );
  INV_X1 npu_inst_pe_1_7_3_U106 ( .A(npu_inst_pe_1_7_3_n6), .ZN(
        npu_inst_pe_1_7_3_n5) );
  INV_X1 npu_inst_pe_1_7_3_U105 ( .A(npu_inst_n34), .ZN(npu_inst_pe_1_7_3_n2)
         );
  AOI22_X1 npu_inst_pe_1_7_3_U104 ( .A1(npu_inst_pe_1_7_3_n38), .A2(
        int_i_data_v_npu[9]), .B1(npu_inst_pe_1_7_3_n113), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_3_n39) );
  INV_X1 npu_inst_pe_1_7_3_U103 ( .A(npu_inst_pe_1_7_3_n39), .ZN(
        npu_inst_pe_1_7_3_n111) );
  AOI22_X1 npu_inst_pe_1_7_3_U102 ( .A1(npu_inst_pe_1_7_3_n38), .A2(
        int_i_data_v_npu[8]), .B1(npu_inst_pe_1_7_3_n113), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_3_n37) );
  INV_X1 npu_inst_pe_1_7_3_U99 ( .A(npu_inst_pe_1_7_3_n37), .ZN(
        npu_inst_pe_1_7_3_n112) );
  AOI22_X1 npu_inst_pe_1_7_3_U98 ( .A1(int_i_data_v_npu[9]), .A2(
        npu_inst_pe_1_7_3_n58), .B1(npu_inst_pe_1_7_3_n118), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_3_n59) );
  INV_X1 npu_inst_pe_1_7_3_U97 ( .A(npu_inst_pe_1_7_3_n59), .ZN(
        npu_inst_pe_1_7_3_n101) );
  AOI22_X1 npu_inst_pe_1_7_3_U96 ( .A1(int_i_data_v_npu[8]), .A2(
        npu_inst_pe_1_7_3_n58), .B1(npu_inst_pe_1_7_3_n118), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_3_n57) );
  INV_X1 npu_inst_pe_1_7_3_U95 ( .A(npu_inst_pe_1_7_3_n57), .ZN(
        npu_inst_pe_1_7_3_n102) );
  AOI22_X1 npu_inst_pe_1_7_3_U94 ( .A1(int_i_data_v_npu[9]), .A2(
        npu_inst_pe_1_7_3_n54), .B1(npu_inst_pe_1_7_3_n117), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_3_n55) );
  INV_X1 npu_inst_pe_1_7_3_U93 ( .A(npu_inst_pe_1_7_3_n55), .ZN(
        npu_inst_pe_1_7_3_n103) );
  AOI22_X1 npu_inst_pe_1_7_3_U92 ( .A1(int_i_data_v_npu[8]), .A2(
        npu_inst_pe_1_7_3_n54), .B1(npu_inst_pe_1_7_3_n117), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_3_n53) );
  INV_X1 npu_inst_pe_1_7_3_U91 ( .A(npu_inst_pe_1_7_3_n53), .ZN(
        npu_inst_pe_1_7_3_n104) );
  AOI22_X1 npu_inst_pe_1_7_3_U90 ( .A1(int_i_data_v_npu[9]), .A2(
        npu_inst_pe_1_7_3_n50), .B1(npu_inst_pe_1_7_3_n116), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_3_n51) );
  INV_X1 npu_inst_pe_1_7_3_U89 ( .A(npu_inst_pe_1_7_3_n51), .ZN(
        npu_inst_pe_1_7_3_n105) );
  AOI22_X1 npu_inst_pe_1_7_3_U88 ( .A1(int_i_data_v_npu[8]), .A2(
        npu_inst_pe_1_7_3_n50), .B1(npu_inst_pe_1_7_3_n116), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_3_n49) );
  INV_X1 npu_inst_pe_1_7_3_U87 ( .A(npu_inst_pe_1_7_3_n49), .ZN(
        npu_inst_pe_1_7_3_n106) );
  AOI22_X1 npu_inst_pe_1_7_3_U86 ( .A1(int_i_data_v_npu[9]), .A2(
        npu_inst_pe_1_7_3_n46), .B1(npu_inst_pe_1_7_3_n115), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_3_n47) );
  INV_X1 npu_inst_pe_1_7_3_U85 ( .A(npu_inst_pe_1_7_3_n47), .ZN(
        npu_inst_pe_1_7_3_n107) );
  AOI22_X1 npu_inst_pe_1_7_3_U84 ( .A1(int_i_data_v_npu[8]), .A2(
        npu_inst_pe_1_7_3_n46), .B1(npu_inst_pe_1_7_3_n115), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_3_n45) );
  INV_X1 npu_inst_pe_1_7_3_U83 ( .A(npu_inst_pe_1_7_3_n45), .ZN(
        npu_inst_pe_1_7_3_n108) );
  AOI22_X1 npu_inst_pe_1_7_3_U82 ( .A1(int_i_data_v_npu[9]), .A2(
        npu_inst_pe_1_7_3_n42), .B1(npu_inst_pe_1_7_3_n114), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_3_n43) );
  INV_X1 npu_inst_pe_1_7_3_U81 ( .A(npu_inst_pe_1_7_3_n43), .ZN(
        npu_inst_pe_1_7_3_n109) );
  AOI22_X1 npu_inst_pe_1_7_3_U80 ( .A1(int_i_data_v_npu[8]), .A2(
        npu_inst_pe_1_7_3_n42), .B1(npu_inst_pe_1_7_3_n114), .B2(
        npu_inst_pe_1_7_3_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_3_n41) );
  INV_X1 npu_inst_pe_1_7_3_U79 ( .A(npu_inst_pe_1_7_3_n41), .ZN(
        npu_inst_pe_1_7_3_n110) );
  AND2_X1 npu_inst_pe_1_7_3_U78 ( .A1(npu_inst_pe_1_7_3_N93), .A2(npu_inst_n34), .ZN(npu_inst_int_data_y_7__3__0_) );
  NAND2_X1 npu_inst_pe_1_7_3_U77 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_3_n60), .ZN(npu_inst_pe_1_7_3_n74) );
  OAI21_X1 npu_inst_pe_1_7_3_U76 ( .B1(npu_inst_pe_1_7_3_n63), .B2(
        npu_inst_pe_1_7_3_n60), .A(npu_inst_pe_1_7_3_n74), .ZN(
        npu_inst_pe_1_7_3_n97) );
  NAND2_X1 npu_inst_pe_1_7_3_U75 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_3_n60), .ZN(npu_inst_pe_1_7_3_n73) );
  OAI21_X1 npu_inst_pe_1_7_3_U74 ( .B1(npu_inst_pe_1_7_3_n61), .B2(
        npu_inst_pe_1_7_3_n60), .A(npu_inst_pe_1_7_3_n73), .ZN(
        npu_inst_pe_1_7_3_n96) );
  NAND2_X1 npu_inst_pe_1_7_3_U73 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_3_n56), .ZN(npu_inst_pe_1_7_3_n72) );
  OAI21_X1 npu_inst_pe_1_7_3_U72 ( .B1(npu_inst_pe_1_7_3_n63), .B2(
        npu_inst_pe_1_7_3_n56), .A(npu_inst_pe_1_7_3_n72), .ZN(
        npu_inst_pe_1_7_3_n95) );
  NAND2_X1 npu_inst_pe_1_7_3_U71 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_3_n56), .ZN(npu_inst_pe_1_7_3_n71) );
  OAI21_X1 npu_inst_pe_1_7_3_U70 ( .B1(npu_inst_pe_1_7_3_n61), .B2(
        npu_inst_pe_1_7_3_n56), .A(npu_inst_pe_1_7_3_n71), .ZN(
        npu_inst_pe_1_7_3_n94) );
  NAND2_X1 npu_inst_pe_1_7_3_U69 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_3_n52), .ZN(npu_inst_pe_1_7_3_n70) );
  OAI21_X1 npu_inst_pe_1_7_3_U68 ( .B1(npu_inst_pe_1_7_3_n63), .B2(
        npu_inst_pe_1_7_3_n52), .A(npu_inst_pe_1_7_3_n70), .ZN(
        npu_inst_pe_1_7_3_n93) );
  NAND2_X1 npu_inst_pe_1_7_3_U67 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_3_n52), .ZN(npu_inst_pe_1_7_3_n69) );
  OAI21_X1 npu_inst_pe_1_7_3_U66 ( .B1(npu_inst_pe_1_7_3_n61), .B2(
        npu_inst_pe_1_7_3_n52), .A(npu_inst_pe_1_7_3_n69), .ZN(
        npu_inst_pe_1_7_3_n92) );
  NAND2_X1 npu_inst_pe_1_7_3_U65 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_3_n48), .ZN(npu_inst_pe_1_7_3_n68) );
  OAI21_X1 npu_inst_pe_1_7_3_U64 ( .B1(npu_inst_pe_1_7_3_n63), .B2(
        npu_inst_pe_1_7_3_n48), .A(npu_inst_pe_1_7_3_n68), .ZN(
        npu_inst_pe_1_7_3_n91) );
  NAND2_X1 npu_inst_pe_1_7_3_U63 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_3_n48), .ZN(npu_inst_pe_1_7_3_n67) );
  OAI21_X1 npu_inst_pe_1_7_3_U62 ( .B1(npu_inst_pe_1_7_3_n61), .B2(
        npu_inst_pe_1_7_3_n48), .A(npu_inst_pe_1_7_3_n67), .ZN(
        npu_inst_pe_1_7_3_n90) );
  NAND2_X1 npu_inst_pe_1_7_3_U61 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_3_n44), .ZN(npu_inst_pe_1_7_3_n66) );
  OAI21_X1 npu_inst_pe_1_7_3_U60 ( .B1(npu_inst_pe_1_7_3_n63), .B2(
        npu_inst_pe_1_7_3_n44), .A(npu_inst_pe_1_7_3_n66), .ZN(
        npu_inst_pe_1_7_3_n89) );
  NAND2_X1 npu_inst_pe_1_7_3_U59 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_3_n44), .ZN(npu_inst_pe_1_7_3_n65) );
  OAI21_X1 npu_inst_pe_1_7_3_U58 ( .B1(npu_inst_pe_1_7_3_n61), .B2(
        npu_inst_pe_1_7_3_n44), .A(npu_inst_pe_1_7_3_n65), .ZN(
        npu_inst_pe_1_7_3_n88) );
  NAND2_X1 npu_inst_pe_1_7_3_U57 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_3_n40), .ZN(npu_inst_pe_1_7_3_n64) );
  OAI21_X1 npu_inst_pe_1_7_3_U56 ( .B1(npu_inst_pe_1_7_3_n63), .B2(
        npu_inst_pe_1_7_3_n40), .A(npu_inst_pe_1_7_3_n64), .ZN(
        npu_inst_pe_1_7_3_n87) );
  NAND2_X1 npu_inst_pe_1_7_3_U55 ( .A1(npu_inst_pe_1_7_3_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_3_n40), .ZN(npu_inst_pe_1_7_3_n62) );
  OAI21_X1 npu_inst_pe_1_7_3_U54 ( .B1(npu_inst_pe_1_7_3_n61), .B2(
        npu_inst_pe_1_7_3_n40), .A(npu_inst_pe_1_7_3_n62), .ZN(
        npu_inst_pe_1_7_3_n86) );
  AND2_X1 npu_inst_pe_1_7_3_U53 ( .A1(npu_inst_n34), .A2(npu_inst_pe_1_7_3_N94), .ZN(npu_inst_int_data_y_7__3__1_) );
  AOI22_X1 npu_inst_pe_1_7_3_U52 ( .A1(npu_inst_n34), .A2(int_i_data_v_npu[9]), 
        .B1(npu_inst_pe_1_7_3_n2), .B2(npu_inst_int_data_x_7__4__1_), .ZN(
        npu_inst_pe_1_7_3_n63) );
  AOI22_X1 npu_inst_pe_1_7_3_U51 ( .A1(npu_inst_n34), .A2(int_i_data_v_npu[8]), 
        .B1(npu_inst_pe_1_7_3_n2), .B2(npu_inst_int_data_x_7__4__0_), .ZN(
        npu_inst_pe_1_7_3_n61) );
  AOI222_X1 npu_inst_pe_1_7_3_U50 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N73), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N65), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n84) );
  INV_X1 npu_inst_pe_1_7_3_U49 ( .A(npu_inst_pe_1_7_3_n84), .ZN(
        npu_inst_pe_1_7_3_n100) );
  AOI222_X1 npu_inst_pe_1_7_3_U48 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N74), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N66), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n83) );
  INV_X1 npu_inst_pe_1_7_3_U47 ( .A(npu_inst_pe_1_7_3_n83), .ZN(
        npu_inst_pe_1_7_3_n99) );
  AOI222_X1 npu_inst_pe_1_7_3_U46 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N75), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N67), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n82) );
  INV_X1 npu_inst_pe_1_7_3_U45 ( .A(npu_inst_pe_1_7_3_n82), .ZN(
        npu_inst_pe_1_7_3_n98) );
  AOI222_X1 npu_inst_pe_1_7_3_U44 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N76), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N68), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n81) );
  INV_X1 npu_inst_pe_1_7_3_U43 ( .A(npu_inst_pe_1_7_3_n81), .ZN(
        npu_inst_pe_1_7_3_n36) );
  AOI222_X1 npu_inst_pe_1_7_3_U42 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N77), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N69), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n80) );
  INV_X1 npu_inst_pe_1_7_3_U41 ( .A(npu_inst_pe_1_7_3_n80), .ZN(
        npu_inst_pe_1_7_3_n35) );
  AOI222_X1 npu_inst_pe_1_7_3_U40 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N78), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N70), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n79) );
  INV_X1 npu_inst_pe_1_7_3_U39 ( .A(npu_inst_pe_1_7_3_n79), .ZN(
        npu_inst_pe_1_7_3_n34) );
  AOI222_X1 npu_inst_pe_1_7_3_U38 ( .A1(1'b0), .A2(npu_inst_pe_1_7_3_n1), .B1(
        npu_inst_pe_1_7_3_N79), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N71), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n78) );
  INV_X1 npu_inst_pe_1_7_3_U37 ( .A(npu_inst_pe_1_7_3_n78), .ZN(
        npu_inst_pe_1_7_3_n33) );
  AOI222_X1 npu_inst_pe_1_7_3_U36 ( .A1(npu_inst_pe_1_7_3_n1), .A2(1'b0), .B1(
        npu_inst_pe_1_7_3_N80), .B2(npu_inst_pe_1_7_3_n76), .C1(
        npu_inst_pe_1_7_3_N72), .C2(npu_inst_pe_1_7_3_n77), .ZN(
        npu_inst_pe_1_7_3_n75) );
  INV_X1 npu_inst_pe_1_7_3_U35 ( .A(npu_inst_pe_1_7_3_n75), .ZN(
        npu_inst_pe_1_7_3_n32) );
  AND2_X1 npu_inst_pe_1_7_3_U34 ( .A1(npu_inst_int_data_x_7__3__1_), .A2(
        npu_inst_pe_1_7_3_int_q_weight_1_), .ZN(npu_inst_pe_1_7_3_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_3_U33 ( .A1(npu_inst_int_data_x_7__3__0_), .A2(
        npu_inst_pe_1_7_3_int_q_weight_1_), .ZN(npu_inst_pe_1_7_3_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_3_U32 ( .A(npu_inst_pe_1_7_3_int_data_1_), .ZN(
        npu_inst_pe_1_7_3_n13) );
  NOR3_X1 npu_inst_pe_1_7_3_U31 ( .A1(npu_inst_pe_1_7_3_n26), .A2(npu_inst_n34), .A3(npu_inst_int_ckg[4]), .ZN(npu_inst_pe_1_7_3_n85) );
  OR2_X1 npu_inst_pe_1_7_3_U30 ( .A1(npu_inst_pe_1_7_3_n85), .A2(
        npu_inst_pe_1_7_3_n1), .ZN(npu_inst_pe_1_7_3_N84) );
  INV_X1 npu_inst_pe_1_7_3_U29 ( .A(npu_inst_pe_1_7_3_int_data_0_), .ZN(
        npu_inst_pe_1_7_3_n12) );
  INV_X1 npu_inst_pe_1_7_3_U28 ( .A(npu_inst_n49), .ZN(npu_inst_pe_1_7_3_n4)
         );
  OR3_X1 npu_inst_pe_1_7_3_U27 ( .A1(npu_inst_pe_1_7_3_n5), .A2(
        npu_inst_pe_1_7_3_n7), .A3(npu_inst_pe_1_7_3_n4), .ZN(
        npu_inst_pe_1_7_3_n56) );
  OR3_X1 npu_inst_pe_1_7_3_U26 ( .A1(npu_inst_pe_1_7_3_n4), .A2(
        npu_inst_pe_1_7_3_n7), .A3(npu_inst_pe_1_7_3_n6), .ZN(
        npu_inst_pe_1_7_3_n48) );
  INV_X1 npu_inst_pe_1_7_3_U25 ( .A(npu_inst_pe_1_7_3_n4), .ZN(
        npu_inst_pe_1_7_3_n3) );
  OR3_X1 npu_inst_pe_1_7_3_U24 ( .A1(npu_inst_pe_1_7_3_n3), .A2(
        npu_inst_pe_1_7_3_n7), .A3(npu_inst_pe_1_7_3_n6), .ZN(
        npu_inst_pe_1_7_3_n52) );
  OR3_X1 npu_inst_pe_1_7_3_U23 ( .A1(npu_inst_pe_1_7_3_n5), .A2(
        npu_inst_pe_1_7_3_n7), .A3(npu_inst_pe_1_7_3_n3), .ZN(
        npu_inst_pe_1_7_3_n60) );
  BUF_X1 npu_inst_pe_1_7_3_U22 ( .A(npu_inst_n12), .Z(npu_inst_pe_1_7_3_n1) );
  NOR2_X1 npu_inst_pe_1_7_3_U21 ( .A1(npu_inst_pe_1_7_3_n60), .A2(
        npu_inst_pe_1_7_3_n2), .ZN(npu_inst_pe_1_7_3_n58) );
  NOR2_X1 npu_inst_pe_1_7_3_U20 ( .A1(npu_inst_pe_1_7_3_n56), .A2(
        npu_inst_pe_1_7_3_n2), .ZN(npu_inst_pe_1_7_3_n54) );
  NOR2_X1 npu_inst_pe_1_7_3_U19 ( .A1(npu_inst_pe_1_7_3_n52), .A2(
        npu_inst_pe_1_7_3_n2), .ZN(npu_inst_pe_1_7_3_n50) );
  NOR2_X1 npu_inst_pe_1_7_3_U18 ( .A1(npu_inst_pe_1_7_3_n48), .A2(
        npu_inst_pe_1_7_3_n2), .ZN(npu_inst_pe_1_7_3_n46) );
  NOR2_X1 npu_inst_pe_1_7_3_U17 ( .A1(npu_inst_pe_1_7_3_n40), .A2(
        npu_inst_pe_1_7_3_n2), .ZN(npu_inst_pe_1_7_3_n38) );
  NOR2_X1 npu_inst_pe_1_7_3_U16 ( .A1(npu_inst_pe_1_7_3_n44), .A2(
        npu_inst_pe_1_7_3_n2), .ZN(npu_inst_pe_1_7_3_n42) );
  BUF_X1 npu_inst_pe_1_7_3_U15 ( .A(npu_inst_n75), .Z(npu_inst_pe_1_7_3_n7) );
  INV_X1 npu_inst_pe_1_7_3_U14 ( .A(npu_inst_n104), .ZN(npu_inst_pe_1_7_3_n11)
         );
  INV_X1 npu_inst_pe_1_7_3_U13 ( .A(npu_inst_pe_1_7_3_n38), .ZN(
        npu_inst_pe_1_7_3_n113) );
  INV_X1 npu_inst_pe_1_7_3_U12 ( .A(npu_inst_pe_1_7_3_n58), .ZN(
        npu_inst_pe_1_7_3_n118) );
  INV_X1 npu_inst_pe_1_7_3_U11 ( .A(npu_inst_pe_1_7_3_n54), .ZN(
        npu_inst_pe_1_7_3_n117) );
  INV_X1 npu_inst_pe_1_7_3_U10 ( .A(npu_inst_pe_1_7_3_n50), .ZN(
        npu_inst_pe_1_7_3_n116) );
  INV_X1 npu_inst_pe_1_7_3_U9 ( .A(npu_inst_pe_1_7_3_n46), .ZN(
        npu_inst_pe_1_7_3_n115) );
  INV_X1 npu_inst_pe_1_7_3_U8 ( .A(npu_inst_pe_1_7_3_n42), .ZN(
        npu_inst_pe_1_7_3_n114) );
  BUF_X1 npu_inst_pe_1_7_3_U7 ( .A(npu_inst_pe_1_7_3_n11), .Z(
        npu_inst_pe_1_7_3_n10) );
  BUF_X1 npu_inst_pe_1_7_3_U6 ( .A(npu_inst_pe_1_7_3_n11), .Z(
        npu_inst_pe_1_7_3_n9) );
  BUF_X1 npu_inst_pe_1_7_3_U5 ( .A(npu_inst_pe_1_7_3_n11), .Z(
        npu_inst_pe_1_7_3_n8) );
  NOR2_X1 npu_inst_pe_1_7_3_U4 ( .A1(npu_inst_pe_1_7_3_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_3_n1), .ZN(npu_inst_pe_1_7_3_n76) );
  NOR2_X1 npu_inst_pe_1_7_3_U3 ( .A1(npu_inst_pe_1_7_3_n27), .A2(
        npu_inst_pe_1_7_3_n1), .ZN(npu_inst_pe_1_7_3_n77) );
  FA_X1 npu_inst_pe_1_7_3_sub_77_U2_1 ( .A(npu_inst_int_data_res_7__3__1_), 
        .B(npu_inst_pe_1_7_3_n13), .CI(npu_inst_pe_1_7_3_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_7_3_sub_77_carry_2_), .S(npu_inst_pe_1_7_3_N66) );
  FA_X1 npu_inst_pe_1_7_3_add_79_U1_1 ( .A(npu_inst_int_data_res_7__3__1_), 
        .B(npu_inst_pe_1_7_3_int_data_1_), .CI(
        npu_inst_pe_1_7_3_add_79_carry_1_), .CO(
        npu_inst_pe_1_7_3_add_79_carry_2_), .S(npu_inst_pe_1_7_3_N74) );
  NAND3_X1 npu_inst_pe_1_7_3_U101 ( .A1(npu_inst_pe_1_7_3_n4), .A2(
        npu_inst_pe_1_7_3_n6), .A3(npu_inst_pe_1_7_3_n7), .ZN(
        npu_inst_pe_1_7_3_n44) );
  NAND3_X1 npu_inst_pe_1_7_3_U100 ( .A1(npu_inst_pe_1_7_3_n3), .A2(
        npu_inst_pe_1_7_3_n6), .A3(npu_inst_pe_1_7_3_n7), .ZN(
        npu_inst_pe_1_7_3_n40) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_3_n33), .CK(
        npu_inst_pe_1_7_3_net3121), .RN(npu_inst_pe_1_7_3_n8), .Q(
        npu_inst_int_data_res_7__3__6_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_3_n34), .CK(
        npu_inst_pe_1_7_3_net3121), .RN(npu_inst_pe_1_7_3_n8), .Q(
        npu_inst_int_data_res_7__3__5_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_3_n35), .CK(
        npu_inst_pe_1_7_3_net3121), .RN(npu_inst_pe_1_7_3_n8), .Q(
        npu_inst_int_data_res_7__3__4_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_3_n36), .CK(
        npu_inst_pe_1_7_3_net3121), .RN(npu_inst_pe_1_7_3_n8), .Q(
        npu_inst_int_data_res_7__3__3_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_3_n98), .CK(
        npu_inst_pe_1_7_3_net3121), .RN(npu_inst_pe_1_7_3_n8), .Q(
        npu_inst_int_data_res_7__3__2_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_3_n99), .CK(
        npu_inst_pe_1_7_3_net3121), .RN(npu_inst_pe_1_7_3_n8), .Q(
        npu_inst_int_data_res_7__3__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_3_n32), .CK(
        npu_inst_pe_1_7_3_net3121), .RN(npu_inst_pe_1_7_3_n8), .Q(
        npu_inst_int_data_res_7__3__7_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_3_n100), 
        .CK(npu_inst_pe_1_7_3_net3121), .RN(npu_inst_pe_1_7_3_n8), .Q(
        npu_inst_int_data_res_7__3__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_weight_reg_0_ ( .D(npu_inst_n90), .CK(
        npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n8), .Q(
        npu_inst_pe_1_7_3_int_q_weight_0_), .QN(npu_inst_pe_1_7_3_n27) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_weight_reg_1_ ( .D(npu_inst_n96), .CK(
        npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n8), .Q(
        npu_inst_pe_1_7_3_int_q_weight_1_), .QN(npu_inst_pe_1_7_3_n26) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_3_n112), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n8), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_3_n111), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n8), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_3_n110), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_3_n109), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_3_n108), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_3_n107), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_3_n106), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_3_n105), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_3_n104), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_3_n103), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_3_n102), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_3_n101), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_3_n86), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_3_n87), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n9), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_3_n88), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_3_n89), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_3_n90), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_3_n91), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_3_n92), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_3_n93), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_3_n94), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_3_n95), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_3_n96), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_3_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_3_n97), 
        .CK(npu_inst_pe_1_7_3_net3127), .RN(npu_inst_pe_1_7_3_n10), .Q(
        npu_inst_pe_1_7_3_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_3_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_3_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_3_net3121) );
  CLKGATETST_X1 npu_inst_pe_1_7_3_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n43), .SE(1'b0), .GCK(npu_inst_pe_1_7_3_net3127) );
  MUX2_X1 npu_inst_pe_1_7_4_U153 ( .A(npu_inst_pe_1_7_4_n31), .B(
        npu_inst_pe_1_7_4_n28), .S(npu_inst_pe_1_7_4_n7), .Z(
        npu_inst_pe_1_7_4_N93) );
  MUX2_X1 npu_inst_pe_1_7_4_U152 ( .A(npu_inst_pe_1_7_4_n30), .B(
        npu_inst_pe_1_7_4_n29), .S(npu_inst_pe_1_7_4_n5), .Z(
        npu_inst_pe_1_7_4_n31) );
  MUX2_X1 npu_inst_pe_1_7_4_U151 ( .A(npu_inst_pe_1_7_4_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_4_n3), .Z(
        npu_inst_pe_1_7_4_n30) );
  MUX2_X1 npu_inst_pe_1_7_4_U150 ( .A(npu_inst_pe_1_7_4_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_4_n3), .Z(
        npu_inst_pe_1_7_4_n29) );
  MUX2_X1 npu_inst_pe_1_7_4_U149 ( .A(npu_inst_pe_1_7_4_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_4_n3), .Z(
        npu_inst_pe_1_7_4_n28) );
  MUX2_X1 npu_inst_pe_1_7_4_U148 ( .A(npu_inst_pe_1_7_4_n25), .B(
        npu_inst_pe_1_7_4_n22), .S(npu_inst_pe_1_7_4_n7), .Z(
        npu_inst_pe_1_7_4_N94) );
  MUX2_X1 npu_inst_pe_1_7_4_U147 ( .A(npu_inst_pe_1_7_4_n24), .B(
        npu_inst_pe_1_7_4_n23), .S(npu_inst_pe_1_7_4_n5), .Z(
        npu_inst_pe_1_7_4_n25) );
  MUX2_X1 npu_inst_pe_1_7_4_U146 ( .A(npu_inst_pe_1_7_4_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_4_n3), .Z(
        npu_inst_pe_1_7_4_n24) );
  MUX2_X1 npu_inst_pe_1_7_4_U145 ( .A(npu_inst_pe_1_7_4_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_4_n3), .Z(
        npu_inst_pe_1_7_4_n23) );
  MUX2_X1 npu_inst_pe_1_7_4_U144 ( .A(npu_inst_pe_1_7_4_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_4_n3), .Z(
        npu_inst_pe_1_7_4_n22) );
  MUX2_X1 npu_inst_pe_1_7_4_U143 ( .A(npu_inst_pe_1_7_4_n21), .B(
        npu_inst_pe_1_7_4_n18), .S(npu_inst_pe_1_7_4_n7), .Z(
        npu_inst_int_data_x_7__4__1_) );
  MUX2_X1 npu_inst_pe_1_7_4_U142 ( .A(npu_inst_pe_1_7_4_n20), .B(
        npu_inst_pe_1_7_4_n19), .S(npu_inst_pe_1_7_4_n5), .Z(
        npu_inst_pe_1_7_4_n21) );
  MUX2_X1 npu_inst_pe_1_7_4_U141 ( .A(npu_inst_pe_1_7_4_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_4_n3), .Z(
        npu_inst_pe_1_7_4_n20) );
  MUX2_X1 npu_inst_pe_1_7_4_U140 ( .A(npu_inst_pe_1_7_4_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_4_n3), .Z(
        npu_inst_pe_1_7_4_n19) );
  MUX2_X1 npu_inst_pe_1_7_4_U139 ( .A(npu_inst_pe_1_7_4_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_4_n3), .Z(
        npu_inst_pe_1_7_4_n18) );
  MUX2_X1 npu_inst_pe_1_7_4_U138 ( .A(npu_inst_pe_1_7_4_n17), .B(
        npu_inst_pe_1_7_4_n14), .S(npu_inst_pe_1_7_4_n7), .Z(
        npu_inst_int_data_x_7__4__0_) );
  MUX2_X1 npu_inst_pe_1_7_4_U137 ( .A(npu_inst_pe_1_7_4_n16), .B(
        npu_inst_pe_1_7_4_n15), .S(npu_inst_pe_1_7_4_n5), .Z(
        npu_inst_pe_1_7_4_n17) );
  MUX2_X1 npu_inst_pe_1_7_4_U136 ( .A(npu_inst_pe_1_7_4_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_4_n3), .Z(
        npu_inst_pe_1_7_4_n16) );
  MUX2_X1 npu_inst_pe_1_7_4_U135 ( .A(npu_inst_pe_1_7_4_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_4_n3), .Z(
        npu_inst_pe_1_7_4_n15) );
  MUX2_X1 npu_inst_pe_1_7_4_U134 ( .A(npu_inst_pe_1_7_4_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_4_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_4_n3), .Z(
        npu_inst_pe_1_7_4_n14) );
  XOR2_X1 npu_inst_pe_1_7_4_U133 ( .A(npu_inst_pe_1_7_4_int_data_0_), .B(
        npu_inst_int_data_res_7__4__0_), .Z(npu_inst_pe_1_7_4_N73) );
  AND2_X1 npu_inst_pe_1_7_4_U132 ( .A1(npu_inst_int_data_res_7__4__0_), .A2(
        npu_inst_pe_1_7_4_int_data_0_), .ZN(npu_inst_pe_1_7_4_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_4_U131 ( .A(npu_inst_int_data_res_7__4__0_), .B(
        npu_inst_pe_1_7_4_n12), .ZN(npu_inst_pe_1_7_4_N65) );
  OR2_X1 npu_inst_pe_1_7_4_U130 ( .A1(npu_inst_pe_1_7_4_n12), .A2(
        npu_inst_int_data_res_7__4__0_), .ZN(npu_inst_pe_1_7_4_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_4_U129 ( .A(npu_inst_int_data_res_7__4__2_), .B(
        npu_inst_pe_1_7_4_add_79_carry_2_), .Z(npu_inst_pe_1_7_4_N75) );
  AND2_X1 npu_inst_pe_1_7_4_U128 ( .A1(npu_inst_pe_1_7_4_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_7__4__2_), .ZN(
        npu_inst_pe_1_7_4_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_4_U127 ( .A(npu_inst_int_data_res_7__4__3_), .B(
        npu_inst_pe_1_7_4_add_79_carry_3_), .Z(npu_inst_pe_1_7_4_N76) );
  AND2_X1 npu_inst_pe_1_7_4_U126 ( .A1(npu_inst_pe_1_7_4_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_7__4__3_), .ZN(
        npu_inst_pe_1_7_4_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_4_U125 ( .A(npu_inst_int_data_res_7__4__4_), .B(
        npu_inst_pe_1_7_4_add_79_carry_4_), .Z(npu_inst_pe_1_7_4_N77) );
  AND2_X1 npu_inst_pe_1_7_4_U124 ( .A1(npu_inst_pe_1_7_4_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_7__4__4_), .ZN(
        npu_inst_pe_1_7_4_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_4_U123 ( .A(npu_inst_int_data_res_7__4__5_), .B(
        npu_inst_pe_1_7_4_add_79_carry_5_), .Z(npu_inst_pe_1_7_4_N78) );
  AND2_X1 npu_inst_pe_1_7_4_U122 ( .A1(npu_inst_pe_1_7_4_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_7__4__5_), .ZN(
        npu_inst_pe_1_7_4_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_4_U121 ( .A(npu_inst_int_data_res_7__4__6_), .B(
        npu_inst_pe_1_7_4_add_79_carry_6_), .Z(npu_inst_pe_1_7_4_N79) );
  AND2_X1 npu_inst_pe_1_7_4_U120 ( .A1(npu_inst_pe_1_7_4_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_7__4__6_), .ZN(
        npu_inst_pe_1_7_4_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_4_U119 ( .A(npu_inst_int_data_res_7__4__7_), .B(
        npu_inst_pe_1_7_4_add_79_carry_7_), .Z(npu_inst_pe_1_7_4_N80) );
  XNOR2_X1 npu_inst_pe_1_7_4_U118 ( .A(npu_inst_pe_1_7_4_sub_77_carry_2_), .B(
        npu_inst_int_data_res_7__4__2_), .ZN(npu_inst_pe_1_7_4_N67) );
  OR2_X1 npu_inst_pe_1_7_4_U117 ( .A1(npu_inst_int_data_res_7__4__2_), .A2(
        npu_inst_pe_1_7_4_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_7_4_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_4_U116 ( .A(npu_inst_pe_1_7_4_sub_77_carry_3_), .B(
        npu_inst_int_data_res_7__4__3_), .ZN(npu_inst_pe_1_7_4_N68) );
  OR2_X1 npu_inst_pe_1_7_4_U115 ( .A1(npu_inst_int_data_res_7__4__3_), .A2(
        npu_inst_pe_1_7_4_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_7_4_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_4_U114 ( .A(npu_inst_pe_1_7_4_sub_77_carry_4_), .B(
        npu_inst_int_data_res_7__4__4_), .ZN(npu_inst_pe_1_7_4_N69) );
  OR2_X1 npu_inst_pe_1_7_4_U113 ( .A1(npu_inst_int_data_res_7__4__4_), .A2(
        npu_inst_pe_1_7_4_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_7_4_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_4_U112 ( .A(npu_inst_pe_1_7_4_sub_77_carry_5_), .B(
        npu_inst_int_data_res_7__4__5_), .ZN(npu_inst_pe_1_7_4_N70) );
  OR2_X1 npu_inst_pe_1_7_4_U111 ( .A1(npu_inst_int_data_res_7__4__5_), .A2(
        npu_inst_pe_1_7_4_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_7_4_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_4_U110 ( .A(npu_inst_pe_1_7_4_sub_77_carry_6_), .B(
        npu_inst_int_data_res_7__4__6_), .ZN(npu_inst_pe_1_7_4_N71) );
  OR2_X1 npu_inst_pe_1_7_4_U109 ( .A1(npu_inst_int_data_res_7__4__6_), .A2(
        npu_inst_pe_1_7_4_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_7_4_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_4_U108 ( .A(npu_inst_int_data_res_7__4__7_), .B(
        npu_inst_pe_1_7_4_sub_77_carry_7_), .ZN(npu_inst_pe_1_7_4_N72) );
  INV_X1 npu_inst_pe_1_7_4_U107 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_7_4_n6)
         );
  INV_X1 npu_inst_pe_1_7_4_U106 ( .A(npu_inst_pe_1_7_4_n6), .ZN(
        npu_inst_pe_1_7_4_n5) );
  INV_X1 npu_inst_pe_1_7_4_U105 ( .A(npu_inst_n34), .ZN(npu_inst_pe_1_7_4_n2)
         );
  AOI22_X1 npu_inst_pe_1_7_4_U104 ( .A1(npu_inst_pe_1_7_4_n38), .A2(
        int_i_data_v_npu[7]), .B1(npu_inst_pe_1_7_4_n113), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_4_n39) );
  INV_X1 npu_inst_pe_1_7_4_U103 ( .A(npu_inst_pe_1_7_4_n39), .ZN(
        npu_inst_pe_1_7_4_n111) );
  AOI22_X1 npu_inst_pe_1_7_4_U102 ( .A1(npu_inst_pe_1_7_4_n38), .A2(
        int_i_data_v_npu[6]), .B1(npu_inst_pe_1_7_4_n113), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_4_n37) );
  INV_X1 npu_inst_pe_1_7_4_U99 ( .A(npu_inst_pe_1_7_4_n37), .ZN(
        npu_inst_pe_1_7_4_n112) );
  AOI22_X1 npu_inst_pe_1_7_4_U98 ( .A1(int_i_data_v_npu[7]), .A2(
        npu_inst_pe_1_7_4_n58), .B1(npu_inst_pe_1_7_4_n118), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_4_n59) );
  INV_X1 npu_inst_pe_1_7_4_U97 ( .A(npu_inst_pe_1_7_4_n59), .ZN(
        npu_inst_pe_1_7_4_n101) );
  AOI22_X1 npu_inst_pe_1_7_4_U96 ( .A1(int_i_data_v_npu[6]), .A2(
        npu_inst_pe_1_7_4_n58), .B1(npu_inst_pe_1_7_4_n118), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_4_n57) );
  INV_X1 npu_inst_pe_1_7_4_U95 ( .A(npu_inst_pe_1_7_4_n57), .ZN(
        npu_inst_pe_1_7_4_n102) );
  AOI22_X1 npu_inst_pe_1_7_4_U94 ( .A1(int_i_data_v_npu[7]), .A2(
        npu_inst_pe_1_7_4_n54), .B1(npu_inst_pe_1_7_4_n117), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_4_n55) );
  INV_X1 npu_inst_pe_1_7_4_U93 ( .A(npu_inst_pe_1_7_4_n55), .ZN(
        npu_inst_pe_1_7_4_n103) );
  AOI22_X1 npu_inst_pe_1_7_4_U92 ( .A1(int_i_data_v_npu[6]), .A2(
        npu_inst_pe_1_7_4_n54), .B1(npu_inst_pe_1_7_4_n117), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_4_n53) );
  INV_X1 npu_inst_pe_1_7_4_U91 ( .A(npu_inst_pe_1_7_4_n53), .ZN(
        npu_inst_pe_1_7_4_n104) );
  AOI22_X1 npu_inst_pe_1_7_4_U90 ( .A1(int_i_data_v_npu[7]), .A2(
        npu_inst_pe_1_7_4_n50), .B1(npu_inst_pe_1_7_4_n116), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_4_n51) );
  INV_X1 npu_inst_pe_1_7_4_U89 ( .A(npu_inst_pe_1_7_4_n51), .ZN(
        npu_inst_pe_1_7_4_n105) );
  AOI22_X1 npu_inst_pe_1_7_4_U88 ( .A1(int_i_data_v_npu[6]), .A2(
        npu_inst_pe_1_7_4_n50), .B1(npu_inst_pe_1_7_4_n116), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_4_n49) );
  INV_X1 npu_inst_pe_1_7_4_U87 ( .A(npu_inst_pe_1_7_4_n49), .ZN(
        npu_inst_pe_1_7_4_n106) );
  AOI22_X1 npu_inst_pe_1_7_4_U86 ( .A1(int_i_data_v_npu[7]), .A2(
        npu_inst_pe_1_7_4_n46), .B1(npu_inst_pe_1_7_4_n115), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_4_n47) );
  INV_X1 npu_inst_pe_1_7_4_U85 ( .A(npu_inst_pe_1_7_4_n47), .ZN(
        npu_inst_pe_1_7_4_n107) );
  AOI22_X1 npu_inst_pe_1_7_4_U84 ( .A1(int_i_data_v_npu[6]), .A2(
        npu_inst_pe_1_7_4_n46), .B1(npu_inst_pe_1_7_4_n115), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_4_n45) );
  INV_X1 npu_inst_pe_1_7_4_U83 ( .A(npu_inst_pe_1_7_4_n45), .ZN(
        npu_inst_pe_1_7_4_n108) );
  AOI22_X1 npu_inst_pe_1_7_4_U82 ( .A1(int_i_data_v_npu[7]), .A2(
        npu_inst_pe_1_7_4_n42), .B1(npu_inst_pe_1_7_4_n114), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_4_n43) );
  INV_X1 npu_inst_pe_1_7_4_U81 ( .A(npu_inst_pe_1_7_4_n43), .ZN(
        npu_inst_pe_1_7_4_n109) );
  AOI22_X1 npu_inst_pe_1_7_4_U80 ( .A1(int_i_data_v_npu[6]), .A2(
        npu_inst_pe_1_7_4_n42), .B1(npu_inst_pe_1_7_4_n114), .B2(
        npu_inst_pe_1_7_4_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_4_n41) );
  INV_X1 npu_inst_pe_1_7_4_U79 ( .A(npu_inst_pe_1_7_4_n41), .ZN(
        npu_inst_pe_1_7_4_n110) );
  AND2_X1 npu_inst_pe_1_7_4_U78 ( .A1(npu_inst_pe_1_7_4_N93), .A2(npu_inst_n34), .ZN(npu_inst_int_data_y_7__4__0_) );
  NAND2_X1 npu_inst_pe_1_7_4_U77 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_4_n60), .ZN(npu_inst_pe_1_7_4_n74) );
  OAI21_X1 npu_inst_pe_1_7_4_U76 ( .B1(npu_inst_pe_1_7_4_n63), .B2(
        npu_inst_pe_1_7_4_n60), .A(npu_inst_pe_1_7_4_n74), .ZN(
        npu_inst_pe_1_7_4_n97) );
  NAND2_X1 npu_inst_pe_1_7_4_U75 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_4_n60), .ZN(npu_inst_pe_1_7_4_n73) );
  OAI21_X1 npu_inst_pe_1_7_4_U74 ( .B1(npu_inst_pe_1_7_4_n61), .B2(
        npu_inst_pe_1_7_4_n60), .A(npu_inst_pe_1_7_4_n73), .ZN(
        npu_inst_pe_1_7_4_n96) );
  NAND2_X1 npu_inst_pe_1_7_4_U73 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_4_n56), .ZN(npu_inst_pe_1_7_4_n72) );
  OAI21_X1 npu_inst_pe_1_7_4_U72 ( .B1(npu_inst_pe_1_7_4_n63), .B2(
        npu_inst_pe_1_7_4_n56), .A(npu_inst_pe_1_7_4_n72), .ZN(
        npu_inst_pe_1_7_4_n95) );
  NAND2_X1 npu_inst_pe_1_7_4_U71 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_4_n56), .ZN(npu_inst_pe_1_7_4_n71) );
  OAI21_X1 npu_inst_pe_1_7_4_U70 ( .B1(npu_inst_pe_1_7_4_n61), .B2(
        npu_inst_pe_1_7_4_n56), .A(npu_inst_pe_1_7_4_n71), .ZN(
        npu_inst_pe_1_7_4_n94) );
  NAND2_X1 npu_inst_pe_1_7_4_U69 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_4_n52), .ZN(npu_inst_pe_1_7_4_n70) );
  OAI21_X1 npu_inst_pe_1_7_4_U68 ( .B1(npu_inst_pe_1_7_4_n63), .B2(
        npu_inst_pe_1_7_4_n52), .A(npu_inst_pe_1_7_4_n70), .ZN(
        npu_inst_pe_1_7_4_n93) );
  NAND2_X1 npu_inst_pe_1_7_4_U67 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_4_n52), .ZN(npu_inst_pe_1_7_4_n69) );
  OAI21_X1 npu_inst_pe_1_7_4_U66 ( .B1(npu_inst_pe_1_7_4_n61), .B2(
        npu_inst_pe_1_7_4_n52), .A(npu_inst_pe_1_7_4_n69), .ZN(
        npu_inst_pe_1_7_4_n92) );
  NAND2_X1 npu_inst_pe_1_7_4_U65 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_4_n48), .ZN(npu_inst_pe_1_7_4_n68) );
  OAI21_X1 npu_inst_pe_1_7_4_U64 ( .B1(npu_inst_pe_1_7_4_n63), .B2(
        npu_inst_pe_1_7_4_n48), .A(npu_inst_pe_1_7_4_n68), .ZN(
        npu_inst_pe_1_7_4_n91) );
  NAND2_X1 npu_inst_pe_1_7_4_U63 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_4_n48), .ZN(npu_inst_pe_1_7_4_n67) );
  OAI21_X1 npu_inst_pe_1_7_4_U62 ( .B1(npu_inst_pe_1_7_4_n61), .B2(
        npu_inst_pe_1_7_4_n48), .A(npu_inst_pe_1_7_4_n67), .ZN(
        npu_inst_pe_1_7_4_n90) );
  NAND2_X1 npu_inst_pe_1_7_4_U61 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_4_n44), .ZN(npu_inst_pe_1_7_4_n66) );
  OAI21_X1 npu_inst_pe_1_7_4_U60 ( .B1(npu_inst_pe_1_7_4_n63), .B2(
        npu_inst_pe_1_7_4_n44), .A(npu_inst_pe_1_7_4_n66), .ZN(
        npu_inst_pe_1_7_4_n89) );
  NAND2_X1 npu_inst_pe_1_7_4_U59 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_4_n44), .ZN(npu_inst_pe_1_7_4_n65) );
  OAI21_X1 npu_inst_pe_1_7_4_U58 ( .B1(npu_inst_pe_1_7_4_n61), .B2(
        npu_inst_pe_1_7_4_n44), .A(npu_inst_pe_1_7_4_n65), .ZN(
        npu_inst_pe_1_7_4_n88) );
  NAND2_X1 npu_inst_pe_1_7_4_U57 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_4_n40), .ZN(npu_inst_pe_1_7_4_n64) );
  OAI21_X1 npu_inst_pe_1_7_4_U56 ( .B1(npu_inst_pe_1_7_4_n63), .B2(
        npu_inst_pe_1_7_4_n40), .A(npu_inst_pe_1_7_4_n64), .ZN(
        npu_inst_pe_1_7_4_n87) );
  NAND2_X1 npu_inst_pe_1_7_4_U55 ( .A1(npu_inst_pe_1_7_4_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_4_n40), .ZN(npu_inst_pe_1_7_4_n62) );
  OAI21_X1 npu_inst_pe_1_7_4_U54 ( .B1(npu_inst_pe_1_7_4_n61), .B2(
        npu_inst_pe_1_7_4_n40), .A(npu_inst_pe_1_7_4_n62), .ZN(
        npu_inst_pe_1_7_4_n86) );
  AND2_X1 npu_inst_pe_1_7_4_U53 ( .A1(npu_inst_n34), .A2(npu_inst_pe_1_7_4_N94), .ZN(npu_inst_int_data_y_7__4__1_) );
  AOI22_X1 npu_inst_pe_1_7_4_U52 ( .A1(npu_inst_n34), .A2(int_i_data_v_npu[7]), 
        .B1(npu_inst_pe_1_7_4_n2), .B2(npu_inst_int_data_x_7__5__1_), .ZN(
        npu_inst_pe_1_7_4_n63) );
  AOI22_X1 npu_inst_pe_1_7_4_U51 ( .A1(npu_inst_n34), .A2(int_i_data_v_npu[6]), 
        .B1(npu_inst_pe_1_7_4_n2), .B2(npu_inst_int_data_x_7__5__0_), .ZN(
        npu_inst_pe_1_7_4_n61) );
  AOI222_X1 npu_inst_pe_1_7_4_U50 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N73), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N65), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n84) );
  INV_X1 npu_inst_pe_1_7_4_U49 ( .A(npu_inst_pe_1_7_4_n84), .ZN(
        npu_inst_pe_1_7_4_n100) );
  AOI222_X1 npu_inst_pe_1_7_4_U48 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N74), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N66), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n83) );
  INV_X1 npu_inst_pe_1_7_4_U47 ( .A(npu_inst_pe_1_7_4_n83), .ZN(
        npu_inst_pe_1_7_4_n99) );
  AOI222_X1 npu_inst_pe_1_7_4_U46 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N75), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N67), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n82) );
  INV_X1 npu_inst_pe_1_7_4_U45 ( .A(npu_inst_pe_1_7_4_n82), .ZN(
        npu_inst_pe_1_7_4_n98) );
  AOI222_X1 npu_inst_pe_1_7_4_U44 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N76), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N68), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n81) );
  INV_X1 npu_inst_pe_1_7_4_U43 ( .A(npu_inst_pe_1_7_4_n81), .ZN(
        npu_inst_pe_1_7_4_n36) );
  AOI222_X1 npu_inst_pe_1_7_4_U42 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N77), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N69), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n80) );
  INV_X1 npu_inst_pe_1_7_4_U41 ( .A(npu_inst_pe_1_7_4_n80), .ZN(
        npu_inst_pe_1_7_4_n35) );
  AOI222_X1 npu_inst_pe_1_7_4_U40 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N78), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N70), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n79) );
  INV_X1 npu_inst_pe_1_7_4_U39 ( .A(npu_inst_pe_1_7_4_n79), .ZN(
        npu_inst_pe_1_7_4_n34) );
  AOI222_X1 npu_inst_pe_1_7_4_U38 ( .A1(1'b0), .A2(npu_inst_pe_1_7_4_n1), .B1(
        npu_inst_pe_1_7_4_N79), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N71), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n78) );
  INV_X1 npu_inst_pe_1_7_4_U37 ( .A(npu_inst_pe_1_7_4_n78), .ZN(
        npu_inst_pe_1_7_4_n33) );
  AOI222_X1 npu_inst_pe_1_7_4_U36 ( .A1(npu_inst_pe_1_7_4_n1), .A2(1'b0), .B1(
        npu_inst_pe_1_7_4_N80), .B2(npu_inst_pe_1_7_4_n76), .C1(
        npu_inst_pe_1_7_4_N72), .C2(npu_inst_pe_1_7_4_n77), .ZN(
        npu_inst_pe_1_7_4_n75) );
  INV_X1 npu_inst_pe_1_7_4_U35 ( .A(npu_inst_pe_1_7_4_n75), .ZN(
        npu_inst_pe_1_7_4_n32) );
  AND2_X1 npu_inst_pe_1_7_4_U34 ( .A1(npu_inst_int_data_x_7__4__1_), .A2(
        npu_inst_pe_1_7_4_int_q_weight_1_), .ZN(npu_inst_pe_1_7_4_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_4_U33 ( .A1(npu_inst_int_data_x_7__4__0_), .A2(
        npu_inst_pe_1_7_4_int_q_weight_1_), .ZN(npu_inst_pe_1_7_4_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_4_U32 ( .A(npu_inst_pe_1_7_4_int_data_1_), .ZN(
        npu_inst_pe_1_7_4_n13) );
  NOR3_X1 npu_inst_pe_1_7_4_U31 ( .A1(npu_inst_pe_1_7_4_n26), .A2(npu_inst_n34), .A3(npu_inst_int_ckg[3]), .ZN(npu_inst_pe_1_7_4_n85) );
  OR2_X1 npu_inst_pe_1_7_4_U30 ( .A1(npu_inst_pe_1_7_4_n85), .A2(
        npu_inst_pe_1_7_4_n1), .ZN(npu_inst_pe_1_7_4_N84) );
  INV_X1 npu_inst_pe_1_7_4_U29 ( .A(npu_inst_pe_1_7_4_int_data_0_), .ZN(
        npu_inst_pe_1_7_4_n12) );
  INV_X1 npu_inst_pe_1_7_4_U28 ( .A(npu_inst_n49), .ZN(npu_inst_pe_1_7_4_n4)
         );
  OR3_X1 npu_inst_pe_1_7_4_U27 ( .A1(npu_inst_pe_1_7_4_n5), .A2(
        npu_inst_pe_1_7_4_n7), .A3(npu_inst_pe_1_7_4_n4), .ZN(
        npu_inst_pe_1_7_4_n56) );
  OR3_X1 npu_inst_pe_1_7_4_U26 ( .A1(npu_inst_pe_1_7_4_n4), .A2(
        npu_inst_pe_1_7_4_n7), .A3(npu_inst_pe_1_7_4_n6), .ZN(
        npu_inst_pe_1_7_4_n48) );
  INV_X1 npu_inst_pe_1_7_4_U25 ( .A(npu_inst_pe_1_7_4_n4), .ZN(
        npu_inst_pe_1_7_4_n3) );
  OR3_X1 npu_inst_pe_1_7_4_U24 ( .A1(npu_inst_pe_1_7_4_n3), .A2(
        npu_inst_pe_1_7_4_n7), .A3(npu_inst_pe_1_7_4_n6), .ZN(
        npu_inst_pe_1_7_4_n52) );
  OR3_X1 npu_inst_pe_1_7_4_U23 ( .A1(npu_inst_pe_1_7_4_n5), .A2(
        npu_inst_pe_1_7_4_n7), .A3(npu_inst_pe_1_7_4_n3), .ZN(
        npu_inst_pe_1_7_4_n60) );
  BUF_X1 npu_inst_pe_1_7_4_U22 ( .A(npu_inst_n12), .Z(npu_inst_pe_1_7_4_n1) );
  NOR2_X1 npu_inst_pe_1_7_4_U21 ( .A1(npu_inst_pe_1_7_4_n60), .A2(
        npu_inst_pe_1_7_4_n2), .ZN(npu_inst_pe_1_7_4_n58) );
  NOR2_X1 npu_inst_pe_1_7_4_U20 ( .A1(npu_inst_pe_1_7_4_n56), .A2(
        npu_inst_pe_1_7_4_n2), .ZN(npu_inst_pe_1_7_4_n54) );
  NOR2_X1 npu_inst_pe_1_7_4_U19 ( .A1(npu_inst_pe_1_7_4_n52), .A2(
        npu_inst_pe_1_7_4_n2), .ZN(npu_inst_pe_1_7_4_n50) );
  NOR2_X1 npu_inst_pe_1_7_4_U18 ( .A1(npu_inst_pe_1_7_4_n48), .A2(
        npu_inst_pe_1_7_4_n2), .ZN(npu_inst_pe_1_7_4_n46) );
  NOR2_X1 npu_inst_pe_1_7_4_U17 ( .A1(npu_inst_pe_1_7_4_n40), .A2(
        npu_inst_pe_1_7_4_n2), .ZN(npu_inst_pe_1_7_4_n38) );
  NOR2_X1 npu_inst_pe_1_7_4_U16 ( .A1(npu_inst_pe_1_7_4_n44), .A2(
        npu_inst_pe_1_7_4_n2), .ZN(npu_inst_pe_1_7_4_n42) );
  BUF_X1 npu_inst_pe_1_7_4_U15 ( .A(npu_inst_n74), .Z(npu_inst_pe_1_7_4_n7) );
  INV_X1 npu_inst_pe_1_7_4_U14 ( .A(npu_inst_n104), .ZN(npu_inst_pe_1_7_4_n11)
         );
  INV_X1 npu_inst_pe_1_7_4_U13 ( .A(npu_inst_pe_1_7_4_n38), .ZN(
        npu_inst_pe_1_7_4_n113) );
  INV_X1 npu_inst_pe_1_7_4_U12 ( .A(npu_inst_pe_1_7_4_n58), .ZN(
        npu_inst_pe_1_7_4_n118) );
  INV_X1 npu_inst_pe_1_7_4_U11 ( .A(npu_inst_pe_1_7_4_n54), .ZN(
        npu_inst_pe_1_7_4_n117) );
  INV_X1 npu_inst_pe_1_7_4_U10 ( .A(npu_inst_pe_1_7_4_n50), .ZN(
        npu_inst_pe_1_7_4_n116) );
  INV_X1 npu_inst_pe_1_7_4_U9 ( .A(npu_inst_pe_1_7_4_n46), .ZN(
        npu_inst_pe_1_7_4_n115) );
  INV_X1 npu_inst_pe_1_7_4_U8 ( .A(npu_inst_pe_1_7_4_n42), .ZN(
        npu_inst_pe_1_7_4_n114) );
  BUF_X1 npu_inst_pe_1_7_4_U7 ( .A(npu_inst_pe_1_7_4_n11), .Z(
        npu_inst_pe_1_7_4_n10) );
  BUF_X1 npu_inst_pe_1_7_4_U6 ( .A(npu_inst_pe_1_7_4_n11), .Z(
        npu_inst_pe_1_7_4_n9) );
  BUF_X1 npu_inst_pe_1_7_4_U5 ( .A(npu_inst_pe_1_7_4_n11), .Z(
        npu_inst_pe_1_7_4_n8) );
  NOR2_X1 npu_inst_pe_1_7_4_U4 ( .A1(npu_inst_pe_1_7_4_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_4_n1), .ZN(npu_inst_pe_1_7_4_n76) );
  NOR2_X1 npu_inst_pe_1_7_4_U3 ( .A1(npu_inst_pe_1_7_4_n27), .A2(
        npu_inst_pe_1_7_4_n1), .ZN(npu_inst_pe_1_7_4_n77) );
  FA_X1 npu_inst_pe_1_7_4_sub_77_U2_1 ( .A(npu_inst_int_data_res_7__4__1_), 
        .B(npu_inst_pe_1_7_4_n13), .CI(npu_inst_pe_1_7_4_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_7_4_sub_77_carry_2_), .S(npu_inst_pe_1_7_4_N66) );
  FA_X1 npu_inst_pe_1_7_4_add_79_U1_1 ( .A(npu_inst_int_data_res_7__4__1_), 
        .B(npu_inst_pe_1_7_4_int_data_1_), .CI(
        npu_inst_pe_1_7_4_add_79_carry_1_), .CO(
        npu_inst_pe_1_7_4_add_79_carry_2_), .S(npu_inst_pe_1_7_4_N74) );
  NAND3_X1 npu_inst_pe_1_7_4_U101 ( .A1(npu_inst_pe_1_7_4_n4), .A2(
        npu_inst_pe_1_7_4_n6), .A3(npu_inst_pe_1_7_4_n7), .ZN(
        npu_inst_pe_1_7_4_n44) );
  NAND3_X1 npu_inst_pe_1_7_4_U100 ( .A1(npu_inst_pe_1_7_4_n3), .A2(
        npu_inst_pe_1_7_4_n6), .A3(npu_inst_pe_1_7_4_n7), .ZN(
        npu_inst_pe_1_7_4_n40) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_4_n33), .CK(
        npu_inst_pe_1_7_4_net3098), .RN(npu_inst_pe_1_7_4_n8), .Q(
        npu_inst_int_data_res_7__4__6_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_4_n34), .CK(
        npu_inst_pe_1_7_4_net3098), .RN(npu_inst_pe_1_7_4_n8), .Q(
        npu_inst_int_data_res_7__4__5_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_4_n35), .CK(
        npu_inst_pe_1_7_4_net3098), .RN(npu_inst_pe_1_7_4_n8), .Q(
        npu_inst_int_data_res_7__4__4_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_4_n36), .CK(
        npu_inst_pe_1_7_4_net3098), .RN(npu_inst_pe_1_7_4_n8), .Q(
        npu_inst_int_data_res_7__4__3_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_4_n98), .CK(
        npu_inst_pe_1_7_4_net3098), .RN(npu_inst_pe_1_7_4_n8), .Q(
        npu_inst_int_data_res_7__4__2_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_4_n99), .CK(
        npu_inst_pe_1_7_4_net3098), .RN(npu_inst_pe_1_7_4_n8), .Q(
        npu_inst_int_data_res_7__4__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_4_n32), .CK(
        npu_inst_pe_1_7_4_net3098), .RN(npu_inst_pe_1_7_4_n8), .Q(
        npu_inst_int_data_res_7__4__7_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_4_n100), 
        .CK(npu_inst_pe_1_7_4_net3098), .RN(npu_inst_pe_1_7_4_n8), .Q(
        npu_inst_int_data_res_7__4__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_weight_reg_0_ ( .D(npu_inst_n90), .CK(
        npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n8), .Q(
        npu_inst_pe_1_7_4_int_q_weight_0_), .QN(npu_inst_pe_1_7_4_n27) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_weight_reg_1_ ( .D(npu_inst_n96), .CK(
        npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n8), .Q(
        npu_inst_pe_1_7_4_int_q_weight_1_), .QN(npu_inst_pe_1_7_4_n26) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_4_n112), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n8), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_4_n111), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n8), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_4_n110), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_4_n109), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_4_n108), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_4_n107), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_4_n106), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_4_n105), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_4_n104), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_4_n103), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_4_n102), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_4_n101), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_4_n86), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_4_n87), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n9), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_4_n88), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_4_n89), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_4_n90), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_4_n91), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_4_n92), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_4_n93), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_4_n94), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_4_n95), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_4_n96), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_4_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_4_n97), 
        .CK(npu_inst_pe_1_7_4_net3104), .RN(npu_inst_pe_1_7_4_n10), .Q(
        npu_inst_pe_1_7_4_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_4_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_4_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_4_net3098) );
  CLKGATETST_X1 npu_inst_pe_1_7_4_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n43), .SE(1'b0), .GCK(npu_inst_pe_1_7_4_net3104) );
  MUX2_X1 npu_inst_pe_1_7_5_U153 ( .A(npu_inst_pe_1_7_5_n31), .B(
        npu_inst_pe_1_7_5_n28), .S(npu_inst_pe_1_7_5_n7), .Z(
        npu_inst_pe_1_7_5_N93) );
  MUX2_X1 npu_inst_pe_1_7_5_U152 ( .A(npu_inst_pe_1_7_5_n30), .B(
        npu_inst_pe_1_7_5_n29), .S(npu_inst_pe_1_7_5_n5), .Z(
        npu_inst_pe_1_7_5_n31) );
  MUX2_X1 npu_inst_pe_1_7_5_U151 ( .A(npu_inst_pe_1_7_5_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_5_n3), .Z(
        npu_inst_pe_1_7_5_n30) );
  MUX2_X1 npu_inst_pe_1_7_5_U150 ( .A(npu_inst_pe_1_7_5_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_5_n3), .Z(
        npu_inst_pe_1_7_5_n29) );
  MUX2_X1 npu_inst_pe_1_7_5_U149 ( .A(npu_inst_pe_1_7_5_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_5_n3), .Z(
        npu_inst_pe_1_7_5_n28) );
  MUX2_X1 npu_inst_pe_1_7_5_U148 ( .A(npu_inst_pe_1_7_5_n25), .B(
        npu_inst_pe_1_7_5_n22), .S(npu_inst_pe_1_7_5_n7), .Z(
        npu_inst_pe_1_7_5_N94) );
  MUX2_X1 npu_inst_pe_1_7_5_U147 ( .A(npu_inst_pe_1_7_5_n24), .B(
        npu_inst_pe_1_7_5_n23), .S(npu_inst_pe_1_7_5_n5), .Z(
        npu_inst_pe_1_7_5_n25) );
  MUX2_X1 npu_inst_pe_1_7_5_U146 ( .A(npu_inst_pe_1_7_5_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_5_n3), .Z(
        npu_inst_pe_1_7_5_n24) );
  MUX2_X1 npu_inst_pe_1_7_5_U145 ( .A(npu_inst_pe_1_7_5_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_5_n3), .Z(
        npu_inst_pe_1_7_5_n23) );
  MUX2_X1 npu_inst_pe_1_7_5_U144 ( .A(npu_inst_pe_1_7_5_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_5_n3), .Z(
        npu_inst_pe_1_7_5_n22) );
  MUX2_X1 npu_inst_pe_1_7_5_U143 ( .A(npu_inst_pe_1_7_5_n21), .B(
        npu_inst_pe_1_7_5_n18), .S(npu_inst_pe_1_7_5_n7), .Z(
        npu_inst_int_data_x_7__5__1_) );
  MUX2_X1 npu_inst_pe_1_7_5_U142 ( .A(npu_inst_pe_1_7_5_n20), .B(
        npu_inst_pe_1_7_5_n19), .S(npu_inst_pe_1_7_5_n5), .Z(
        npu_inst_pe_1_7_5_n21) );
  MUX2_X1 npu_inst_pe_1_7_5_U141 ( .A(npu_inst_pe_1_7_5_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_5_n3), .Z(
        npu_inst_pe_1_7_5_n20) );
  MUX2_X1 npu_inst_pe_1_7_5_U140 ( .A(npu_inst_pe_1_7_5_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_5_n3), .Z(
        npu_inst_pe_1_7_5_n19) );
  MUX2_X1 npu_inst_pe_1_7_5_U139 ( .A(npu_inst_pe_1_7_5_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_5_n3), .Z(
        npu_inst_pe_1_7_5_n18) );
  MUX2_X1 npu_inst_pe_1_7_5_U138 ( .A(npu_inst_pe_1_7_5_n17), .B(
        npu_inst_pe_1_7_5_n14), .S(npu_inst_pe_1_7_5_n7), .Z(
        npu_inst_int_data_x_7__5__0_) );
  MUX2_X1 npu_inst_pe_1_7_5_U137 ( .A(npu_inst_pe_1_7_5_n16), .B(
        npu_inst_pe_1_7_5_n15), .S(npu_inst_pe_1_7_5_n5), .Z(
        npu_inst_pe_1_7_5_n17) );
  MUX2_X1 npu_inst_pe_1_7_5_U136 ( .A(npu_inst_pe_1_7_5_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_5_n3), .Z(
        npu_inst_pe_1_7_5_n16) );
  MUX2_X1 npu_inst_pe_1_7_5_U135 ( .A(npu_inst_pe_1_7_5_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_5_n3), .Z(
        npu_inst_pe_1_7_5_n15) );
  MUX2_X1 npu_inst_pe_1_7_5_U134 ( .A(npu_inst_pe_1_7_5_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_5_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_5_n3), .Z(
        npu_inst_pe_1_7_5_n14) );
  XOR2_X1 npu_inst_pe_1_7_5_U133 ( .A(npu_inst_pe_1_7_5_int_data_0_), .B(
        npu_inst_int_data_res_7__5__0_), .Z(npu_inst_pe_1_7_5_N73) );
  AND2_X1 npu_inst_pe_1_7_5_U132 ( .A1(npu_inst_int_data_res_7__5__0_), .A2(
        npu_inst_pe_1_7_5_int_data_0_), .ZN(npu_inst_pe_1_7_5_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_5_U131 ( .A(npu_inst_int_data_res_7__5__0_), .B(
        npu_inst_pe_1_7_5_n12), .ZN(npu_inst_pe_1_7_5_N65) );
  OR2_X1 npu_inst_pe_1_7_5_U130 ( .A1(npu_inst_pe_1_7_5_n12), .A2(
        npu_inst_int_data_res_7__5__0_), .ZN(npu_inst_pe_1_7_5_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_5_U129 ( .A(npu_inst_int_data_res_7__5__2_), .B(
        npu_inst_pe_1_7_5_add_79_carry_2_), .Z(npu_inst_pe_1_7_5_N75) );
  AND2_X1 npu_inst_pe_1_7_5_U128 ( .A1(npu_inst_pe_1_7_5_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_7__5__2_), .ZN(
        npu_inst_pe_1_7_5_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_5_U127 ( .A(npu_inst_int_data_res_7__5__3_), .B(
        npu_inst_pe_1_7_5_add_79_carry_3_), .Z(npu_inst_pe_1_7_5_N76) );
  AND2_X1 npu_inst_pe_1_7_5_U126 ( .A1(npu_inst_pe_1_7_5_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_7__5__3_), .ZN(
        npu_inst_pe_1_7_5_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_5_U125 ( .A(npu_inst_int_data_res_7__5__4_), .B(
        npu_inst_pe_1_7_5_add_79_carry_4_), .Z(npu_inst_pe_1_7_5_N77) );
  AND2_X1 npu_inst_pe_1_7_5_U124 ( .A1(npu_inst_pe_1_7_5_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_7__5__4_), .ZN(
        npu_inst_pe_1_7_5_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_5_U123 ( .A(npu_inst_int_data_res_7__5__5_), .B(
        npu_inst_pe_1_7_5_add_79_carry_5_), .Z(npu_inst_pe_1_7_5_N78) );
  AND2_X1 npu_inst_pe_1_7_5_U122 ( .A1(npu_inst_pe_1_7_5_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_7__5__5_), .ZN(
        npu_inst_pe_1_7_5_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_5_U121 ( .A(npu_inst_int_data_res_7__5__6_), .B(
        npu_inst_pe_1_7_5_add_79_carry_6_), .Z(npu_inst_pe_1_7_5_N79) );
  AND2_X1 npu_inst_pe_1_7_5_U120 ( .A1(npu_inst_pe_1_7_5_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_7__5__6_), .ZN(
        npu_inst_pe_1_7_5_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_5_U119 ( .A(npu_inst_int_data_res_7__5__7_), .B(
        npu_inst_pe_1_7_5_add_79_carry_7_), .Z(npu_inst_pe_1_7_5_N80) );
  XNOR2_X1 npu_inst_pe_1_7_5_U118 ( .A(npu_inst_pe_1_7_5_sub_77_carry_2_), .B(
        npu_inst_int_data_res_7__5__2_), .ZN(npu_inst_pe_1_7_5_N67) );
  OR2_X1 npu_inst_pe_1_7_5_U117 ( .A1(npu_inst_int_data_res_7__5__2_), .A2(
        npu_inst_pe_1_7_5_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_7_5_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_5_U116 ( .A(npu_inst_pe_1_7_5_sub_77_carry_3_), .B(
        npu_inst_int_data_res_7__5__3_), .ZN(npu_inst_pe_1_7_5_N68) );
  OR2_X1 npu_inst_pe_1_7_5_U115 ( .A1(npu_inst_int_data_res_7__5__3_), .A2(
        npu_inst_pe_1_7_5_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_7_5_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_5_U114 ( .A(npu_inst_pe_1_7_5_sub_77_carry_4_), .B(
        npu_inst_int_data_res_7__5__4_), .ZN(npu_inst_pe_1_7_5_N69) );
  OR2_X1 npu_inst_pe_1_7_5_U113 ( .A1(npu_inst_int_data_res_7__5__4_), .A2(
        npu_inst_pe_1_7_5_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_7_5_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_5_U112 ( .A(npu_inst_pe_1_7_5_sub_77_carry_5_), .B(
        npu_inst_int_data_res_7__5__5_), .ZN(npu_inst_pe_1_7_5_N70) );
  OR2_X1 npu_inst_pe_1_7_5_U111 ( .A1(npu_inst_int_data_res_7__5__5_), .A2(
        npu_inst_pe_1_7_5_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_7_5_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_5_U110 ( .A(npu_inst_pe_1_7_5_sub_77_carry_6_), .B(
        npu_inst_int_data_res_7__5__6_), .ZN(npu_inst_pe_1_7_5_N71) );
  OR2_X1 npu_inst_pe_1_7_5_U109 ( .A1(npu_inst_int_data_res_7__5__6_), .A2(
        npu_inst_pe_1_7_5_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_7_5_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_5_U108 ( .A(npu_inst_int_data_res_7__5__7_), .B(
        npu_inst_pe_1_7_5_sub_77_carry_7_), .ZN(npu_inst_pe_1_7_5_N72) );
  INV_X1 npu_inst_pe_1_7_5_U107 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_7_5_n6)
         );
  INV_X1 npu_inst_pe_1_7_5_U106 ( .A(npu_inst_pe_1_7_5_n6), .ZN(
        npu_inst_pe_1_7_5_n5) );
  INV_X1 npu_inst_pe_1_7_5_U105 ( .A(npu_inst_n34), .ZN(npu_inst_pe_1_7_5_n2)
         );
  AOI22_X1 npu_inst_pe_1_7_5_U104 ( .A1(npu_inst_pe_1_7_5_n38), .A2(
        int_i_data_v_npu[5]), .B1(npu_inst_pe_1_7_5_n113), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_5_n39) );
  INV_X1 npu_inst_pe_1_7_5_U103 ( .A(npu_inst_pe_1_7_5_n39), .ZN(
        npu_inst_pe_1_7_5_n111) );
  AOI22_X1 npu_inst_pe_1_7_5_U102 ( .A1(npu_inst_pe_1_7_5_n38), .A2(
        int_i_data_v_npu[4]), .B1(npu_inst_pe_1_7_5_n113), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_5_n37) );
  INV_X1 npu_inst_pe_1_7_5_U99 ( .A(npu_inst_pe_1_7_5_n37), .ZN(
        npu_inst_pe_1_7_5_n112) );
  AOI22_X1 npu_inst_pe_1_7_5_U98 ( .A1(int_i_data_v_npu[5]), .A2(
        npu_inst_pe_1_7_5_n58), .B1(npu_inst_pe_1_7_5_n118), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_5_n59) );
  INV_X1 npu_inst_pe_1_7_5_U97 ( .A(npu_inst_pe_1_7_5_n59), .ZN(
        npu_inst_pe_1_7_5_n101) );
  AOI22_X1 npu_inst_pe_1_7_5_U96 ( .A1(int_i_data_v_npu[4]), .A2(
        npu_inst_pe_1_7_5_n58), .B1(npu_inst_pe_1_7_5_n118), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_5_n57) );
  INV_X1 npu_inst_pe_1_7_5_U95 ( .A(npu_inst_pe_1_7_5_n57), .ZN(
        npu_inst_pe_1_7_5_n102) );
  AOI22_X1 npu_inst_pe_1_7_5_U94 ( .A1(int_i_data_v_npu[5]), .A2(
        npu_inst_pe_1_7_5_n54), .B1(npu_inst_pe_1_7_5_n117), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_5_n55) );
  INV_X1 npu_inst_pe_1_7_5_U93 ( .A(npu_inst_pe_1_7_5_n55), .ZN(
        npu_inst_pe_1_7_5_n103) );
  AOI22_X1 npu_inst_pe_1_7_5_U92 ( .A1(int_i_data_v_npu[4]), .A2(
        npu_inst_pe_1_7_5_n54), .B1(npu_inst_pe_1_7_5_n117), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_5_n53) );
  INV_X1 npu_inst_pe_1_7_5_U91 ( .A(npu_inst_pe_1_7_5_n53), .ZN(
        npu_inst_pe_1_7_5_n104) );
  AOI22_X1 npu_inst_pe_1_7_5_U90 ( .A1(int_i_data_v_npu[5]), .A2(
        npu_inst_pe_1_7_5_n50), .B1(npu_inst_pe_1_7_5_n116), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_5_n51) );
  INV_X1 npu_inst_pe_1_7_5_U89 ( .A(npu_inst_pe_1_7_5_n51), .ZN(
        npu_inst_pe_1_7_5_n105) );
  AOI22_X1 npu_inst_pe_1_7_5_U88 ( .A1(int_i_data_v_npu[4]), .A2(
        npu_inst_pe_1_7_5_n50), .B1(npu_inst_pe_1_7_5_n116), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_5_n49) );
  INV_X1 npu_inst_pe_1_7_5_U87 ( .A(npu_inst_pe_1_7_5_n49), .ZN(
        npu_inst_pe_1_7_5_n106) );
  AOI22_X1 npu_inst_pe_1_7_5_U86 ( .A1(int_i_data_v_npu[5]), .A2(
        npu_inst_pe_1_7_5_n46), .B1(npu_inst_pe_1_7_5_n115), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_5_n47) );
  INV_X1 npu_inst_pe_1_7_5_U85 ( .A(npu_inst_pe_1_7_5_n47), .ZN(
        npu_inst_pe_1_7_5_n107) );
  AOI22_X1 npu_inst_pe_1_7_5_U84 ( .A1(int_i_data_v_npu[4]), .A2(
        npu_inst_pe_1_7_5_n46), .B1(npu_inst_pe_1_7_5_n115), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_5_n45) );
  INV_X1 npu_inst_pe_1_7_5_U83 ( .A(npu_inst_pe_1_7_5_n45), .ZN(
        npu_inst_pe_1_7_5_n108) );
  AOI22_X1 npu_inst_pe_1_7_5_U82 ( .A1(int_i_data_v_npu[5]), .A2(
        npu_inst_pe_1_7_5_n42), .B1(npu_inst_pe_1_7_5_n114), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_5_n43) );
  INV_X1 npu_inst_pe_1_7_5_U81 ( .A(npu_inst_pe_1_7_5_n43), .ZN(
        npu_inst_pe_1_7_5_n109) );
  AOI22_X1 npu_inst_pe_1_7_5_U80 ( .A1(int_i_data_v_npu[4]), .A2(
        npu_inst_pe_1_7_5_n42), .B1(npu_inst_pe_1_7_5_n114), .B2(
        npu_inst_pe_1_7_5_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_5_n41) );
  INV_X1 npu_inst_pe_1_7_5_U79 ( .A(npu_inst_pe_1_7_5_n41), .ZN(
        npu_inst_pe_1_7_5_n110) );
  AND2_X1 npu_inst_pe_1_7_5_U78 ( .A1(npu_inst_pe_1_7_5_N93), .A2(npu_inst_n34), .ZN(npu_inst_int_data_y_7__5__0_) );
  NAND2_X1 npu_inst_pe_1_7_5_U77 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_5_n60), .ZN(npu_inst_pe_1_7_5_n74) );
  OAI21_X1 npu_inst_pe_1_7_5_U76 ( .B1(npu_inst_pe_1_7_5_n63), .B2(
        npu_inst_pe_1_7_5_n60), .A(npu_inst_pe_1_7_5_n74), .ZN(
        npu_inst_pe_1_7_5_n97) );
  NAND2_X1 npu_inst_pe_1_7_5_U75 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_5_n60), .ZN(npu_inst_pe_1_7_5_n73) );
  OAI21_X1 npu_inst_pe_1_7_5_U74 ( .B1(npu_inst_pe_1_7_5_n61), .B2(
        npu_inst_pe_1_7_5_n60), .A(npu_inst_pe_1_7_5_n73), .ZN(
        npu_inst_pe_1_7_5_n96) );
  NAND2_X1 npu_inst_pe_1_7_5_U73 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_5_n56), .ZN(npu_inst_pe_1_7_5_n72) );
  OAI21_X1 npu_inst_pe_1_7_5_U72 ( .B1(npu_inst_pe_1_7_5_n63), .B2(
        npu_inst_pe_1_7_5_n56), .A(npu_inst_pe_1_7_5_n72), .ZN(
        npu_inst_pe_1_7_5_n95) );
  NAND2_X1 npu_inst_pe_1_7_5_U71 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_5_n56), .ZN(npu_inst_pe_1_7_5_n71) );
  OAI21_X1 npu_inst_pe_1_7_5_U70 ( .B1(npu_inst_pe_1_7_5_n61), .B2(
        npu_inst_pe_1_7_5_n56), .A(npu_inst_pe_1_7_5_n71), .ZN(
        npu_inst_pe_1_7_5_n94) );
  NAND2_X1 npu_inst_pe_1_7_5_U69 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_5_n52), .ZN(npu_inst_pe_1_7_5_n70) );
  OAI21_X1 npu_inst_pe_1_7_5_U68 ( .B1(npu_inst_pe_1_7_5_n63), .B2(
        npu_inst_pe_1_7_5_n52), .A(npu_inst_pe_1_7_5_n70), .ZN(
        npu_inst_pe_1_7_5_n93) );
  NAND2_X1 npu_inst_pe_1_7_5_U67 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_5_n52), .ZN(npu_inst_pe_1_7_5_n69) );
  OAI21_X1 npu_inst_pe_1_7_5_U66 ( .B1(npu_inst_pe_1_7_5_n61), .B2(
        npu_inst_pe_1_7_5_n52), .A(npu_inst_pe_1_7_5_n69), .ZN(
        npu_inst_pe_1_7_5_n92) );
  NAND2_X1 npu_inst_pe_1_7_5_U65 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_5_n48), .ZN(npu_inst_pe_1_7_5_n68) );
  OAI21_X1 npu_inst_pe_1_7_5_U64 ( .B1(npu_inst_pe_1_7_5_n63), .B2(
        npu_inst_pe_1_7_5_n48), .A(npu_inst_pe_1_7_5_n68), .ZN(
        npu_inst_pe_1_7_5_n91) );
  NAND2_X1 npu_inst_pe_1_7_5_U63 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_5_n48), .ZN(npu_inst_pe_1_7_5_n67) );
  OAI21_X1 npu_inst_pe_1_7_5_U62 ( .B1(npu_inst_pe_1_7_5_n61), .B2(
        npu_inst_pe_1_7_5_n48), .A(npu_inst_pe_1_7_5_n67), .ZN(
        npu_inst_pe_1_7_5_n90) );
  NAND2_X1 npu_inst_pe_1_7_5_U61 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_5_n44), .ZN(npu_inst_pe_1_7_5_n66) );
  OAI21_X1 npu_inst_pe_1_7_5_U60 ( .B1(npu_inst_pe_1_7_5_n63), .B2(
        npu_inst_pe_1_7_5_n44), .A(npu_inst_pe_1_7_5_n66), .ZN(
        npu_inst_pe_1_7_5_n89) );
  NAND2_X1 npu_inst_pe_1_7_5_U59 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_5_n44), .ZN(npu_inst_pe_1_7_5_n65) );
  OAI21_X1 npu_inst_pe_1_7_5_U58 ( .B1(npu_inst_pe_1_7_5_n61), .B2(
        npu_inst_pe_1_7_5_n44), .A(npu_inst_pe_1_7_5_n65), .ZN(
        npu_inst_pe_1_7_5_n88) );
  NAND2_X1 npu_inst_pe_1_7_5_U57 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_5_n40), .ZN(npu_inst_pe_1_7_5_n64) );
  OAI21_X1 npu_inst_pe_1_7_5_U56 ( .B1(npu_inst_pe_1_7_5_n63), .B2(
        npu_inst_pe_1_7_5_n40), .A(npu_inst_pe_1_7_5_n64), .ZN(
        npu_inst_pe_1_7_5_n87) );
  NAND2_X1 npu_inst_pe_1_7_5_U55 ( .A1(npu_inst_pe_1_7_5_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_5_n40), .ZN(npu_inst_pe_1_7_5_n62) );
  OAI21_X1 npu_inst_pe_1_7_5_U54 ( .B1(npu_inst_pe_1_7_5_n61), .B2(
        npu_inst_pe_1_7_5_n40), .A(npu_inst_pe_1_7_5_n62), .ZN(
        npu_inst_pe_1_7_5_n86) );
  AND2_X1 npu_inst_pe_1_7_5_U53 ( .A1(npu_inst_n34), .A2(npu_inst_pe_1_7_5_N94), .ZN(npu_inst_int_data_y_7__5__1_) );
  AOI22_X1 npu_inst_pe_1_7_5_U52 ( .A1(npu_inst_n34), .A2(int_i_data_v_npu[5]), 
        .B1(npu_inst_pe_1_7_5_n2), .B2(npu_inst_int_data_x_7__6__1_), .ZN(
        npu_inst_pe_1_7_5_n63) );
  AOI22_X1 npu_inst_pe_1_7_5_U51 ( .A1(npu_inst_n34), .A2(int_i_data_v_npu[4]), 
        .B1(npu_inst_pe_1_7_5_n2), .B2(npu_inst_int_data_x_7__6__0_), .ZN(
        npu_inst_pe_1_7_5_n61) );
  AOI222_X1 npu_inst_pe_1_7_5_U50 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N73), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N65), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n84) );
  INV_X1 npu_inst_pe_1_7_5_U49 ( .A(npu_inst_pe_1_7_5_n84), .ZN(
        npu_inst_pe_1_7_5_n100) );
  AOI222_X1 npu_inst_pe_1_7_5_U48 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N74), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N66), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n83) );
  INV_X1 npu_inst_pe_1_7_5_U47 ( .A(npu_inst_pe_1_7_5_n83), .ZN(
        npu_inst_pe_1_7_5_n99) );
  AOI222_X1 npu_inst_pe_1_7_5_U46 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N75), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N67), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n82) );
  INV_X1 npu_inst_pe_1_7_5_U45 ( .A(npu_inst_pe_1_7_5_n82), .ZN(
        npu_inst_pe_1_7_5_n98) );
  AOI222_X1 npu_inst_pe_1_7_5_U44 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N76), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N68), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n81) );
  INV_X1 npu_inst_pe_1_7_5_U43 ( .A(npu_inst_pe_1_7_5_n81), .ZN(
        npu_inst_pe_1_7_5_n36) );
  AOI222_X1 npu_inst_pe_1_7_5_U42 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N77), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N69), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n80) );
  INV_X1 npu_inst_pe_1_7_5_U41 ( .A(npu_inst_pe_1_7_5_n80), .ZN(
        npu_inst_pe_1_7_5_n35) );
  AOI222_X1 npu_inst_pe_1_7_5_U40 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N78), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N70), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n79) );
  INV_X1 npu_inst_pe_1_7_5_U39 ( .A(npu_inst_pe_1_7_5_n79), .ZN(
        npu_inst_pe_1_7_5_n34) );
  AOI222_X1 npu_inst_pe_1_7_5_U38 ( .A1(1'b0), .A2(npu_inst_pe_1_7_5_n1), .B1(
        npu_inst_pe_1_7_5_N79), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N71), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n78) );
  INV_X1 npu_inst_pe_1_7_5_U37 ( .A(npu_inst_pe_1_7_5_n78), .ZN(
        npu_inst_pe_1_7_5_n33) );
  AOI222_X1 npu_inst_pe_1_7_5_U36 ( .A1(npu_inst_pe_1_7_5_n1), .A2(1'b0), .B1(
        npu_inst_pe_1_7_5_N80), .B2(npu_inst_pe_1_7_5_n76), .C1(
        npu_inst_pe_1_7_5_N72), .C2(npu_inst_pe_1_7_5_n77), .ZN(
        npu_inst_pe_1_7_5_n75) );
  INV_X1 npu_inst_pe_1_7_5_U35 ( .A(npu_inst_pe_1_7_5_n75), .ZN(
        npu_inst_pe_1_7_5_n32) );
  AND2_X1 npu_inst_pe_1_7_5_U34 ( .A1(npu_inst_int_data_x_7__5__1_), .A2(
        npu_inst_pe_1_7_5_int_q_weight_1_), .ZN(npu_inst_pe_1_7_5_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_5_U33 ( .A1(npu_inst_int_data_x_7__5__0_), .A2(
        npu_inst_pe_1_7_5_int_q_weight_1_), .ZN(npu_inst_pe_1_7_5_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_5_U32 ( .A(npu_inst_pe_1_7_5_int_data_1_), .ZN(
        npu_inst_pe_1_7_5_n13) );
  NOR3_X1 npu_inst_pe_1_7_5_U31 ( .A1(npu_inst_pe_1_7_5_n26), .A2(npu_inst_n34), .A3(npu_inst_int_ckg[2]), .ZN(npu_inst_pe_1_7_5_n85) );
  OR2_X1 npu_inst_pe_1_7_5_U30 ( .A1(npu_inst_pe_1_7_5_n85), .A2(
        npu_inst_pe_1_7_5_n1), .ZN(npu_inst_pe_1_7_5_N84) );
  INV_X1 npu_inst_pe_1_7_5_U29 ( .A(npu_inst_pe_1_7_5_int_data_0_), .ZN(
        npu_inst_pe_1_7_5_n12) );
  INV_X1 npu_inst_pe_1_7_5_U28 ( .A(npu_inst_n49), .ZN(npu_inst_pe_1_7_5_n4)
         );
  OR3_X1 npu_inst_pe_1_7_5_U27 ( .A1(npu_inst_pe_1_7_5_n5), .A2(
        npu_inst_pe_1_7_5_n7), .A3(npu_inst_pe_1_7_5_n4), .ZN(
        npu_inst_pe_1_7_5_n56) );
  OR3_X1 npu_inst_pe_1_7_5_U26 ( .A1(npu_inst_pe_1_7_5_n4), .A2(
        npu_inst_pe_1_7_5_n7), .A3(npu_inst_pe_1_7_5_n6), .ZN(
        npu_inst_pe_1_7_5_n48) );
  INV_X1 npu_inst_pe_1_7_5_U25 ( .A(npu_inst_pe_1_7_5_n4), .ZN(
        npu_inst_pe_1_7_5_n3) );
  OR3_X1 npu_inst_pe_1_7_5_U24 ( .A1(npu_inst_pe_1_7_5_n3), .A2(
        npu_inst_pe_1_7_5_n7), .A3(npu_inst_pe_1_7_5_n6), .ZN(
        npu_inst_pe_1_7_5_n52) );
  OR3_X1 npu_inst_pe_1_7_5_U23 ( .A1(npu_inst_pe_1_7_5_n5), .A2(
        npu_inst_pe_1_7_5_n7), .A3(npu_inst_pe_1_7_5_n3), .ZN(
        npu_inst_pe_1_7_5_n60) );
  BUF_X1 npu_inst_pe_1_7_5_U22 ( .A(npu_inst_n11), .Z(npu_inst_pe_1_7_5_n1) );
  NOR2_X1 npu_inst_pe_1_7_5_U21 ( .A1(npu_inst_pe_1_7_5_n60), .A2(
        npu_inst_pe_1_7_5_n2), .ZN(npu_inst_pe_1_7_5_n58) );
  NOR2_X1 npu_inst_pe_1_7_5_U20 ( .A1(npu_inst_pe_1_7_5_n56), .A2(
        npu_inst_pe_1_7_5_n2), .ZN(npu_inst_pe_1_7_5_n54) );
  NOR2_X1 npu_inst_pe_1_7_5_U19 ( .A1(npu_inst_pe_1_7_5_n52), .A2(
        npu_inst_pe_1_7_5_n2), .ZN(npu_inst_pe_1_7_5_n50) );
  NOR2_X1 npu_inst_pe_1_7_5_U18 ( .A1(npu_inst_pe_1_7_5_n48), .A2(
        npu_inst_pe_1_7_5_n2), .ZN(npu_inst_pe_1_7_5_n46) );
  NOR2_X1 npu_inst_pe_1_7_5_U17 ( .A1(npu_inst_pe_1_7_5_n40), .A2(
        npu_inst_pe_1_7_5_n2), .ZN(npu_inst_pe_1_7_5_n38) );
  NOR2_X1 npu_inst_pe_1_7_5_U16 ( .A1(npu_inst_pe_1_7_5_n44), .A2(
        npu_inst_pe_1_7_5_n2), .ZN(npu_inst_pe_1_7_5_n42) );
  BUF_X1 npu_inst_pe_1_7_5_U15 ( .A(npu_inst_n74), .Z(npu_inst_pe_1_7_5_n7) );
  INV_X1 npu_inst_pe_1_7_5_U14 ( .A(npu_inst_n104), .ZN(npu_inst_pe_1_7_5_n11)
         );
  INV_X1 npu_inst_pe_1_7_5_U13 ( .A(npu_inst_pe_1_7_5_n38), .ZN(
        npu_inst_pe_1_7_5_n113) );
  INV_X1 npu_inst_pe_1_7_5_U12 ( .A(npu_inst_pe_1_7_5_n58), .ZN(
        npu_inst_pe_1_7_5_n118) );
  INV_X1 npu_inst_pe_1_7_5_U11 ( .A(npu_inst_pe_1_7_5_n54), .ZN(
        npu_inst_pe_1_7_5_n117) );
  INV_X1 npu_inst_pe_1_7_5_U10 ( .A(npu_inst_pe_1_7_5_n50), .ZN(
        npu_inst_pe_1_7_5_n116) );
  INV_X1 npu_inst_pe_1_7_5_U9 ( .A(npu_inst_pe_1_7_5_n46), .ZN(
        npu_inst_pe_1_7_5_n115) );
  INV_X1 npu_inst_pe_1_7_5_U8 ( .A(npu_inst_pe_1_7_5_n42), .ZN(
        npu_inst_pe_1_7_5_n114) );
  BUF_X1 npu_inst_pe_1_7_5_U7 ( .A(npu_inst_pe_1_7_5_n11), .Z(
        npu_inst_pe_1_7_5_n10) );
  BUF_X1 npu_inst_pe_1_7_5_U6 ( .A(npu_inst_pe_1_7_5_n11), .Z(
        npu_inst_pe_1_7_5_n9) );
  BUF_X1 npu_inst_pe_1_7_5_U5 ( .A(npu_inst_pe_1_7_5_n11), .Z(
        npu_inst_pe_1_7_5_n8) );
  NOR2_X1 npu_inst_pe_1_7_5_U4 ( .A1(npu_inst_pe_1_7_5_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_5_n1), .ZN(npu_inst_pe_1_7_5_n76) );
  NOR2_X1 npu_inst_pe_1_7_5_U3 ( .A1(npu_inst_pe_1_7_5_n27), .A2(
        npu_inst_pe_1_7_5_n1), .ZN(npu_inst_pe_1_7_5_n77) );
  FA_X1 npu_inst_pe_1_7_5_sub_77_U2_1 ( .A(npu_inst_int_data_res_7__5__1_), 
        .B(npu_inst_pe_1_7_5_n13), .CI(npu_inst_pe_1_7_5_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_7_5_sub_77_carry_2_), .S(npu_inst_pe_1_7_5_N66) );
  FA_X1 npu_inst_pe_1_7_5_add_79_U1_1 ( .A(npu_inst_int_data_res_7__5__1_), 
        .B(npu_inst_pe_1_7_5_int_data_1_), .CI(
        npu_inst_pe_1_7_5_add_79_carry_1_), .CO(
        npu_inst_pe_1_7_5_add_79_carry_2_), .S(npu_inst_pe_1_7_5_N74) );
  NAND3_X1 npu_inst_pe_1_7_5_U101 ( .A1(npu_inst_pe_1_7_5_n4), .A2(
        npu_inst_pe_1_7_5_n6), .A3(npu_inst_pe_1_7_5_n7), .ZN(
        npu_inst_pe_1_7_5_n44) );
  NAND3_X1 npu_inst_pe_1_7_5_U100 ( .A1(npu_inst_pe_1_7_5_n3), .A2(
        npu_inst_pe_1_7_5_n6), .A3(npu_inst_pe_1_7_5_n7), .ZN(
        npu_inst_pe_1_7_5_n40) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_5_n33), .CK(
        npu_inst_pe_1_7_5_net3075), .RN(npu_inst_pe_1_7_5_n8), .Q(
        npu_inst_int_data_res_7__5__6_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_5_n34), .CK(
        npu_inst_pe_1_7_5_net3075), .RN(npu_inst_pe_1_7_5_n8), .Q(
        npu_inst_int_data_res_7__5__5_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_5_n35), .CK(
        npu_inst_pe_1_7_5_net3075), .RN(npu_inst_pe_1_7_5_n8), .Q(
        npu_inst_int_data_res_7__5__4_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_5_n36), .CK(
        npu_inst_pe_1_7_5_net3075), .RN(npu_inst_pe_1_7_5_n8), .Q(
        npu_inst_int_data_res_7__5__3_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_5_n98), .CK(
        npu_inst_pe_1_7_5_net3075), .RN(npu_inst_pe_1_7_5_n8), .Q(
        npu_inst_int_data_res_7__5__2_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_5_n99), .CK(
        npu_inst_pe_1_7_5_net3075), .RN(npu_inst_pe_1_7_5_n8), .Q(
        npu_inst_int_data_res_7__5__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_5_n32), .CK(
        npu_inst_pe_1_7_5_net3075), .RN(npu_inst_pe_1_7_5_n8), .Q(
        npu_inst_int_data_res_7__5__7_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_5_n100), 
        .CK(npu_inst_pe_1_7_5_net3075), .RN(npu_inst_pe_1_7_5_n8), .Q(
        npu_inst_int_data_res_7__5__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_weight_reg_0_ ( .D(npu_inst_n90), .CK(
        npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n8), .Q(
        npu_inst_pe_1_7_5_int_q_weight_0_), .QN(npu_inst_pe_1_7_5_n27) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_weight_reg_1_ ( .D(npu_inst_n96), .CK(
        npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n8), .Q(
        npu_inst_pe_1_7_5_int_q_weight_1_), .QN(npu_inst_pe_1_7_5_n26) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_5_n112), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n8), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_5_n111), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n8), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_5_n110), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_5_n109), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_5_n108), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_5_n107), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_5_n106), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_5_n105), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_5_n104), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_5_n103), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_5_n102), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_5_n101), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_5_n86), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_5_n87), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n9), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_5_n88), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_5_n89), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_5_n90), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_5_n91), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_5_n92), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_5_n93), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_5_n94), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_5_n95), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_5_n96), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_5_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_5_n97), 
        .CK(npu_inst_pe_1_7_5_net3081), .RN(npu_inst_pe_1_7_5_n10), .Q(
        npu_inst_pe_1_7_5_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_5_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_5_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_5_net3075) );
  CLKGATETST_X1 npu_inst_pe_1_7_5_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n43), .SE(1'b0), .GCK(npu_inst_pe_1_7_5_net3081) );
  MUX2_X1 npu_inst_pe_1_7_6_U153 ( .A(npu_inst_pe_1_7_6_n31), .B(
        npu_inst_pe_1_7_6_n28), .S(npu_inst_pe_1_7_6_n7), .Z(
        npu_inst_pe_1_7_6_N93) );
  MUX2_X1 npu_inst_pe_1_7_6_U152 ( .A(npu_inst_pe_1_7_6_n30), .B(
        npu_inst_pe_1_7_6_n29), .S(npu_inst_pe_1_7_6_n5), .Z(
        npu_inst_pe_1_7_6_n31) );
  MUX2_X1 npu_inst_pe_1_7_6_U151 ( .A(npu_inst_pe_1_7_6_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_6_n3), .Z(
        npu_inst_pe_1_7_6_n30) );
  MUX2_X1 npu_inst_pe_1_7_6_U150 ( .A(npu_inst_pe_1_7_6_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_6_n3), .Z(
        npu_inst_pe_1_7_6_n29) );
  MUX2_X1 npu_inst_pe_1_7_6_U149 ( .A(npu_inst_pe_1_7_6_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_6_n3), .Z(
        npu_inst_pe_1_7_6_n28) );
  MUX2_X1 npu_inst_pe_1_7_6_U148 ( .A(npu_inst_pe_1_7_6_n25), .B(
        npu_inst_pe_1_7_6_n22), .S(npu_inst_pe_1_7_6_n7), .Z(
        npu_inst_pe_1_7_6_N94) );
  MUX2_X1 npu_inst_pe_1_7_6_U147 ( .A(npu_inst_pe_1_7_6_n24), .B(
        npu_inst_pe_1_7_6_n23), .S(npu_inst_pe_1_7_6_n5), .Z(
        npu_inst_pe_1_7_6_n25) );
  MUX2_X1 npu_inst_pe_1_7_6_U146 ( .A(npu_inst_pe_1_7_6_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_6_n3), .Z(
        npu_inst_pe_1_7_6_n24) );
  MUX2_X1 npu_inst_pe_1_7_6_U145 ( .A(npu_inst_pe_1_7_6_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_6_n3), .Z(
        npu_inst_pe_1_7_6_n23) );
  MUX2_X1 npu_inst_pe_1_7_6_U144 ( .A(npu_inst_pe_1_7_6_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_6_n3), .Z(
        npu_inst_pe_1_7_6_n22) );
  MUX2_X1 npu_inst_pe_1_7_6_U143 ( .A(npu_inst_pe_1_7_6_n21), .B(
        npu_inst_pe_1_7_6_n18), .S(npu_inst_pe_1_7_6_n7), .Z(
        npu_inst_int_data_x_7__6__1_) );
  MUX2_X1 npu_inst_pe_1_7_6_U142 ( .A(npu_inst_pe_1_7_6_n20), .B(
        npu_inst_pe_1_7_6_n19), .S(npu_inst_pe_1_7_6_n5), .Z(
        npu_inst_pe_1_7_6_n21) );
  MUX2_X1 npu_inst_pe_1_7_6_U141 ( .A(npu_inst_pe_1_7_6_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_6_n3), .Z(
        npu_inst_pe_1_7_6_n20) );
  MUX2_X1 npu_inst_pe_1_7_6_U140 ( .A(npu_inst_pe_1_7_6_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_6_n3), .Z(
        npu_inst_pe_1_7_6_n19) );
  MUX2_X1 npu_inst_pe_1_7_6_U139 ( .A(npu_inst_pe_1_7_6_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_6_n3), .Z(
        npu_inst_pe_1_7_6_n18) );
  MUX2_X1 npu_inst_pe_1_7_6_U138 ( .A(npu_inst_pe_1_7_6_n17), .B(
        npu_inst_pe_1_7_6_n14), .S(npu_inst_pe_1_7_6_n7), .Z(
        npu_inst_int_data_x_7__6__0_) );
  MUX2_X1 npu_inst_pe_1_7_6_U137 ( .A(npu_inst_pe_1_7_6_n16), .B(
        npu_inst_pe_1_7_6_n15), .S(npu_inst_pe_1_7_6_n5), .Z(
        npu_inst_pe_1_7_6_n17) );
  MUX2_X1 npu_inst_pe_1_7_6_U136 ( .A(npu_inst_pe_1_7_6_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_6_n3), .Z(
        npu_inst_pe_1_7_6_n16) );
  MUX2_X1 npu_inst_pe_1_7_6_U135 ( .A(npu_inst_pe_1_7_6_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_6_n3), .Z(
        npu_inst_pe_1_7_6_n15) );
  MUX2_X1 npu_inst_pe_1_7_6_U134 ( .A(npu_inst_pe_1_7_6_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_6_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_6_n3), .Z(
        npu_inst_pe_1_7_6_n14) );
  XOR2_X1 npu_inst_pe_1_7_6_U133 ( .A(npu_inst_pe_1_7_6_int_data_0_), .B(
        npu_inst_int_data_res_7__6__0_), .Z(npu_inst_pe_1_7_6_N73) );
  AND2_X1 npu_inst_pe_1_7_6_U132 ( .A1(npu_inst_int_data_res_7__6__0_), .A2(
        npu_inst_pe_1_7_6_int_data_0_), .ZN(npu_inst_pe_1_7_6_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_6_U131 ( .A(npu_inst_int_data_res_7__6__0_), .B(
        npu_inst_pe_1_7_6_n12), .ZN(npu_inst_pe_1_7_6_N65) );
  OR2_X1 npu_inst_pe_1_7_6_U130 ( .A1(npu_inst_pe_1_7_6_n12), .A2(
        npu_inst_int_data_res_7__6__0_), .ZN(npu_inst_pe_1_7_6_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_6_U129 ( .A(npu_inst_int_data_res_7__6__2_), .B(
        npu_inst_pe_1_7_6_add_79_carry_2_), .Z(npu_inst_pe_1_7_6_N75) );
  AND2_X1 npu_inst_pe_1_7_6_U128 ( .A1(npu_inst_pe_1_7_6_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_7__6__2_), .ZN(
        npu_inst_pe_1_7_6_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_6_U127 ( .A(npu_inst_int_data_res_7__6__3_), .B(
        npu_inst_pe_1_7_6_add_79_carry_3_), .Z(npu_inst_pe_1_7_6_N76) );
  AND2_X1 npu_inst_pe_1_7_6_U126 ( .A1(npu_inst_pe_1_7_6_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_7__6__3_), .ZN(
        npu_inst_pe_1_7_6_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_6_U125 ( .A(npu_inst_int_data_res_7__6__4_), .B(
        npu_inst_pe_1_7_6_add_79_carry_4_), .Z(npu_inst_pe_1_7_6_N77) );
  AND2_X1 npu_inst_pe_1_7_6_U124 ( .A1(npu_inst_pe_1_7_6_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_7__6__4_), .ZN(
        npu_inst_pe_1_7_6_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_6_U123 ( .A(npu_inst_int_data_res_7__6__5_), .B(
        npu_inst_pe_1_7_6_add_79_carry_5_), .Z(npu_inst_pe_1_7_6_N78) );
  AND2_X1 npu_inst_pe_1_7_6_U122 ( .A1(npu_inst_pe_1_7_6_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_7__6__5_), .ZN(
        npu_inst_pe_1_7_6_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_6_U121 ( .A(npu_inst_int_data_res_7__6__6_), .B(
        npu_inst_pe_1_7_6_add_79_carry_6_), .Z(npu_inst_pe_1_7_6_N79) );
  AND2_X1 npu_inst_pe_1_7_6_U120 ( .A1(npu_inst_pe_1_7_6_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_7__6__6_), .ZN(
        npu_inst_pe_1_7_6_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_6_U119 ( .A(npu_inst_int_data_res_7__6__7_), .B(
        npu_inst_pe_1_7_6_add_79_carry_7_), .Z(npu_inst_pe_1_7_6_N80) );
  XNOR2_X1 npu_inst_pe_1_7_6_U118 ( .A(npu_inst_pe_1_7_6_sub_77_carry_2_), .B(
        npu_inst_int_data_res_7__6__2_), .ZN(npu_inst_pe_1_7_6_N67) );
  OR2_X1 npu_inst_pe_1_7_6_U117 ( .A1(npu_inst_int_data_res_7__6__2_), .A2(
        npu_inst_pe_1_7_6_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_7_6_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_6_U116 ( .A(npu_inst_pe_1_7_6_sub_77_carry_3_), .B(
        npu_inst_int_data_res_7__6__3_), .ZN(npu_inst_pe_1_7_6_N68) );
  OR2_X1 npu_inst_pe_1_7_6_U115 ( .A1(npu_inst_int_data_res_7__6__3_), .A2(
        npu_inst_pe_1_7_6_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_7_6_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_6_U114 ( .A(npu_inst_pe_1_7_6_sub_77_carry_4_), .B(
        npu_inst_int_data_res_7__6__4_), .ZN(npu_inst_pe_1_7_6_N69) );
  OR2_X1 npu_inst_pe_1_7_6_U113 ( .A1(npu_inst_int_data_res_7__6__4_), .A2(
        npu_inst_pe_1_7_6_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_7_6_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_6_U112 ( .A(npu_inst_pe_1_7_6_sub_77_carry_5_), .B(
        npu_inst_int_data_res_7__6__5_), .ZN(npu_inst_pe_1_7_6_N70) );
  OR2_X1 npu_inst_pe_1_7_6_U111 ( .A1(npu_inst_int_data_res_7__6__5_), .A2(
        npu_inst_pe_1_7_6_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_7_6_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_6_U110 ( .A(npu_inst_pe_1_7_6_sub_77_carry_6_), .B(
        npu_inst_int_data_res_7__6__6_), .ZN(npu_inst_pe_1_7_6_N71) );
  OR2_X1 npu_inst_pe_1_7_6_U109 ( .A1(npu_inst_int_data_res_7__6__6_), .A2(
        npu_inst_pe_1_7_6_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_7_6_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_6_U108 ( .A(npu_inst_int_data_res_7__6__7_), .B(
        npu_inst_pe_1_7_6_sub_77_carry_7_), .ZN(npu_inst_pe_1_7_6_N72) );
  INV_X1 npu_inst_pe_1_7_6_U107 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_7_6_n6)
         );
  INV_X1 npu_inst_pe_1_7_6_U106 ( .A(npu_inst_pe_1_7_6_n6), .ZN(
        npu_inst_pe_1_7_6_n5) );
  INV_X1 npu_inst_pe_1_7_6_U105 ( .A(npu_inst_n34), .ZN(npu_inst_pe_1_7_6_n2)
         );
  AOI22_X1 npu_inst_pe_1_7_6_U104 ( .A1(npu_inst_pe_1_7_6_n38), .A2(
        int_i_data_v_npu[3]), .B1(npu_inst_pe_1_7_6_n113), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_6_n39) );
  INV_X1 npu_inst_pe_1_7_6_U103 ( .A(npu_inst_pe_1_7_6_n39), .ZN(
        npu_inst_pe_1_7_6_n111) );
  AOI22_X1 npu_inst_pe_1_7_6_U102 ( .A1(npu_inst_pe_1_7_6_n38), .A2(
        int_i_data_v_npu[2]), .B1(npu_inst_pe_1_7_6_n113), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_6_n37) );
  INV_X1 npu_inst_pe_1_7_6_U99 ( .A(npu_inst_pe_1_7_6_n37), .ZN(
        npu_inst_pe_1_7_6_n112) );
  AOI22_X1 npu_inst_pe_1_7_6_U98 ( .A1(int_i_data_v_npu[3]), .A2(
        npu_inst_pe_1_7_6_n58), .B1(npu_inst_pe_1_7_6_n118), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_6_n59) );
  INV_X1 npu_inst_pe_1_7_6_U97 ( .A(npu_inst_pe_1_7_6_n59), .ZN(
        npu_inst_pe_1_7_6_n101) );
  AOI22_X1 npu_inst_pe_1_7_6_U96 ( .A1(int_i_data_v_npu[2]), .A2(
        npu_inst_pe_1_7_6_n58), .B1(npu_inst_pe_1_7_6_n118), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_6_n57) );
  INV_X1 npu_inst_pe_1_7_6_U95 ( .A(npu_inst_pe_1_7_6_n57), .ZN(
        npu_inst_pe_1_7_6_n102) );
  AOI22_X1 npu_inst_pe_1_7_6_U94 ( .A1(int_i_data_v_npu[3]), .A2(
        npu_inst_pe_1_7_6_n54), .B1(npu_inst_pe_1_7_6_n117), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_6_n55) );
  INV_X1 npu_inst_pe_1_7_6_U93 ( .A(npu_inst_pe_1_7_6_n55), .ZN(
        npu_inst_pe_1_7_6_n103) );
  AOI22_X1 npu_inst_pe_1_7_6_U92 ( .A1(int_i_data_v_npu[2]), .A2(
        npu_inst_pe_1_7_6_n54), .B1(npu_inst_pe_1_7_6_n117), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_6_n53) );
  INV_X1 npu_inst_pe_1_7_6_U91 ( .A(npu_inst_pe_1_7_6_n53), .ZN(
        npu_inst_pe_1_7_6_n104) );
  AOI22_X1 npu_inst_pe_1_7_6_U90 ( .A1(int_i_data_v_npu[3]), .A2(
        npu_inst_pe_1_7_6_n50), .B1(npu_inst_pe_1_7_6_n116), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_6_n51) );
  INV_X1 npu_inst_pe_1_7_6_U89 ( .A(npu_inst_pe_1_7_6_n51), .ZN(
        npu_inst_pe_1_7_6_n105) );
  AOI22_X1 npu_inst_pe_1_7_6_U88 ( .A1(int_i_data_v_npu[2]), .A2(
        npu_inst_pe_1_7_6_n50), .B1(npu_inst_pe_1_7_6_n116), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_6_n49) );
  INV_X1 npu_inst_pe_1_7_6_U87 ( .A(npu_inst_pe_1_7_6_n49), .ZN(
        npu_inst_pe_1_7_6_n106) );
  AOI22_X1 npu_inst_pe_1_7_6_U86 ( .A1(int_i_data_v_npu[3]), .A2(
        npu_inst_pe_1_7_6_n46), .B1(npu_inst_pe_1_7_6_n115), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_6_n47) );
  INV_X1 npu_inst_pe_1_7_6_U85 ( .A(npu_inst_pe_1_7_6_n47), .ZN(
        npu_inst_pe_1_7_6_n107) );
  AOI22_X1 npu_inst_pe_1_7_6_U84 ( .A1(int_i_data_v_npu[2]), .A2(
        npu_inst_pe_1_7_6_n46), .B1(npu_inst_pe_1_7_6_n115), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_6_n45) );
  INV_X1 npu_inst_pe_1_7_6_U83 ( .A(npu_inst_pe_1_7_6_n45), .ZN(
        npu_inst_pe_1_7_6_n108) );
  AOI22_X1 npu_inst_pe_1_7_6_U82 ( .A1(int_i_data_v_npu[3]), .A2(
        npu_inst_pe_1_7_6_n42), .B1(npu_inst_pe_1_7_6_n114), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_6_n43) );
  INV_X1 npu_inst_pe_1_7_6_U81 ( .A(npu_inst_pe_1_7_6_n43), .ZN(
        npu_inst_pe_1_7_6_n109) );
  AOI22_X1 npu_inst_pe_1_7_6_U80 ( .A1(int_i_data_v_npu[2]), .A2(
        npu_inst_pe_1_7_6_n42), .B1(npu_inst_pe_1_7_6_n114), .B2(
        npu_inst_pe_1_7_6_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_6_n41) );
  INV_X1 npu_inst_pe_1_7_6_U79 ( .A(npu_inst_pe_1_7_6_n41), .ZN(
        npu_inst_pe_1_7_6_n110) );
  AND2_X1 npu_inst_pe_1_7_6_U78 ( .A1(npu_inst_pe_1_7_6_N93), .A2(npu_inst_n34), .ZN(npu_inst_int_data_y_7__6__0_) );
  NAND2_X1 npu_inst_pe_1_7_6_U77 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_6_n60), .ZN(npu_inst_pe_1_7_6_n74) );
  OAI21_X1 npu_inst_pe_1_7_6_U76 ( .B1(npu_inst_pe_1_7_6_n63), .B2(
        npu_inst_pe_1_7_6_n60), .A(npu_inst_pe_1_7_6_n74), .ZN(
        npu_inst_pe_1_7_6_n97) );
  NAND2_X1 npu_inst_pe_1_7_6_U75 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_6_n60), .ZN(npu_inst_pe_1_7_6_n73) );
  OAI21_X1 npu_inst_pe_1_7_6_U74 ( .B1(npu_inst_pe_1_7_6_n61), .B2(
        npu_inst_pe_1_7_6_n60), .A(npu_inst_pe_1_7_6_n73), .ZN(
        npu_inst_pe_1_7_6_n96) );
  NAND2_X1 npu_inst_pe_1_7_6_U73 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_6_n56), .ZN(npu_inst_pe_1_7_6_n72) );
  OAI21_X1 npu_inst_pe_1_7_6_U72 ( .B1(npu_inst_pe_1_7_6_n63), .B2(
        npu_inst_pe_1_7_6_n56), .A(npu_inst_pe_1_7_6_n72), .ZN(
        npu_inst_pe_1_7_6_n95) );
  NAND2_X1 npu_inst_pe_1_7_6_U71 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_6_n56), .ZN(npu_inst_pe_1_7_6_n71) );
  OAI21_X1 npu_inst_pe_1_7_6_U70 ( .B1(npu_inst_pe_1_7_6_n61), .B2(
        npu_inst_pe_1_7_6_n56), .A(npu_inst_pe_1_7_6_n71), .ZN(
        npu_inst_pe_1_7_6_n94) );
  NAND2_X1 npu_inst_pe_1_7_6_U69 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_6_n52), .ZN(npu_inst_pe_1_7_6_n70) );
  OAI21_X1 npu_inst_pe_1_7_6_U68 ( .B1(npu_inst_pe_1_7_6_n63), .B2(
        npu_inst_pe_1_7_6_n52), .A(npu_inst_pe_1_7_6_n70), .ZN(
        npu_inst_pe_1_7_6_n93) );
  NAND2_X1 npu_inst_pe_1_7_6_U67 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_6_n52), .ZN(npu_inst_pe_1_7_6_n69) );
  OAI21_X1 npu_inst_pe_1_7_6_U66 ( .B1(npu_inst_pe_1_7_6_n61), .B2(
        npu_inst_pe_1_7_6_n52), .A(npu_inst_pe_1_7_6_n69), .ZN(
        npu_inst_pe_1_7_6_n92) );
  NAND2_X1 npu_inst_pe_1_7_6_U65 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_6_n48), .ZN(npu_inst_pe_1_7_6_n68) );
  OAI21_X1 npu_inst_pe_1_7_6_U64 ( .B1(npu_inst_pe_1_7_6_n63), .B2(
        npu_inst_pe_1_7_6_n48), .A(npu_inst_pe_1_7_6_n68), .ZN(
        npu_inst_pe_1_7_6_n91) );
  NAND2_X1 npu_inst_pe_1_7_6_U63 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_6_n48), .ZN(npu_inst_pe_1_7_6_n67) );
  OAI21_X1 npu_inst_pe_1_7_6_U62 ( .B1(npu_inst_pe_1_7_6_n61), .B2(
        npu_inst_pe_1_7_6_n48), .A(npu_inst_pe_1_7_6_n67), .ZN(
        npu_inst_pe_1_7_6_n90) );
  NAND2_X1 npu_inst_pe_1_7_6_U61 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_6_n44), .ZN(npu_inst_pe_1_7_6_n66) );
  OAI21_X1 npu_inst_pe_1_7_6_U60 ( .B1(npu_inst_pe_1_7_6_n63), .B2(
        npu_inst_pe_1_7_6_n44), .A(npu_inst_pe_1_7_6_n66), .ZN(
        npu_inst_pe_1_7_6_n89) );
  NAND2_X1 npu_inst_pe_1_7_6_U59 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_6_n44), .ZN(npu_inst_pe_1_7_6_n65) );
  OAI21_X1 npu_inst_pe_1_7_6_U58 ( .B1(npu_inst_pe_1_7_6_n61), .B2(
        npu_inst_pe_1_7_6_n44), .A(npu_inst_pe_1_7_6_n65), .ZN(
        npu_inst_pe_1_7_6_n88) );
  NAND2_X1 npu_inst_pe_1_7_6_U57 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_6_n40), .ZN(npu_inst_pe_1_7_6_n64) );
  OAI21_X1 npu_inst_pe_1_7_6_U56 ( .B1(npu_inst_pe_1_7_6_n63), .B2(
        npu_inst_pe_1_7_6_n40), .A(npu_inst_pe_1_7_6_n64), .ZN(
        npu_inst_pe_1_7_6_n87) );
  NAND2_X1 npu_inst_pe_1_7_6_U55 ( .A1(npu_inst_pe_1_7_6_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_6_n40), .ZN(npu_inst_pe_1_7_6_n62) );
  OAI21_X1 npu_inst_pe_1_7_6_U54 ( .B1(npu_inst_pe_1_7_6_n61), .B2(
        npu_inst_pe_1_7_6_n40), .A(npu_inst_pe_1_7_6_n62), .ZN(
        npu_inst_pe_1_7_6_n86) );
  AND2_X1 npu_inst_pe_1_7_6_U53 ( .A1(npu_inst_n34), .A2(npu_inst_pe_1_7_6_N94), .ZN(npu_inst_int_data_y_7__6__1_) );
  AOI22_X1 npu_inst_pe_1_7_6_U52 ( .A1(npu_inst_n34), .A2(int_i_data_v_npu[3]), 
        .B1(npu_inst_pe_1_7_6_n2), .B2(npu_inst_int_data_x_7__7__1_), .ZN(
        npu_inst_pe_1_7_6_n63) );
  AOI22_X1 npu_inst_pe_1_7_6_U51 ( .A1(npu_inst_n34), .A2(int_i_data_v_npu[2]), 
        .B1(npu_inst_pe_1_7_6_n2), .B2(npu_inst_int_data_x_7__7__0_), .ZN(
        npu_inst_pe_1_7_6_n61) );
  AOI222_X1 npu_inst_pe_1_7_6_U50 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N73), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N65), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n84) );
  INV_X1 npu_inst_pe_1_7_6_U49 ( .A(npu_inst_pe_1_7_6_n84), .ZN(
        npu_inst_pe_1_7_6_n100) );
  AOI222_X1 npu_inst_pe_1_7_6_U48 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N74), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N66), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n83) );
  INV_X1 npu_inst_pe_1_7_6_U47 ( .A(npu_inst_pe_1_7_6_n83), .ZN(
        npu_inst_pe_1_7_6_n99) );
  AOI222_X1 npu_inst_pe_1_7_6_U46 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N75), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N67), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n82) );
  INV_X1 npu_inst_pe_1_7_6_U45 ( .A(npu_inst_pe_1_7_6_n82), .ZN(
        npu_inst_pe_1_7_6_n98) );
  AOI222_X1 npu_inst_pe_1_7_6_U44 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N76), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N68), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n81) );
  INV_X1 npu_inst_pe_1_7_6_U43 ( .A(npu_inst_pe_1_7_6_n81), .ZN(
        npu_inst_pe_1_7_6_n36) );
  AOI222_X1 npu_inst_pe_1_7_6_U42 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N77), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N69), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n80) );
  INV_X1 npu_inst_pe_1_7_6_U41 ( .A(npu_inst_pe_1_7_6_n80), .ZN(
        npu_inst_pe_1_7_6_n35) );
  AOI222_X1 npu_inst_pe_1_7_6_U40 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N78), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N70), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n79) );
  INV_X1 npu_inst_pe_1_7_6_U39 ( .A(npu_inst_pe_1_7_6_n79), .ZN(
        npu_inst_pe_1_7_6_n34) );
  AOI222_X1 npu_inst_pe_1_7_6_U38 ( .A1(1'b0), .A2(npu_inst_pe_1_7_6_n1), .B1(
        npu_inst_pe_1_7_6_N79), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N71), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n78) );
  INV_X1 npu_inst_pe_1_7_6_U37 ( .A(npu_inst_pe_1_7_6_n78), .ZN(
        npu_inst_pe_1_7_6_n33) );
  AOI222_X1 npu_inst_pe_1_7_6_U36 ( .A1(npu_inst_pe_1_7_6_n1), .A2(1'b0), .B1(
        npu_inst_pe_1_7_6_N80), .B2(npu_inst_pe_1_7_6_n76), .C1(
        npu_inst_pe_1_7_6_N72), .C2(npu_inst_pe_1_7_6_n77), .ZN(
        npu_inst_pe_1_7_6_n75) );
  INV_X1 npu_inst_pe_1_7_6_U35 ( .A(npu_inst_pe_1_7_6_n75), .ZN(
        npu_inst_pe_1_7_6_n32) );
  AND2_X1 npu_inst_pe_1_7_6_U34 ( .A1(npu_inst_int_data_x_7__6__1_), .A2(
        npu_inst_pe_1_7_6_int_q_weight_1_), .ZN(npu_inst_pe_1_7_6_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_6_U33 ( .A1(npu_inst_int_data_x_7__6__0_), .A2(
        npu_inst_pe_1_7_6_int_q_weight_1_), .ZN(npu_inst_pe_1_7_6_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_6_U32 ( .A(npu_inst_pe_1_7_6_int_data_1_), .ZN(
        npu_inst_pe_1_7_6_n13) );
  NOR3_X1 npu_inst_pe_1_7_6_U31 ( .A1(npu_inst_pe_1_7_6_n26), .A2(npu_inst_n34), .A3(npu_inst_int_ckg[1]), .ZN(npu_inst_pe_1_7_6_n85) );
  OR2_X1 npu_inst_pe_1_7_6_U30 ( .A1(npu_inst_pe_1_7_6_n85), .A2(
        npu_inst_pe_1_7_6_n1), .ZN(npu_inst_pe_1_7_6_N84) );
  INV_X1 npu_inst_pe_1_7_6_U29 ( .A(npu_inst_pe_1_7_6_int_data_0_), .ZN(
        npu_inst_pe_1_7_6_n12) );
  INV_X1 npu_inst_pe_1_7_6_U28 ( .A(npu_inst_n49), .ZN(npu_inst_pe_1_7_6_n4)
         );
  OR3_X1 npu_inst_pe_1_7_6_U27 ( .A1(npu_inst_pe_1_7_6_n5), .A2(
        npu_inst_pe_1_7_6_n7), .A3(npu_inst_pe_1_7_6_n4), .ZN(
        npu_inst_pe_1_7_6_n56) );
  OR3_X1 npu_inst_pe_1_7_6_U26 ( .A1(npu_inst_pe_1_7_6_n4), .A2(
        npu_inst_pe_1_7_6_n7), .A3(npu_inst_pe_1_7_6_n6), .ZN(
        npu_inst_pe_1_7_6_n48) );
  INV_X1 npu_inst_pe_1_7_6_U25 ( .A(npu_inst_pe_1_7_6_n4), .ZN(
        npu_inst_pe_1_7_6_n3) );
  OR3_X1 npu_inst_pe_1_7_6_U24 ( .A1(npu_inst_pe_1_7_6_n3), .A2(
        npu_inst_pe_1_7_6_n7), .A3(npu_inst_pe_1_7_6_n6), .ZN(
        npu_inst_pe_1_7_6_n52) );
  OR3_X1 npu_inst_pe_1_7_6_U23 ( .A1(npu_inst_pe_1_7_6_n5), .A2(
        npu_inst_pe_1_7_6_n7), .A3(npu_inst_pe_1_7_6_n3), .ZN(
        npu_inst_pe_1_7_6_n60) );
  BUF_X1 npu_inst_pe_1_7_6_U22 ( .A(npu_inst_n11), .Z(npu_inst_pe_1_7_6_n1) );
  NOR2_X1 npu_inst_pe_1_7_6_U21 ( .A1(npu_inst_pe_1_7_6_n60), .A2(
        npu_inst_pe_1_7_6_n2), .ZN(npu_inst_pe_1_7_6_n58) );
  NOR2_X1 npu_inst_pe_1_7_6_U20 ( .A1(npu_inst_pe_1_7_6_n56), .A2(
        npu_inst_pe_1_7_6_n2), .ZN(npu_inst_pe_1_7_6_n54) );
  NOR2_X1 npu_inst_pe_1_7_6_U19 ( .A1(npu_inst_pe_1_7_6_n52), .A2(
        npu_inst_pe_1_7_6_n2), .ZN(npu_inst_pe_1_7_6_n50) );
  NOR2_X1 npu_inst_pe_1_7_6_U18 ( .A1(npu_inst_pe_1_7_6_n48), .A2(
        npu_inst_pe_1_7_6_n2), .ZN(npu_inst_pe_1_7_6_n46) );
  NOR2_X1 npu_inst_pe_1_7_6_U17 ( .A1(npu_inst_pe_1_7_6_n40), .A2(
        npu_inst_pe_1_7_6_n2), .ZN(npu_inst_pe_1_7_6_n38) );
  NOR2_X1 npu_inst_pe_1_7_6_U16 ( .A1(npu_inst_pe_1_7_6_n44), .A2(
        npu_inst_pe_1_7_6_n2), .ZN(npu_inst_pe_1_7_6_n42) );
  BUF_X1 npu_inst_pe_1_7_6_U15 ( .A(npu_inst_n74), .Z(npu_inst_pe_1_7_6_n7) );
  INV_X1 npu_inst_pe_1_7_6_U14 ( .A(npu_inst_n104), .ZN(npu_inst_pe_1_7_6_n11)
         );
  INV_X1 npu_inst_pe_1_7_6_U13 ( .A(npu_inst_pe_1_7_6_n38), .ZN(
        npu_inst_pe_1_7_6_n113) );
  INV_X1 npu_inst_pe_1_7_6_U12 ( .A(npu_inst_pe_1_7_6_n58), .ZN(
        npu_inst_pe_1_7_6_n118) );
  INV_X1 npu_inst_pe_1_7_6_U11 ( .A(npu_inst_pe_1_7_6_n54), .ZN(
        npu_inst_pe_1_7_6_n117) );
  INV_X1 npu_inst_pe_1_7_6_U10 ( .A(npu_inst_pe_1_7_6_n50), .ZN(
        npu_inst_pe_1_7_6_n116) );
  INV_X1 npu_inst_pe_1_7_6_U9 ( .A(npu_inst_pe_1_7_6_n46), .ZN(
        npu_inst_pe_1_7_6_n115) );
  INV_X1 npu_inst_pe_1_7_6_U8 ( .A(npu_inst_pe_1_7_6_n42), .ZN(
        npu_inst_pe_1_7_6_n114) );
  BUF_X1 npu_inst_pe_1_7_6_U7 ( .A(npu_inst_pe_1_7_6_n11), .Z(
        npu_inst_pe_1_7_6_n10) );
  BUF_X1 npu_inst_pe_1_7_6_U6 ( .A(npu_inst_pe_1_7_6_n11), .Z(
        npu_inst_pe_1_7_6_n9) );
  BUF_X1 npu_inst_pe_1_7_6_U5 ( .A(npu_inst_pe_1_7_6_n11), .Z(
        npu_inst_pe_1_7_6_n8) );
  NOR2_X1 npu_inst_pe_1_7_6_U4 ( .A1(npu_inst_pe_1_7_6_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_6_n1), .ZN(npu_inst_pe_1_7_6_n76) );
  NOR2_X1 npu_inst_pe_1_7_6_U3 ( .A1(npu_inst_pe_1_7_6_n27), .A2(
        npu_inst_pe_1_7_6_n1), .ZN(npu_inst_pe_1_7_6_n77) );
  FA_X1 npu_inst_pe_1_7_6_sub_77_U2_1 ( .A(npu_inst_int_data_res_7__6__1_), 
        .B(npu_inst_pe_1_7_6_n13), .CI(npu_inst_pe_1_7_6_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_7_6_sub_77_carry_2_), .S(npu_inst_pe_1_7_6_N66) );
  FA_X1 npu_inst_pe_1_7_6_add_79_U1_1 ( .A(npu_inst_int_data_res_7__6__1_), 
        .B(npu_inst_pe_1_7_6_int_data_1_), .CI(
        npu_inst_pe_1_7_6_add_79_carry_1_), .CO(
        npu_inst_pe_1_7_6_add_79_carry_2_), .S(npu_inst_pe_1_7_6_N74) );
  NAND3_X1 npu_inst_pe_1_7_6_U101 ( .A1(npu_inst_pe_1_7_6_n4), .A2(
        npu_inst_pe_1_7_6_n6), .A3(npu_inst_pe_1_7_6_n7), .ZN(
        npu_inst_pe_1_7_6_n44) );
  NAND3_X1 npu_inst_pe_1_7_6_U100 ( .A1(npu_inst_pe_1_7_6_n3), .A2(
        npu_inst_pe_1_7_6_n6), .A3(npu_inst_pe_1_7_6_n7), .ZN(
        npu_inst_pe_1_7_6_n40) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_6_n33), .CK(
        npu_inst_pe_1_7_6_net3052), .RN(npu_inst_pe_1_7_6_n8), .Q(
        npu_inst_int_data_res_7__6__6_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_6_n34), .CK(
        npu_inst_pe_1_7_6_net3052), .RN(npu_inst_pe_1_7_6_n8), .Q(
        npu_inst_int_data_res_7__6__5_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_6_n35), .CK(
        npu_inst_pe_1_7_6_net3052), .RN(npu_inst_pe_1_7_6_n8), .Q(
        npu_inst_int_data_res_7__6__4_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_6_n36), .CK(
        npu_inst_pe_1_7_6_net3052), .RN(npu_inst_pe_1_7_6_n8), .Q(
        npu_inst_int_data_res_7__6__3_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_6_n98), .CK(
        npu_inst_pe_1_7_6_net3052), .RN(npu_inst_pe_1_7_6_n8), .Q(
        npu_inst_int_data_res_7__6__2_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_6_n99), .CK(
        npu_inst_pe_1_7_6_net3052), .RN(npu_inst_pe_1_7_6_n8), .Q(
        npu_inst_int_data_res_7__6__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_6_n32), .CK(
        npu_inst_pe_1_7_6_net3052), .RN(npu_inst_pe_1_7_6_n8), .Q(
        npu_inst_int_data_res_7__6__7_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_6_n100), 
        .CK(npu_inst_pe_1_7_6_net3052), .RN(npu_inst_pe_1_7_6_n8), .Q(
        npu_inst_int_data_res_7__6__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_weight_reg_0_ ( .D(npu_inst_n90), .CK(
        npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n8), .Q(
        npu_inst_pe_1_7_6_int_q_weight_0_), .QN(npu_inst_pe_1_7_6_n27) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_weight_reg_1_ ( .D(npu_inst_n96), .CK(
        npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n8), .Q(
        npu_inst_pe_1_7_6_int_q_weight_1_), .QN(npu_inst_pe_1_7_6_n26) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_6_n112), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n8), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_6_n111), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n8), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_6_n110), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_6_n109), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_6_n108), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_6_n107), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_6_n106), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_6_n105), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_6_n104), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_6_n103), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_6_n102), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_6_n101), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_6_n86), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_6_n87), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n9), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_6_n88), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_6_n89), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_6_n90), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_6_n91), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_6_n92), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_6_n93), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_6_n94), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_6_n95), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_6_n96), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_6_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_6_n97), 
        .CK(npu_inst_pe_1_7_6_net3058), .RN(npu_inst_pe_1_7_6_n10), .Q(
        npu_inst_pe_1_7_6_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_6_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_6_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_6_net3052) );
  CLKGATETST_X1 npu_inst_pe_1_7_6_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n43), .SE(1'b0), .GCK(npu_inst_pe_1_7_6_net3058) );
  MUX2_X1 npu_inst_pe_1_7_7_U153 ( .A(npu_inst_pe_1_7_7_n31), .B(
        npu_inst_pe_1_7_7_n28), .S(npu_inst_pe_1_7_7_n7), .Z(
        npu_inst_pe_1_7_7_N93) );
  MUX2_X1 npu_inst_pe_1_7_7_U152 ( .A(npu_inst_pe_1_7_7_n30), .B(
        npu_inst_pe_1_7_7_n29), .S(npu_inst_pe_1_7_7_n5), .Z(
        npu_inst_pe_1_7_7_n31) );
  MUX2_X1 npu_inst_pe_1_7_7_U151 ( .A(npu_inst_pe_1_7_7_int_q_reg_v_0__0_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_v_1__0_), .S(npu_inst_pe_1_7_7_n3), .Z(
        npu_inst_pe_1_7_7_n30) );
  MUX2_X1 npu_inst_pe_1_7_7_U150 ( .A(npu_inst_pe_1_7_7_int_q_reg_v_2__0_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_v_3__0_), .S(npu_inst_pe_1_7_7_n3), .Z(
        npu_inst_pe_1_7_7_n29) );
  MUX2_X1 npu_inst_pe_1_7_7_U149 ( .A(npu_inst_pe_1_7_7_int_q_reg_v_4__0_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_v_5__0_), .S(npu_inst_pe_1_7_7_n3), .Z(
        npu_inst_pe_1_7_7_n28) );
  MUX2_X1 npu_inst_pe_1_7_7_U148 ( .A(npu_inst_pe_1_7_7_n25), .B(
        npu_inst_pe_1_7_7_n22), .S(npu_inst_pe_1_7_7_n7), .Z(
        npu_inst_pe_1_7_7_N94) );
  MUX2_X1 npu_inst_pe_1_7_7_U147 ( .A(npu_inst_pe_1_7_7_n24), .B(
        npu_inst_pe_1_7_7_n23), .S(npu_inst_pe_1_7_7_n5), .Z(
        npu_inst_pe_1_7_7_n25) );
  MUX2_X1 npu_inst_pe_1_7_7_U146 ( .A(npu_inst_pe_1_7_7_int_q_reg_v_0__1_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_v_1__1_), .S(npu_inst_pe_1_7_7_n3), .Z(
        npu_inst_pe_1_7_7_n24) );
  MUX2_X1 npu_inst_pe_1_7_7_U145 ( .A(npu_inst_pe_1_7_7_int_q_reg_v_2__1_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_v_3__1_), .S(npu_inst_pe_1_7_7_n3), .Z(
        npu_inst_pe_1_7_7_n23) );
  MUX2_X1 npu_inst_pe_1_7_7_U144 ( .A(npu_inst_pe_1_7_7_int_q_reg_v_4__1_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_v_5__1_), .S(npu_inst_pe_1_7_7_n3), .Z(
        npu_inst_pe_1_7_7_n22) );
  MUX2_X1 npu_inst_pe_1_7_7_U143 ( .A(npu_inst_pe_1_7_7_n21), .B(
        npu_inst_pe_1_7_7_n18), .S(npu_inst_pe_1_7_7_n7), .Z(
        npu_inst_int_data_x_7__7__1_) );
  MUX2_X1 npu_inst_pe_1_7_7_U142 ( .A(npu_inst_pe_1_7_7_n20), .B(
        npu_inst_pe_1_7_7_n19), .S(npu_inst_pe_1_7_7_n5), .Z(
        npu_inst_pe_1_7_7_n21) );
  MUX2_X1 npu_inst_pe_1_7_7_U141 ( .A(npu_inst_pe_1_7_7_int_q_reg_h_0__1_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_h_1__1_), .S(npu_inst_pe_1_7_7_n3), .Z(
        npu_inst_pe_1_7_7_n20) );
  MUX2_X1 npu_inst_pe_1_7_7_U140 ( .A(npu_inst_pe_1_7_7_int_q_reg_h_2__1_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_h_3__1_), .S(npu_inst_pe_1_7_7_n3), .Z(
        npu_inst_pe_1_7_7_n19) );
  MUX2_X1 npu_inst_pe_1_7_7_U139 ( .A(npu_inst_pe_1_7_7_int_q_reg_h_4__1_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_h_5__1_), .S(npu_inst_pe_1_7_7_n3), .Z(
        npu_inst_pe_1_7_7_n18) );
  MUX2_X1 npu_inst_pe_1_7_7_U138 ( .A(npu_inst_pe_1_7_7_n17), .B(
        npu_inst_pe_1_7_7_n14), .S(npu_inst_pe_1_7_7_n7), .Z(
        npu_inst_int_data_x_7__7__0_) );
  MUX2_X1 npu_inst_pe_1_7_7_U137 ( .A(npu_inst_pe_1_7_7_n16), .B(
        npu_inst_pe_1_7_7_n15), .S(npu_inst_pe_1_7_7_n5), .Z(
        npu_inst_pe_1_7_7_n17) );
  MUX2_X1 npu_inst_pe_1_7_7_U136 ( .A(npu_inst_pe_1_7_7_int_q_reg_h_0__0_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_h_1__0_), .S(npu_inst_pe_1_7_7_n3), .Z(
        npu_inst_pe_1_7_7_n16) );
  MUX2_X1 npu_inst_pe_1_7_7_U135 ( .A(npu_inst_pe_1_7_7_int_q_reg_h_2__0_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_h_3__0_), .S(npu_inst_pe_1_7_7_n3), .Z(
        npu_inst_pe_1_7_7_n15) );
  MUX2_X1 npu_inst_pe_1_7_7_U134 ( .A(npu_inst_pe_1_7_7_int_q_reg_h_4__0_), 
        .B(npu_inst_pe_1_7_7_int_q_reg_h_5__0_), .S(npu_inst_pe_1_7_7_n3), .Z(
        npu_inst_pe_1_7_7_n14) );
  XOR2_X1 npu_inst_pe_1_7_7_U133 ( .A(npu_inst_pe_1_7_7_int_data_0_), .B(
        npu_inst_int_data_res_7__7__0_), .Z(npu_inst_pe_1_7_7_N73) );
  AND2_X1 npu_inst_pe_1_7_7_U132 ( .A1(npu_inst_int_data_res_7__7__0_), .A2(
        npu_inst_pe_1_7_7_int_data_0_), .ZN(npu_inst_pe_1_7_7_add_79_carry_1_)
         );
  XNOR2_X1 npu_inst_pe_1_7_7_U131 ( .A(npu_inst_int_data_res_7__7__0_), .B(
        npu_inst_pe_1_7_7_n12), .ZN(npu_inst_pe_1_7_7_N65) );
  OR2_X1 npu_inst_pe_1_7_7_U130 ( .A1(npu_inst_pe_1_7_7_n12), .A2(
        npu_inst_int_data_res_7__7__0_), .ZN(npu_inst_pe_1_7_7_sub_77_carry_1_) );
  XOR2_X1 npu_inst_pe_1_7_7_U129 ( .A(npu_inst_int_data_res_7__7__2_), .B(
        npu_inst_pe_1_7_7_add_79_carry_2_), .Z(npu_inst_pe_1_7_7_N75) );
  AND2_X1 npu_inst_pe_1_7_7_U128 ( .A1(npu_inst_pe_1_7_7_add_79_carry_2_), 
        .A2(npu_inst_int_data_res_7__7__2_), .ZN(
        npu_inst_pe_1_7_7_add_79_carry_3_) );
  XOR2_X1 npu_inst_pe_1_7_7_U127 ( .A(npu_inst_int_data_res_7__7__3_), .B(
        npu_inst_pe_1_7_7_add_79_carry_3_), .Z(npu_inst_pe_1_7_7_N76) );
  AND2_X1 npu_inst_pe_1_7_7_U126 ( .A1(npu_inst_pe_1_7_7_add_79_carry_3_), 
        .A2(npu_inst_int_data_res_7__7__3_), .ZN(
        npu_inst_pe_1_7_7_add_79_carry_4_) );
  XOR2_X1 npu_inst_pe_1_7_7_U125 ( .A(npu_inst_int_data_res_7__7__4_), .B(
        npu_inst_pe_1_7_7_add_79_carry_4_), .Z(npu_inst_pe_1_7_7_N77) );
  AND2_X1 npu_inst_pe_1_7_7_U124 ( .A1(npu_inst_pe_1_7_7_add_79_carry_4_), 
        .A2(npu_inst_int_data_res_7__7__4_), .ZN(
        npu_inst_pe_1_7_7_add_79_carry_5_) );
  XOR2_X1 npu_inst_pe_1_7_7_U123 ( .A(npu_inst_int_data_res_7__7__5_), .B(
        npu_inst_pe_1_7_7_add_79_carry_5_), .Z(npu_inst_pe_1_7_7_N78) );
  AND2_X1 npu_inst_pe_1_7_7_U122 ( .A1(npu_inst_pe_1_7_7_add_79_carry_5_), 
        .A2(npu_inst_int_data_res_7__7__5_), .ZN(
        npu_inst_pe_1_7_7_add_79_carry_6_) );
  XOR2_X1 npu_inst_pe_1_7_7_U121 ( .A(npu_inst_int_data_res_7__7__6_), .B(
        npu_inst_pe_1_7_7_add_79_carry_6_), .Z(npu_inst_pe_1_7_7_N79) );
  AND2_X1 npu_inst_pe_1_7_7_U120 ( .A1(npu_inst_pe_1_7_7_add_79_carry_6_), 
        .A2(npu_inst_int_data_res_7__7__6_), .ZN(
        npu_inst_pe_1_7_7_add_79_carry_7_) );
  XOR2_X1 npu_inst_pe_1_7_7_U119 ( .A(npu_inst_int_data_res_7__7__7_), .B(
        npu_inst_pe_1_7_7_add_79_carry_7_), .Z(npu_inst_pe_1_7_7_N80) );
  XNOR2_X1 npu_inst_pe_1_7_7_U118 ( .A(npu_inst_pe_1_7_7_sub_77_carry_2_), .B(
        npu_inst_int_data_res_7__7__2_), .ZN(npu_inst_pe_1_7_7_N67) );
  OR2_X1 npu_inst_pe_1_7_7_U117 ( .A1(npu_inst_int_data_res_7__7__2_), .A2(
        npu_inst_pe_1_7_7_sub_77_carry_2_), .ZN(
        npu_inst_pe_1_7_7_sub_77_carry_3_) );
  XNOR2_X1 npu_inst_pe_1_7_7_U116 ( .A(npu_inst_pe_1_7_7_sub_77_carry_3_), .B(
        npu_inst_int_data_res_7__7__3_), .ZN(npu_inst_pe_1_7_7_N68) );
  OR2_X1 npu_inst_pe_1_7_7_U115 ( .A1(npu_inst_int_data_res_7__7__3_), .A2(
        npu_inst_pe_1_7_7_sub_77_carry_3_), .ZN(
        npu_inst_pe_1_7_7_sub_77_carry_4_) );
  XNOR2_X1 npu_inst_pe_1_7_7_U114 ( .A(npu_inst_pe_1_7_7_sub_77_carry_4_), .B(
        npu_inst_int_data_res_7__7__4_), .ZN(npu_inst_pe_1_7_7_N69) );
  OR2_X1 npu_inst_pe_1_7_7_U113 ( .A1(npu_inst_int_data_res_7__7__4_), .A2(
        npu_inst_pe_1_7_7_sub_77_carry_4_), .ZN(
        npu_inst_pe_1_7_7_sub_77_carry_5_) );
  XNOR2_X1 npu_inst_pe_1_7_7_U112 ( .A(npu_inst_pe_1_7_7_sub_77_carry_5_), .B(
        npu_inst_int_data_res_7__7__5_), .ZN(npu_inst_pe_1_7_7_N70) );
  OR2_X1 npu_inst_pe_1_7_7_U111 ( .A1(npu_inst_int_data_res_7__7__5_), .A2(
        npu_inst_pe_1_7_7_sub_77_carry_5_), .ZN(
        npu_inst_pe_1_7_7_sub_77_carry_6_) );
  XNOR2_X1 npu_inst_pe_1_7_7_U110 ( .A(npu_inst_pe_1_7_7_sub_77_carry_6_), .B(
        npu_inst_int_data_res_7__7__6_), .ZN(npu_inst_pe_1_7_7_N71) );
  OR2_X1 npu_inst_pe_1_7_7_U109 ( .A1(npu_inst_int_data_res_7__7__6_), .A2(
        npu_inst_pe_1_7_7_sub_77_carry_6_), .ZN(
        npu_inst_pe_1_7_7_sub_77_carry_7_) );
  XNOR2_X1 npu_inst_pe_1_7_7_U108 ( .A(npu_inst_int_data_res_7__7__7_), .B(
        npu_inst_pe_1_7_7_sub_77_carry_7_), .ZN(npu_inst_pe_1_7_7_N72) );
  INV_X1 npu_inst_pe_1_7_7_U107 ( .A(npu_inst_n57), .ZN(npu_inst_pe_1_7_7_n6)
         );
  INV_X1 npu_inst_pe_1_7_7_U106 ( .A(npu_inst_pe_1_7_7_n6), .ZN(
        npu_inst_pe_1_7_7_n5) );
  INV_X1 npu_inst_pe_1_7_7_U105 ( .A(npu_inst_n34), .ZN(npu_inst_pe_1_7_7_n2)
         );
  AOI22_X1 npu_inst_pe_1_7_7_U104 ( .A1(npu_inst_pe_1_7_7_n38), .A2(
        int_i_data_v_npu[1]), .B1(npu_inst_pe_1_7_7_n113), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_5__1_), .ZN(npu_inst_pe_1_7_7_n39) );
  INV_X1 npu_inst_pe_1_7_7_U103 ( .A(npu_inst_pe_1_7_7_n39), .ZN(
        npu_inst_pe_1_7_7_n111) );
  AOI22_X1 npu_inst_pe_1_7_7_U102 ( .A1(npu_inst_pe_1_7_7_n38), .A2(
        int_i_data_v_npu[0]), .B1(npu_inst_pe_1_7_7_n113), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_5__0_), .ZN(npu_inst_pe_1_7_7_n37) );
  INV_X1 npu_inst_pe_1_7_7_U99 ( .A(npu_inst_pe_1_7_7_n37), .ZN(
        npu_inst_pe_1_7_7_n112) );
  AOI22_X1 npu_inst_pe_1_7_7_U98 ( .A1(int_i_data_v_npu[1]), .A2(
        npu_inst_pe_1_7_7_n58), .B1(npu_inst_pe_1_7_7_n118), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_0__1_), .ZN(npu_inst_pe_1_7_7_n59) );
  INV_X1 npu_inst_pe_1_7_7_U97 ( .A(npu_inst_pe_1_7_7_n59), .ZN(
        npu_inst_pe_1_7_7_n101) );
  AOI22_X1 npu_inst_pe_1_7_7_U96 ( .A1(int_i_data_v_npu[0]), .A2(
        npu_inst_pe_1_7_7_n58), .B1(npu_inst_pe_1_7_7_n118), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_0__0_), .ZN(npu_inst_pe_1_7_7_n57) );
  INV_X1 npu_inst_pe_1_7_7_U95 ( .A(npu_inst_pe_1_7_7_n57), .ZN(
        npu_inst_pe_1_7_7_n102) );
  AOI22_X1 npu_inst_pe_1_7_7_U94 ( .A1(int_i_data_v_npu[1]), .A2(
        npu_inst_pe_1_7_7_n54), .B1(npu_inst_pe_1_7_7_n117), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_1__1_), .ZN(npu_inst_pe_1_7_7_n55) );
  INV_X1 npu_inst_pe_1_7_7_U93 ( .A(npu_inst_pe_1_7_7_n55), .ZN(
        npu_inst_pe_1_7_7_n103) );
  AOI22_X1 npu_inst_pe_1_7_7_U92 ( .A1(int_i_data_v_npu[0]), .A2(
        npu_inst_pe_1_7_7_n54), .B1(npu_inst_pe_1_7_7_n117), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_1__0_), .ZN(npu_inst_pe_1_7_7_n53) );
  INV_X1 npu_inst_pe_1_7_7_U91 ( .A(npu_inst_pe_1_7_7_n53), .ZN(
        npu_inst_pe_1_7_7_n104) );
  AOI22_X1 npu_inst_pe_1_7_7_U90 ( .A1(int_i_data_v_npu[1]), .A2(
        npu_inst_pe_1_7_7_n50), .B1(npu_inst_pe_1_7_7_n116), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_2__1_), .ZN(npu_inst_pe_1_7_7_n51) );
  INV_X1 npu_inst_pe_1_7_7_U89 ( .A(npu_inst_pe_1_7_7_n51), .ZN(
        npu_inst_pe_1_7_7_n105) );
  AOI22_X1 npu_inst_pe_1_7_7_U88 ( .A1(int_i_data_v_npu[0]), .A2(
        npu_inst_pe_1_7_7_n50), .B1(npu_inst_pe_1_7_7_n116), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_2__0_), .ZN(npu_inst_pe_1_7_7_n49) );
  INV_X1 npu_inst_pe_1_7_7_U87 ( .A(npu_inst_pe_1_7_7_n49), .ZN(
        npu_inst_pe_1_7_7_n106) );
  AOI22_X1 npu_inst_pe_1_7_7_U86 ( .A1(int_i_data_v_npu[1]), .A2(
        npu_inst_pe_1_7_7_n46), .B1(npu_inst_pe_1_7_7_n115), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_3__1_), .ZN(npu_inst_pe_1_7_7_n47) );
  INV_X1 npu_inst_pe_1_7_7_U85 ( .A(npu_inst_pe_1_7_7_n47), .ZN(
        npu_inst_pe_1_7_7_n107) );
  AOI22_X1 npu_inst_pe_1_7_7_U84 ( .A1(int_i_data_v_npu[0]), .A2(
        npu_inst_pe_1_7_7_n46), .B1(npu_inst_pe_1_7_7_n115), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_3__0_), .ZN(npu_inst_pe_1_7_7_n45) );
  INV_X1 npu_inst_pe_1_7_7_U83 ( .A(npu_inst_pe_1_7_7_n45), .ZN(
        npu_inst_pe_1_7_7_n108) );
  AOI22_X1 npu_inst_pe_1_7_7_U82 ( .A1(int_i_data_v_npu[1]), .A2(
        npu_inst_pe_1_7_7_n42), .B1(npu_inst_pe_1_7_7_n114), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_4__1_), .ZN(npu_inst_pe_1_7_7_n43) );
  INV_X1 npu_inst_pe_1_7_7_U81 ( .A(npu_inst_pe_1_7_7_n43), .ZN(
        npu_inst_pe_1_7_7_n109) );
  AOI22_X1 npu_inst_pe_1_7_7_U80 ( .A1(int_i_data_v_npu[0]), .A2(
        npu_inst_pe_1_7_7_n42), .B1(npu_inst_pe_1_7_7_n114), .B2(
        npu_inst_pe_1_7_7_int_q_reg_v_4__0_), .ZN(npu_inst_pe_1_7_7_n41) );
  INV_X1 npu_inst_pe_1_7_7_U79 ( .A(npu_inst_pe_1_7_7_n41), .ZN(
        npu_inst_pe_1_7_7_n110) );
  AND2_X1 npu_inst_pe_1_7_7_U78 ( .A1(npu_inst_pe_1_7_7_N93), .A2(npu_inst_n34), .ZN(npu_inst_int_data_y_7__7__0_) );
  AND2_X1 npu_inst_pe_1_7_7_U77 ( .A1(npu_inst_n34), .A2(npu_inst_pe_1_7_7_N94), .ZN(npu_inst_int_data_y_7__7__1_) );
  AOI222_X1 npu_inst_pe_1_7_7_U76 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N73), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N65), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n84) );
  INV_X1 npu_inst_pe_1_7_7_U75 ( .A(npu_inst_pe_1_7_7_n84), .ZN(
        npu_inst_pe_1_7_7_n100) );
  AOI222_X1 npu_inst_pe_1_7_7_U74 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N74), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N66), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n83) );
  INV_X1 npu_inst_pe_1_7_7_U73 ( .A(npu_inst_pe_1_7_7_n83), .ZN(
        npu_inst_pe_1_7_7_n99) );
  AOI222_X1 npu_inst_pe_1_7_7_U72 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N75), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N67), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n82) );
  INV_X1 npu_inst_pe_1_7_7_U71 ( .A(npu_inst_pe_1_7_7_n82), .ZN(
        npu_inst_pe_1_7_7_n98) );
  AOI222_X1 npu_inst_pe_1_7_7_U70 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N76), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N68), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n81) );
  INV_X1 npu_inst_pe_1_7_7_U69 ( .A(npu_inst_pe_1_7_7_n81), .ZN(
        npu_inst_pe_1_7_7_n36) );
  AOI222_X1 npu_inst_pe_1_7_7_U68 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N77), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N69), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n80) );
  INV_X1 npu_inst_pe_1_7_7_U67 ( .A(npu_inst_pe_1_7_7_n80), .ZN(
        npu_inst_pe_1_7_7_n35) );
  AOI222_X1 npu_inst_pe_1_7_7_U66 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N78), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N70), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n79) );
  INV_X1 npu_inst_pe_1_7_7_U65 ( .A(npu_inst_pe_1_7_7_n79), .ZN(
        npu_inst_pe_1_7_7_n34) );
  AOI222_X1 npu_inst_pe_1_7_7_U64 ( .A1(1'b0), .A2(npu_inst_pe_1_7_7_n1), .B1(
        npu_inst_pe_1_7_7_N79), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N71), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n78) );
  INV_X1 npu_inst_pe_1_7_7_U63 ( .A(npu_inst_pe_1_7_7_n78), .ZN(
        npu_inst_pe_1_7_7_n33) );
  AOI222_X1 npu_inst_pe_1_7_7_U62 ( .A1(npu_inst_pe_1_7_7_n1), .A2(1'b0), .B1(
        npu_inst_pe_1_7_7_N80), .B2(npu_inst_pe_1_7_7_n76), .C1(
        npu_inst_pe_1_7_7_N72), .C2(npu_inst_pe_1_7_7_n77), .ZN(
        npu_inst_pe_1_7_7_n75) );
  INV_X1 npu_inst_pe_1_7_7_U61 ( .A(npu_inst_pe_1_7_7_n75), .ZN(
        npu_inst_pe_1_7_7_n32) );
  AND2_X1 npu_inst_pe_1_7_7_U60 ( .A1(npu_inst_int_data_x_7__7__1_), .A2(
        npu_inst_pe_1_7_7_int_q_weight_1_), .ZN(npu_inst_pe_1_7_7_int_data_1_)
         );
  AND2_X1 npu_inst_pe_1_7_7_U59 ( .A1(npu_inst_int_data_x_7__7__0_), .A2(
        npu_inst_pe_1_7_7_int_q_weight_1_), .ZN(npu_inst_pe_1_7_7_int_data_0_)
         );
  INV_X1 npu_inst_pe_1_7_7_U58 ( .A(npu_inst_pe_1_7_7_int_data_1_), .ZN(
        npu_inst_pe_1_7_7_n13) );
  NAND2_X1 npu_inst_pe_1_7_7_U57 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_0__1_), 
        .A2(npu_inst_pe_1_7_7_n60), .ZN(npu_inst_pe_1_7_7_n74) );
  OAI21_X1 npu_inst_pe_1_7_7_U56 ( .B1(npu_inst_pe_1_7_7_n63), .B2(
        npu_inst_pe_1_7_7_n60), .A(npu_inst_pe_1_7_7_n74), .ZN(
        npu_inst_pe_1_7_7_n97) );
  NAND2_X1 npu_inst_pe_1_7_7_U55 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_0__0_), 
        .A2(npu_inst_pe_1_7_7_n60), .ZN(npu_inst_pe_1_7_7_n73) );
  OAI21_X1 npu_inst_pe_1_7_7_U54 ( .B1(npu_inst_pe_1_7_7_n61), .B2(
        npu_inst_pe_1_7_7_n60), .A(npu_inst_pe_1_7_7_n73), .ZN(
        npu_inst_pe_1_7_7_n96) );
  NAND2_X1 npu_inst_pe_1_7_7_U53 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_1__1_), 
        .A2(npu_inst_pe_1_7_7_n56), .ZN(npu_inst_pe_1_7_7_n72) );
  OAI21_X1 npu_inst_pe_1_7_7_U52 ( .B1(npu_inst_pe_1_7_7_n63), .B2(
        npu_inst_pe_1_7_7_n56), .A(npu_inst_pe_1_7_7_n72), .ZN(
        npu_inst_pe_1_7_7_n95) );
  NAND2_X1 npu_inst_pe_1_7_7_U51 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_1__0_), 
        .A2(npu_inst_pe_1_7_7_n56), .ZN(npu_inst_pe_1_7_7_n71) );
  OAI21_X1 npu_inst_pe_1_7_7_U50 ( .B1(npu_inst_pe_1_7_7_n61), .B2(
        npu_inst_pe_1_7_7_n56), .A(npu_inst_pe_1_7_7_n71), .ZN(
        npu_inst_pe_1_7_7_n94) );
  NAND2_X1 npu_inst_pe_1_7_7_U49 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_2__1_), 
        .A2(npu_inst_pe_1_7_7_n52), .ZN(npu_inst_pe_1_7_7_n70) );
  OAI21_X1 npu_inst_pe_1_7_7_U48 ( .B1(npu_inst_pe_1_7_7_n63), .B2(
        npu_inst_pe_1_7_7_n52), .A(npu_inst_pe_1_7_7_n70), .ZN(
        npu_inst_pe_1_7_7_n93) );
  NAND2_X1 npu_inst_pe_1_7_7_U47 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_2__0_), 
        .A2(npu_inst_pe_1_7_7_n52), .ZN(npu_inst_pe_1_7_7_n69) );
  OAI21_X1 npu_inst_pe_1_7_7_U46 ( .B1(npu_inst_pe_1_7_7_n61), .B2(
        npu_inst_pe_1_7_7_n52), .A(npu_inst_pe_1_7_7_n69), .ZN(
        npu_inst_pe_1_7_7_n92) );
  NAND2_X1 npu_inst_pe_1_7_7_U45 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_3__1_), 
        .A2(npu_inst_pe_1_7_7_n48), .ZN(npu_inst_pe_1_7_7_n68) );
  OAI21_X1 npu_inst_pe_1_7_7_U44 ( .B1(npu_inst_pe_1_7_7_n63), .B2(
        npu_inst_pe_1_7_7_n48), .A(npu_inst_pe_1_7_7_n68), .ZN(
        npu_inst_pe_1_7_7_n91) );
  NAND2_X1 npu_inst_pe_1_7_7_U43 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_3__0_), 
        .A2(npu_inst_pe_1_7_7_n48), .ZN(npu_inst_pe_1_7_7_n67) );
  OAI21_X1 npu_inst_pe_1_7_7_U42 ( .B1(npu_inst_pe_1_7_7_n61), .B2(
        npu_inst_pe_1_7_7_n48), .A(npu_inst_pe_1_7_7_n67), .ZN(
        npu_inst_pe_1_7_7_n90) );
  NAND2_X1 npu_inst_pe_1_7_7_U41 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_4__1_), 
        .A2(npu_inst_pe_1_7_7_n44), .ZN(npu_inst_pe_1_7_7_n66) );
  OAI21_X1 npu_inst_pe_1_7_7_U40 ( .B1(npu_inst_pe_1_7_7_n63), .B2(
        npu_inst_pe_1_7_7_n44), .A(npu_inst_pe_1_7_7_n66), .ZN(
        npu_inst_pe_1_7_7_n89) );
  NAND2_X1 npu_inst_pe_1_7_7_U39 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_4__0_), 
        .A2(npu_inst_pe_1_7_7_n44), .ZN(npu_inst_pe_1_7_7_n65) );
  OAI21_X1 npu_inst_pe_1_7_7_U38 ( .B1(npu_inst_pe_1_7_7_n61), .B2(
        npu_inst_pe_1_7_7_n44), .A(npu_inst_pe_1_7_7_n65), .ZN(
        npu_inst_pe_1_7_7_n88) );
  NAND2_X1 npu_inst_pe_1_7_7_U37 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_5__1_), 
        .A2(npu_inst_pe_1_7_7_n40), .ZN(npu_inst_pe_1_7_7_n64) );
  OAI21_X1 npu_inst_pe_1_7_7_U36 ( .B1(npu_inst_pe_1_7_7_n63), .B2(
        npu_inst_pe_1_7_7_n40), .A(npu_inst_pe_1_7_7_n64), .ZN(
        npu_inst_pe_1_7_7_n87) );
  NAND2_X1 npu_inst_pe_1_7_7_U35 ( .A1(npu_inst_pe_1_7_7_int_q_reg_h_5__0_), 
        .A2(npu_inst_pe_1_7_7_n40), .ZN(npu_inst_pe_1_7_7_n62) );
  OAI21_X1 npu_inst_pe_1_7_7_U34 ( .B1(npu_inst_pe_1_7_7_n61), .B2(
        npu_inst_pe_1_7_7_n40), .A(npu_inst_pe_1_7_7_n62), .ZN(
        npu_inst_pe_1_7_7_n86) );
  NOR3_X1 npu_inst_pe_1_7_7_U33 ( .A1(npu_inst_pe_1_7_7_n26), .A2(npu_inst_n34), .A3(npu_inst_int_ckg[0]), .ZN(npu_inst_pe_1_7_7_n85) );
  OR2_X1 npu_inst_pe_1_7_7_U32 ( .A1(npu_inst_pe_1_7_7_n85), .A2(
        npu_inst_pe_1_7_7_n1), .ZN(npu_inst_pe_1_7_7_N84) );
  AOI22_X1 npu_inst_pe_1_7_7_U31 ( .A1(npu_inst_n34), .A2(int_i_data_v_npu[1]), 
        .B1(npu_inst_pe_1_7_7_n2), .B2(int_i_data_h_npu[1]), .ZN(
        npu_inst_pe_1_7_7_n63) );
  AOI22_X1 npu_inst_pe_1_7_7_U30 ( .A1(npu_inst_n34), .A2(int_i_data_v_npu[0]), 
        .B1(npu_inst_pe_1_7_7_n2), .B2(int_i_data_h_npu[0]), .ZN(
        npu_inst_pe_1_7_7_n61) );
  INV_X1 npu_inst_pe_1_7_7_U29 ( .A(npu_inst_pe_1_7_7_int_data_0_), .ZN(
        npu_inst_pe_1_7_7_n12) );
  INV_X1 npu_inst_pe_1_7_7_U28 ( .A(npu_inst_n49), .ZN(npu_inst_pe_1_7_7_n4)
         );
  OR3_X1 npu_inst_pe_1_7_7_U27 ( .A1(npu_inst_pe_1_7_7_n5), .A2(
        npu_inst_pe_1_7_7_n7), .A3(npu_inst_pe_1_7_7_n4), .ZN(
        npu_inst_pe_1_7_7_n56) );
  OR3_X1 npu_inst_pe_1_7_7_U26 ( .A1(npu_inst_pe_1_7_7_n4), .A2(
        npu_inst_pe_1_7_7_n7), .A3(npu_inst_pe_1_7_7_n6), .ZN(
        npu_inst_pe_1_7_7_n48) );
  INV_X1 npu_inst_pe_1_7_7_U25 ( .A(npu_inst_pe_1_7_7_n4), .ZN(
        npu_inst_pe_1_7_7_n3) );
  OR3_X1 npu_inst_pe_1_7_7_U24 ( .A1(npu_inst_pe_1_7_7_n3), .A2(
        npu_inst_pe_1_7_7_n7), .A3(npu_inst_pe_1_7_7_n6), .ZN(
        npu_inst_pe_1_7_7_n52) );
  OR3_X1 npu_inst_pe_1_7_7_U23 ( .A1(npu_inst_pe_1_7_7_n5), .A2(
        npu_inst_pe_1_7_7_n7), .A3(npu_inst_pe_1_7_7_n3), .ZN(
        npu_inst_pe_1_7_7_n60) );
  BUF_X1 npu_inst_pe_1_7_7_U22 ( .A(npu_inst_n11), .Z(npu_inst_pe_1_7_7_n1) );
  NOR2_X1 npu_inst_pe_1_7_7_U21 ( .A1(npu_inst_pe_1_7_7_n60), .A2(
        npu_inst_pe_1_7_7_n2), .ZN(npu_inst_pe_1_7_7_n58) );
  NOR2_X1 npu_inst_pe_1_7_7_U20 ( .A1(npu_inst_pe_1_7_7_n56), .A2(
        npu_inst_pe_1_7_7_n2), .ZN(npu_inst_pe_1_7_7_n54) );
  NOR2_X1 npu_inst_pe_1_7_7_U19 ( .A1(npu_inst_pe_1_7_7_n52), .A2(
        npu_inst_pe_1_7_7_n2), .ZN(npu_inst_pe_1_7_7_n50) );
  NOR2_X1 npu_inst_pe_1_7_7_U18 ( .A1(npu_inst_pe_1_7_7_n48), .A2(
        npu_inst_pe_1_7_7_n2), .ZN(npu_inst_pe_1_7_7_n46) );
  NOR2_X1 npu_inst_pe_1_7_7_U17 ( .A1(npu_inst_pe_1_7_7_n40), .A2(
        npu_inst_pe_1_7_7_n2), .ZN(npu_inst_pe_1_7_7_n38) );
  NOR2_X1 npu_inst_pe_1_7_7_U16 ( .A1(npu_inst_pe_1_7_7_n44), .A2(
        npu_inst_pe_1_7_7_n2), .ZN(npu_inst_pe_1_7_7_n42) );
  BUF_X1 npu_inst_pe_1_7_7_U15 ( .A(npu_inst_n74), .Z(npu_inst_pe_1_7_7_n7) );
  INV_X1 npu_inst_pe_1_7_7_U14 ( .A(npu_inst_n104), .ZN(npu_inst_pe_1_7_7_n11)
         );
  INV_X1 npu_inst_pe_1_7_7_U13 ( .A(npu_inst_pe_1_7_7_n38), .ZN(
        npu_inst_pe_1_7_7_n113) );
  INV_X1 npu_inst_pe_1_7_7_U12 ( .A(npu_inst_pe_1_7_7_n58), .ZN(
        npu_inst_pe_1_7_7_n118) );
  INV_X1 npu_inst_pe_1_7_7_U11 ( .A(npu_inst_pe_1_7_7_n54), .ZN(
        npu_inst_pe_1_7_7_n117) );
  INV_X1 npu_inst_pe_1_7_7_U10 ( .A(npu_inst_pe_1_7_7_n50), .ZN(
        npu_inst_pe_1_7_7_n116) );
  INV_X1 npu_inst_pe_1_7_7_U9 ( .A(npu_inst_pe_1_7_7_n46), .ZN(
        npu_inst_pe_1_7_7_n115) );
  INV_X1 npu_inst_pe_1_7_7_U8 ( .A(npu_inst_pe_1_7_7_n42), .ZN(
        npu_inst_pe_1_7_7_n114) );
  BUF_X1 npu_inst_pe_1_7_7_U7 ( .A(npu_inst_pe_1_7_7_n11), .Z(
        npu_inst_pe_1_7_7_n10) );
  BUF_X1 npu_inst_pe_1_7_7_U6 ( .A(npu_inst_pe_1_7_7_n11), .Z(
        npu_inst_pe_1_7_7_n9) );
  BUF_X1 npu_inst_pe_1_7_7_U5 ( .A(npu_inst_pe_1_7_7_n11), .Z(
        npu_inst_pe_1_7_7_n8) );
  NOR2_X1 npu_inst_pe_1_7_7_U4 ( .A1(npu_inst_pe_1_7_7_int_q_weight_0_), .A2(
        npu_inst_pe_1_7_7_n1), .ZN(npu_inst_pe_1_7_7_n76) );
  NOR2_X1 npu_inst_pe_1_7_7_U3 ( .A1(npu_inst_pe_1_7_7_n27), .A2(
        npu_inst_pe_1_7_7_n1), .ZN(npu_inst_pe_1_7_7_n77) );
  FA_X1 npu_inst_pe_1_7_7_sub_77_U2_1 ( .A(npu_inst_int_data_res_7__7__1_), 
        .B(npu_inst_pe_1_7_7_n13), .CI(npu_inst_pe_1_7_7_sub_77_carry_1_), 
        .CO(npu_inst_pe_1_7_7_sub_77_carry_2_), .S(npu_inst_pe_1_7_7_N66) );
  FA_X1 npu_inst_pe_1_7_7_add_79_U1_1 ( .A(npu_inst_int_data_res_7__7__1_), 
        .B(npu_inst_pe_1_7_7_int_data_1_), .CI(
        npu_inst_pe_1_7_7_add_79_carry_1_), .CO(
        npu_inst_pe_1_7_7_add_79_carry_2_), .S(npu_inst_pe_1_7_7_N74) );
  NAND3_X1 npu_inst_pe_1_7_7_U101 ( .A1(npu_inst_pe_1_7_7_n4), .A2(
        npu_inst_pe_1_7_7_n6), .A3(npu_inst_pe_1_7_7_n7), .ZN(
        npu_inst_pe_1_7_7_n44) );
  NAND3_X1 npu_inst_pe_1_7_7_U100 ( .A1(npu_inst_pe_1_7_7_n3), .A2(
        npu_inst_pe_1_7_7_n6), .A3(npu_inst_pe_1_7_7_n7), .ZN(
        npu_inst_pe_1_7_7_n40) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_6_ ( .D(npu_inst_pe_1_7_7_n33), .CK(
        npu_inst_pe_1_7_7_net3029), .RN(npu_inst_pe_1_7_7_n8), .Q(
        npu_inst_int_data_res_7__7__6_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_5_ ( .D(npu_inst_pe_1_7_7_n34), .CK(
        npu_inst_pe_1_7_7_net3029), .RN(npu_inst_pe_1_7_7_n8), .Q(
        npu_inst_int_data_res_7__7__5_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_4_ ( .D(npu_inst_pe_1_7_7_n35), .CK(
        npu_inst_pe_1_7_7_net3029), .RN(npu_inst_pe_1_7_7_n8), .Q(
        npu_inst_int_data_res_7__7__4_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_3_ ( .D(npu_inst_pe_1_7_7_n36), .CK(
        npu_inst_pe_1_7_7_net3029), .RN(npu_inst_pe_1_7_7_n8), .Q(
        npu_inst_int_data_res_7__7__3_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_2_ ( .D(npu_inst_pe_1_7_7_n98), .CK(
        npu_inst_pe_1_7_7_net3029), .RN(npu_inst_pe_1_7_7_n8), .Q(
        npu_inst_int_data_res_7__7__2_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_1_ ( .D(npu_inst_pe_1_7_7_n99), .CK(
        npu_inst_pe_1_7_7_net3029), .RN(npu_inst_pe_1_7_7_n8), .Q(
        npu_inst_int_data_res_7__7__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_7_ ( .D(npu_inst_pe_1_7_7_n32), .CK(
        npu_inst_pe_1_7_7_net3029), .RN(npu_inst_pe_1_7_7_n8), .Q(
        npu_inst_int_data_res_7__7__7_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_acc_reg_0_ ( .D(npu_inst_pe_1_7_7_n100), 
        .CK(npu_inst_pe_1_7_7_net3029), .RN(npu_inst_pe_1_7_7_n8), .Q(
        npu_inst_int_data_res_7__7__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_weight_reg_0_ ( .D(npu_inst_n90), .CK(
        npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n8), .Q(
        npu_inst_pe_1_7_7_int_q_weight_0_), .QN(npu_inst_pe_1_7_7_n27) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_weight_reg_1_ ( .D(npu_inst_n96), .CK(
        npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n8), .Q(
        npu_inst_pe_1_7_7_int_q_weight_1_), .QN(npu_inst_pe_1_7_7_n26) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_5__0_ ( .D(npu_inst_pe_1_7_7_n112), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n8), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_5__1_ ( .D(npu_inst_pe_1_7_7_n111), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n8), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_4__0_ ( .D(npu_inst_pe_1_7_7_n110), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_4__1_ ( .D(npu_inst_pe_1_7_7_n109), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_3__0_ ( .D(npu_inst_pe_1_7_7_n108), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_3__1_ ( .D(npu_inst_pe_1_7_7_n107), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_2__0_ ( .D(npu_inst_pe_1_7_7_n106), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_2__1_ ( .D(npu_inst_pe_1_7_7_n105), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_1__0_ ( .D(npu_inst_pe_1_7_7_n104), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_1__1_ ( .D(npu_inst_pe_1_7_7_n103), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_0__0_ ( .D(npu_inst_pe_1_7_7_n102), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_v_reg_0__1_ ( .D(npu_inst_pe_1_7_7_n101), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_reg_v_0__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_5__0_ ( .D(npu_inst_pe_1_7_7_n86), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_5__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_5__1_ ( .D(npu_inst_pe_1_7_7_n87), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n9), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_5__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_4__0_ ( .D(npu_inst_pe_1_7_7_n88), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_4__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_4__1_ ( .D(npu_inst_pe_1_7_7_n89), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_4__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_3__0_ ( .D(npu_inst_pe_1_7_7_n90), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_3__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_3__1_ ( .D(npu_inst_pe_1_7_7_n91), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_3__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_2__0_ ( .D(npu_inst_pe_1_7_7_n92), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_2__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_2__1_ ( .D(npu_inst_pe_1_7_7_n93), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_2__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_1__0_ ( .D(npu_inst_pe_1_7_7_n94), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_1__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_1__1_ ( .D(npu_inst_pe_1_7_7_n95), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_1__1_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_0__0_ ( .D(npu_inst_pe_1_7_7_n96), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_0__0_) );
  DFFR_X1 npu_inst_pe_1_7_7_int_q_reg_h_reg_0__1_ ( .D(npu_inst_pe_1_7_7_n97), 
        .CK(npu_inst_pe_1_7_7_net3035), .RN(npu_inst_pe_1_7_7_n10), .Q(
        npu_inst_pe_1_7_7_int_q_reg_h_0__1_) );
  CLKGATETST_X1 npu_inst_pe_1_7_7_clk_gate_int_q_acc_reg_latch ( .CK(ck), .E(
        npu_inst_pe_1_7_7_N84), .SE(1'b0), .GCK(npu_inst_pe_1_7_7_net3029) );
  CLKGATETST_X1 npu_inst_pe_1_7_7_clk_gate_int_q_reg_h_reg_0__latch ( .CK(ck), 
        .E(npu_inst_n43), .SE(1'b0), .GCK(npu_inst_pe_1_7_7_net3035) );
  OR3_X1 qrelu_i_0_U8 ( .A1(int_o_data_npu[62]), .A2(int_o_data_npu[61]), .A3(
        int_o_data_npu[60]), .ZN(qrelu_i_0_n5) );
  OR2_X1 qrelu_i_0_U7 ( .A1(int_o_data_npu[59]), .A2(int_o_data_npu[58]), .ZN(
        qrelu_i_0_n6) );
  INV_X1 qrelu_i_0_U6 ( .A(int_o_data_npu[63]), .ZN(qrelu_i_0_n2) );
  OAI21_X1 qrelu_i_0_U5 ( .B1(qrelu_i_0_n5), .B2(qrelu_i_0_n6), .A(
        qrelu_i_0_n2), .ZN(qrelu_i_0_n4) );
  INV_X1 qrelu_i_0_U4 ( .A(int_o_data_npu[57]), .ZN(qrelu_i_0_n3) );
  OAI21_X1 qrelu_i_0_U3 ( .B1(qrelu_i_0_n3), .B2(int_o_data_npu[63]), .A(
        qrelu_i_0_n4), .ZN(o_data_relu[15]) );
  INV_X1 qrelu_i_0_U2 ( .A(int_o_data_npu[56]), .ZN(qrelu_i_0_n1) );
  OAI21_X1 qrelu_i_0_U1 ( .B1(qrelu_i_0_n1), .B2(int_o_data_npu[63]), .A(
        qrelu_i_0_n4), .ZN(o_data_relu[14]) );
  OR3_X1 qrelu_i_1_U8 ( .A1(int_o_data_npu[54]), .A2(int_o_data_npu[53]), .A3(
        int_o_data_npu[52]), .ZN(qrelu_i_1_n8) );
  OR2_X1 qrelu_i_1_U7 ( .A1(int_o_data_npu[51]), .A2(int_o_data_npu[50]), .ZN(
        qrelu_i_1_n7) );
  INV_X1 qrelu_i_1_U6 ( .A(int_o_data_npu[55]), .ZN(qrelu_i_1_n2) );
  OAI21_X1 qrelu_i_1_U5 ( .B1(qrelu_i_1_n8), .B2(qrelu_i_1_n7), .A(
        qrelu_i_1_n2), .ZN(qrelu_i_1_n9) );
  INV_X1 qrelu_i_1_U4 ( .A(int_o_data_npu[49]), .ZN(qrelu_i_1_n3) );
  OAI21_X1 qrelu_i_1_U3 ( .B1(qrelu_i_1_n3), .B2(int_o_data_npu[55]), .A(
        qrelu_i_1_n9), .ZN(o_data_relu[13]) );
  INV_X1 qrelu_i_1_U2 ( .A(int_o_data_npu[48]), .ZN(qrelu_i_1_n1) );
  OAI21_X1 qrelu_i_1_U1 ( .B1(qrelu_i_1_n1), .B2(int_o_data_npu[55]), .A(
        qrelu_i_1_n9), .ZN(o_data_relu[12]) );
  OR3_X1 qrelu_i_2_U8 ( .A1(int_o_data_npu[46]), .A2(int_o_data_npu[45]), .A3(
        int_o_data_npu[44]), .ZN(qrelu_i_2_n8) );
  OR2_X1 qrelu_i_2_U7 ( .A1(int_o_data_npu[43]), .A2(int_o_data_npu[42]), .ZN(
        qrelu_i_2_n7) );
  INV_X1 qrelu_i_2_U6 ( .A(int_o_data_npu[47]), .ZN(qrelu_i_2_n2) );
  OAI21_X1 qrelu_i_2_U5 ( .B1(qrelu_i_2_n8), .B2(qrelu_i_2_n7), .A(
        qrelu_i_2_n2), .ZN(qrelu_i_2_n9) );
  INV_X1 qrelu_i_2_U4 ( .A(int_o_data_npu[41]), .ZN(qrelu_i_2_n3) );
  OAI21_X1 qrelu_i_2_U3 ( .B1(qrelu_i_2_n3), .B2(int_o_data_npu[47]), .A(
        qrelu_i_2_n9), .ZN(o_data_relu[11]) );
  INV_X1 qrelu_i_2_U2 ( .A(int_o_data_npu[40]), .ZN(qrelu_i_2_n1) );
  OAI21_X1 qrelu_i_2_U1 ( .B1(qrelu_i_2_n1), .B2(int_o_data_npu[47]), .A(
        qrelu_i_2_n9), .ZN(o_data_relu[10]) );
  OR3_X1 qrelu_i_3_U8 ( .A1(int_o_data_npu[38]), .A2(int_o_data_npu[37]), .A3(
        int_o_data_npu[36]), .ZN(qrelu_i_3_n8) );
  OR2_X1 qrelu_i_3_U7 ( .A1(int_o_data_npu[35]), .A2(int_o_data_npu[34]), .ZN(
        qrelu_i_3_n7) );
  INV_X1 qrelu_i_3_U6 ( .A(int_o_data_npu[39]), .ZN(qrelu_i_3_n2) );
  OAI21_X1 qrelu_i_3_U5 ( .B1(qrelu_i_3_n8), .B2(qrelu_i_3_n7), .A(
        qrelu_i_3_n2), .ZN(qrelu_i_3_n9) );
  INV_X1 qrelu_i_3_U4 ( .A(int_o_data_npu[33]), .ZN(qrelu_i_3_n3) );
  OAI21_X1 qrelu_i_3_U3 ( .B1(qrelu_i_3_n3), .B2(int_o_data_npu[39]), .A(
        qrelu_i_3_n9), .ZN(o_data_relu[9]) );
  INV_X1 qrelu_i_3_U2 ( .A(int_o_data_npu[32]), .ZN(qrelu_i_3_n1) );
  OAI21_X1 qrelu_i_3_U1 ( .B1(qrelu_i_3_n1), .B2(int_o_data_npu[39]), .A(
        qrelu_i_3_n9), .ZN(o_data_relu[8]) );
  OR3_X1 qrelu_i_4_U8 ( .A1(int_o_data_npu[30]), .A2(int_o_data_npu[29]), .A3(
        int_o_data_npu[28]), .ZN(qrelu_i_4_n8) );
  OR2_X1 qrelu_i_4_U7 ( .A1(int_o_data_npu[27]), .A2(int_o_data_npu[26]), .ZN(
        qrelu_i_4_n7) );
  INV_X1 qrelu_i_4_U6 ( .A(int_o_data_npu[31]), .ZN(qrelu_i_4_n2) );
  OAI21_X1 qrelu_i_4_U5 ( .B1(qrelu_i_4_n8), .B2(qrelu_i_4_n7), .A(
        qrelu_i_4_n2), .ZN(qrelu_i_4_n9) );
  INV_X1 qrelu_i_4_U4 ( .A(int_o_data_npu[25]), .ZN(qrelu_i_4_n3) );
  OAI21_X1 qrelu_i_4_U3 ( .B1(qrelu_i_4_n3), .B2(int_o_data_npu[31]), .A(
        qrelu_i_4_n9), .ZN(o_data_relu[7]) );
  INV_X1 qrelu_i_4_U2 ( .A(int_o_data_npu[24]), .ZN(qrelu_i_4_n1) );
  OAI21_X1 qrelu_i_4_U1 ( .B1(qrelu_i_4_n1), .B2(int_o_data_npu[31]), .A(
        qrelu_i_4_n9), .ZN(o_data_relu[6]) );
  OR3_X1 qrelu_i_5_U8 ( .A1(int_o_data_npu[22]), .A2(int_o_data_npu[21]), .A3(
        int_o_data_npu[20]), .ZN(qrelu_i_5_n8) );
  OR2_X1 qrelu_i_5_U7 ( .A1(int_o_data_npu[19]), .A2(int_o_data_npu[18]), .ZN(
        qrelu_i_5_n7) );
  INV_X1 qrelu_i_5_U6 ( .A(int_o_data_npu[23]), .ZN(qrelu_i_5_n2) );
  OAI21_X1 qrelu_i_5_U5 ( .B1(qrelu_i_5_n8), .B2(qrelu_i_5_n7), .A(
        qrelu_i_5_n2), .ZN(qrelu_i_5_n9) );
  INV_X1 qrelu_i_5_U4 ( .A(int_o_data_npu[17]), .ZN(qrelu_i_5_n3) );
  OAI21_X1 qrelu_i_5_U3 ( .B1(qrelu_i_5_n3), .B2(int_o_data_npu[23]), .A(
        qrelu_i_5_n9), .ZN(o_data_relu[5]) );
  INV_X1 qrelu_i_5_U2 ( .A(int_o_data_npu[16]), .ZN(qrelu_i_5_n1) );
  OAI21_X1 qrelu_i_5_U1 ( .B1(qrelu_i_5_n1), .B2(int_o_data_npu[23]), .A(
        qrelu_i_5_n9), .ZN(o_data_relu[4]) );
  OR3_X1 qrelu_i_6_U8 ( .A1(int_o_data_npu[14]), .A2(int_o_data_npu[13]), .A3(
        int_o_data_npu[12]), .ZN(qrelu_i_6_n8) );
  OR2_X1 qrelu_i_6_U7 ( .A1(int_o_data_npu[11]), .A2(int_o_data_npu[10]), .ZN(
        qrelu_i_6_n7) );
  INV_X1 qrelu_i_6_U6 ( .A(int_o_data_npu[15]), .ZN(qrelu_i_6_n2) );
  OAI21_X1 qrelu_i_6_U5 ( .B1(qrelu_i_6_n8), .B2(qrelu_i_6_n7), .A(
        qrelu_i_6_n2), .ZN(qrelu_i_6_n9) );
  INV_X1 qrelu_i_6_U4 ( .A(int_o_data_npu[9]), .ZN(qrelu_i_6_n3) );
  OAI21_X1 qrelu_i_6_U3 ( .B1(qrelu_i_6_n3), .B2(int_o_data_npu[15]), .A(
        qrelu_i_6_n9), .ZN(o_data_relu[3]) );
  INV_X1 qrelu_i_6_U2 ( .A(int_o_data_npu[8]), .ZN(qrelu_i_6_n1) );
  OAI21_X1 qrelu_i_6_U1 ( .B1(qrelu_i_6_n1), .B2(int_o_data_npu[15]), .A(
        qrelu_i_6_n9), .ZN(o_data_relu[2]) );
  OR3_X1 qrelu_i_7_U8 ( .A1(int_o_data_npu[6]), .A2(int_o_data_npu[5]), .A3(
        int_o_data_npu[4]), .ZN(qrelu_i_7_n8) );
  OR2_X1 qrelu_i_7_U7 ( .A1(int_o_data_npu[3]), .A2(int_o_data_npu[2]), .ZN(
        qrelu_i_7_n7) );
  INV_X1 qrelu_i_7_U6 ( .A(int_o_data_npu[7]), .ZN(qrelu_i_7_n2) );
  OAI21_X1 qrelu_i_7_U5 ( .B1(qrelu_i_7_n8), .B2(qrelu_i_7_n7), .A(
        qrelu_i_7_n2), .ZN(qrelu_i_7_n9) );
  INV_X1 qrelu_i_7_U4 ( .A(int_o_data_npu[1]), .ZN(qrelu_i_7_n3) );
  OAI21_X1 qrelu_i_7_U3 ( .B1(qrelu_i_7_n3), .B2(int_o_data_npu[7]), .A(
        qrelu_i_7_n9), .ZN(o_data_relu[1]) );
  INV_X1 qrelu_i_7_U2 ( .A(int_o_data_npu[0]), .ZN(qrelu_i_7_n1) );
  OAI21_X1 qrelu_i_7_U1 ( .B1(qrelu_i_7_n1), .B2(int_o_data_npu[7]), .A(
        qrelu_i_7_n9), .ZN(o_data_relu[0]) );
  INV_X1 p_unit_i_0_U18 ( .A(n48), .ZN(p_unit_i_0_n11) );
  INV_X1 p_unit_i_0_U17 ( .A(p_unit_i_0_n8), .ZN(p_unit_i_0_n16) );
  NOR2_X1 p_unit_i_0_U15 ( .A1(p_unit_i_0_int_ps0_2_), .A2(p_unit_i_0_n16), 
        .ZN(p_unit_i_0_n6) );
  OAI22_X1 p_unit_i_0_U14 ( .A1(p_unit_i_0_n8), .A2(p_unit_i_0_n5), .B1(
        p_unit_i_0_n6), .B2(p_unit_i_0_n7), .ZN(p_unit_i_0_n4) );
  XNOR2_X1 p_unit_i_0_U13 ( .A(p_unit_i_0_n8), .B(p_unit_i_0_n9), .ZN(
        p_unit_i_0_N7) );
  XNOR2_X1 p_unit_i_0_U12 ( .A(p_unit_i_0_int_ps1_1_), .B(
        p_unit_i_0_int_ps0_1_), .ZN(p_unit_i_0_n3) );
  NAND2_X1 p_unit_i_0_U11 ( .A1(p_unit_i_0_int_ps0_0_), .A2(
        p_unit_i_0_int_ps1_0_), .ZN(p_unit_i_0_n2) );
  XOR2_X1 p_unit_i_0_U10 ( .A(p_unit_i_0_n2), .B(p_unit_i_0_n3), .Z(
        p_unit_i_0_N6) );
  OAI211_X1 p_unit_i_0_U9 ( .C1(p_unit_i_0_int_ps0_1_), .C2(
        p_unit_i_0_int_ps1_1_), .A(p_unit_i_0_int_ps0_0_), .B(
        p_unit_i_0_int_ps1_0_), .ZN(p_unit_i_0_n10) );
  INV_X1 p_unit_i_0_U8 ( .A(p_unit_i_0_n10), .ZN(p_unit_i_0_n17) );
  AOI21_X1 p_unit_i_0_U7 ( .B1(p_unit_i_0_int_ps0_1_), .B2(
        p_unit_i_0_int_ps1_1_), .A(p_unit_i_0_n17), .ZN(p_unit_i_0_n8) );
  AND3_X1 p_unit_i_0_U6 ( .A1(o_data_relu[14]), .A2(p_unit_i_0_n15), .A3(
        o_data_relu[12]), .ZN(p_unit_i_0_n14) );
  AOI21_X1 p_unit_i_0_U5 ( .B1(o_data_relu[13]), .B2(o_data_relu[15]), .A(
        p_unit_i_0_n14), .ZN(p_unit_i_0_n13) );
  INV_X1 p_unit_i_0_U4 ( .A(p_unit_i_0_n13), .ZN(p_unit_i_0_n12) );
  NAND2_X1 p_unit_i_0_U3 ( .A1(o_data_relu[14]), .A2(o_data_relu[12]), .ZN(
        p_unit_i_0_n1) );
  XNOR2_X1 p_unit_i_0_U2 ( .A(p_unit_i_0_n1), .B(p_unit_i_0_n15), .ZN(
        p_unit_i_0_N3) );
  XOR2_X1 p_unit_i_0_U22 ( .A(o_data_relu[12]), .B(o_data_relu[14]), .Z(
        p_unit_i_0_N2) );
  XOR2_X1 p_unit_i_0_U21 ( .A(o_data_relu[15]), .B(o_data_relu[13]), .Z(
        p_unit_i_0_n15) );
  XOR2_X1 p_unit_i_0_U19 ( .A(p_unit_i_0_int_ps1_0_), .B(p_unit_i_0_int_ps0_0_), .Z(p_unit_i_0_N5) );
  XOR2_X1 p_unit_i_0_U16 ( .A(p_unit_i_0_int_ps1_2_), .B(p_unit_i_0_int_ps0_2_), .Z(p_unit_i_0_n9) );
  DFFR_X1 p_unit_i_0_o_data_reg_1_ ( .D(p_unit_i_0_N6), .CK(p_unit_i_0_net3011), .RN(p_unit_i_0_n11), .Q(int_o_data_p[13]) );
  DFFR_X1 p_unit_i_0_o_data_reg_2_ ( .D(p_unit_i_0_N7), .CK(p_unit_i_0_net3011), .RN(p_unit_i_0_n11), .Q(int_o_data_p[14]) );
  DFFR_X1 p_unit_i_0_o_data_reg_3_ ( .D(p_unit_i_0_n4), .CK(p_unit_i_0_net3011), .RN(p_unit_i_0_n11), .Q(int_o_data_p[15]) );
  DFFR_X1 p_unit_i_0_o_data_reg_0_ ( .D(p_unit_i_0_N5), .CK(p_unit_i_0_net3011), .RN(p_unit_i_0_n11), .Q(int_o_data_p[12]) );
  DFFR_X1 p_unit_i_0_int_ps1_reg_0_ ( .D(p_unit_i_0_int_ps0_0_), .CK(
        p_unit_i_0_net3011), .RN(p_unit_i_0_n11), .Q(p_unit_i_0_int_ps1_0_) );
  DFFR_X1 p_unit_i_0_int_ps1_reg_1_ ( .D(p_unit_i_0_int_ps0_1_), .CK(
        p_unit_i_0_net3011), .RN(p_unit_i_0_n11), .Q(p_unit_i_0_int_ps1_1_) );
  DFFR_X1 p_unit_i_0_int_ps1_reg_2_ ( .D(p_unit_i_0_int_ps0_2_), .CK(
        p_unit_i_0_net3011), .RN(p_unit_i_0_n11), .Q(p_unit_i_0_int_ps1_2_), 
        .QN(p_unit_i_0_n7) );
  DFFR_X1 p_unit_i_0_int_ps0_reg_0_ ( .D(p_unit_i_0_N2), .CK(
        p_unit_i_0_net3011), .RN(p_unit_i_0_n11), .Q(p_unit_i_0_int_ps0_0_) );
  DFFR_X1 p_unit_i_0_int_ps0_reg_1_ ( .D(p_unit_i_0_N3), .CK(
        p_unit_i_0_net3011), .RN(p_unit_i_0_n11), .Q(p_unit_i_0_int_ps0_1_) );
  DFFR_X1 p_unit_i_0_int_ps0_reg_2_ ( .D(p_unit_i_0_n12), .CK(
        p_unit_i_0_net3011), .RN(p_unit_i_0_n11), .Q(p_unit_i_0_int_ps0_2_), 
        .QN(p_unit_i_0_n5) );
  CLKGATETST_X1 p_unit_i_0_clk_gate_o_data_reg_latch ( .CK(ck), .E(
        ps_ctrl_en_p), .SE(1'b0), .GCK(p_unit_i_0_net3011) );
  INV_X1 p_unit_i_1_U18 ( .A(n48), .ZN(p_unit_i_1_n11) );
  INV_X1 p_unit_i_1_U17 ( .A(p_unit_i_1_n8), .ZN(p_unit_i_1_n16) );
  NOR2_X1 p_unit_i_1_U15 ( .A1(p_unit_i_1_int_ps0_2_), .A2(p_unit_i_1_n16), 
        .ZN(p_unit_i_1_n6) );
  OAI22_X1 p_unit_i_1_U14 ( .A1(p_unit_i_1_n8), .A2(p_unit_i_1_n5), .B1(
        p_unit_i_1_n6), .B2(p_unit_i_1_n7), .ZN(p_unit_i_1_n4) );
  XNOR2_X1 p_unit_i_1_U13 ( .A(p_unit_i_1_n8), .B(p_unit_i_1_n9), .ZN(
        p_unit_i_1_N7) );
  XNOR2_X1 p_unit_i_1_U12 ( .A(p_unit_i_1_int_ps1_1_), .B(
        p_unit_i_1_int_ps0_1_), .ZN(p_unit_i_1_n3) );
  NAND2_X1 p_unit_i_1_U11 ( .A1(p_unit_i_1_int_ps0_0_), .A2(
        p_unit_i_1_int_ps1_0_), .ZN(p_unit_i_1_n2) );
  XOR2_X1 p_unit_i_1_U10 ( .A(p_unit_i_1_n2), .B(p_unit_i_1_n3), .Z(
        p_unit_i_1_N6) );
  OAI211_X1 p_unit_i_1_U9 ( .C1(p_unit_i_1_int_ps0_1_), .C2(
        p_unit_i_1_int_ps1_1_), .A(p_unit_i_1_int_ps0_0_), .B(
        p_unit_i_1_int_ps1_0_), .ZN(p_unit_i_1_n10) );
  INV_X1 p_unit_i_1_U8 ( .A(p_unit_i_1_n10), .ZN(p_unit_i_1_n17) );
  AOI21_X1 p_unit_i_1_U7 ( .B1(p_unit_i_1_int_ps0_1_), .B2(
        p_unit_i_1_int_ps1_1_), .A(p_unit_i_1_n17), .ZN(p_unit_i_1_n8) );
  AND3_X1 p_unit_i_1_U6 ( .A1(o_data_relu[10]), .A2(p_unit_i_1_n15), .A3(
        o_data_relu[8]), .ZN(p_unit_i_1_n14) );
  AOI21_X1 p_unit_i_1_U5 ( .B1(o_data_relu[9]), .B2(o_data_relu[11]), .A(
        p_unit_i_1_n14), .ZN(p_unit_i_1_n13) );
  INV_X1 p_unit_i_1_U4 ( .A(p_unit_i_1_n13), .ZN(p_unit_i_1_n12) );
  NAND2_X1 p_unit_i_1_U3 ( .A1(o_data_relu[10]), .A2(o_data_relu[8]), .ZN(
        p_unit_i_1_n1) );
  XNOR2_X1 p_unit_i_1_U2 ( .A(p_unit_i_1_n1), .B(p_unit_i_1_n15), .ZN(
        p_unit_i_1_N3) );
  XOR2_X1 p_unit_i_1_U22 ( .A(o_data_relu[8]), .B(o_data_relu[10]), .Z(
        p_unit_i_1_N2) );
  XOR2_X1 p_unit_i_1_U21 ( .A(o_data_relu[11]), .B(o_data_relu[9]), .Z(
        p_unit_i_1_n15) );
  XOR2_X1 p_unit_i_1_U19 ( .A(p_unit_i_1_int_ps1_0_), .B(p_unit_i_1_int_ps0_0_), .Z(p_unit_i_1_N5) );
  XOR2_X1 p_unit_i_1_U16 ( .A(p_unit_i_1_int_ps1_2_), .B(p_unit_i_1_int_ps0_2_), .Z(p_unit_i_1_n9) );
  DFFR_X1 p_unit_i_1_o_data_reg_1_ ( .D(p_unit_i_1_N6), .CK(p_unit_i_1_net2993), .RN(p_unit_i_1_n11), .Q(int_o_data_p[9]) );
  DFFR_X1 p_unit_i_1_o_data_reg_2_ ( .D(p_unit_i_1_N7), .CK(p_unit_i_1_net2993), .RN(p_unit_i_1_n11), .Q(int_o_data_p[10]) );
  DFFR_X1 p_unit_i_1_o_data_reg_3_ ( .D(p_unit_i_1_n4), .CK(p_unit_i_1_net2993), .RN(p_unit_i_1_n11), .Q(int_o_data_p[11]) );
  DFFR_X1 p_unit_i_1_o_data_reg_0_ ( .D(p_unit_i_1_N5), .CK(p_unit_i_1_net2993), .RN(p_unit_i_1_n11), .Q(int_o_data_p[8]) );
  DFFR_X1 p_unit_i_1_int_ps1_reg_0_ ( .D(p_unit_i_1_int_ps0_0_), .CK(
        p_unit_i_1_net2993), .RN(p_unit_i_1_n11), .Q(p_unit_i_1_int_ps1_0_) );
  DFFR_X1 p_unit_i_1_int_ps1_reg_1_ ( .D(p_unit_i_1_int_ps0_1_), .CK(
        p_unit_i_1_net2993), .RN(p_unit_i_1_n11), .Q(p_unit_i_1_int_ps1_1_) );
  DFFR_X1 p_unit_i_1_int_ps1_reg_2_ ( .D(p_unit_i_1_int_ps0_2_), .CK(
        p_unit_i_1_net2993), .RN(p_unit_i_1_n11), .Q(p_unit_i_1_int_ps1_2_), 
        .QN(p_unit_i_1_n7) );
  DFFR_X1 p_unit_i_1_int_ps0_reg_0_ ( .D(p_unit_i_1_N2), .CK(
        p_unit_i_1_net2993), .RN(p_unit_i_1_n11), .Q(p_unit_i_1_int_ps0_0_) );
  DFFR_X1 p_unit_i_1_int_ps0_reg_1_ ( .D(p_unit_i_1_N3), .CK(
        p_unit_i_1_net2993), .RN(p_unit_i_1_n11), .Q(p_unit_i_1_int_ps0_1_) );
  DFFR_X1 p_unit_i_1_int_ps0_reg_2_ ( .D(p_unit_i_1_n12), .CK(
        p_unit_i_1_net2993), .RN(p_unit_i_1_n11), .Q(p_unit_i_1_int_ps0_2_), 
        .QN(p_unit_i_1_n5) );
  CLKGATETST_X1 p_unit_i_1_clk_gate_o_data_reg_latch ( .CK(ck), .E(
        ps_ctrl_en_p), .SE(1'b0), .GCK(p_unit_i_1_net2993) );
  INV_X1 p_unit_i_2_U18 ( .A(n48), .ZN(p_unit_i_2_n11) );
  INV_X1 p_unit_i_2_U17 ( .A(p_unit_i_2_n8), .ZN(p_unit_i_2_n16) );
  NOR2_X1 p_unit_i_2_U15 ( .A1(p_unit_i_2_int_ps0_2_), .A2(p_unit_i_2_n16), 
        .ZN(p_unit_i_2_n6) );
  OAI22_X1 p_unit_i_2_U14 ( .A1(p_unit_i_2_n8), .A2(p_unit_i_2_n5), .B1(
        p_unit_i_2_n6), .B2(p_unit_i_2_n7), .ZN(p_unit_i_2_n4) );
  XNOR2_X1 p_unit_i_2_U13 ( .A(p_unit_i_2_n8), .B(p_unit_i_2_n9), .ZN(
        p_unit_i_2_N7) );
  XNOR2_X1 p_unit_i_2_U12 ( .A(p_unit_i_2_int_ps1_1_), .B(
        p_unit_i_2_int_ps0_1_), .ZN(p_unit_i_2_n3) );
  NAND2_X1 p_unit_i_2_U11 ( .A1(p_unit_i_2_int_ps0_0_), .A2(
        p_unit_i_2_int_ps1_0_), .ZN(p_unit_i_2_n2) );
  XOR2_X1 p_unit_i_2_U10 ( .A(p_unit_i_2_n2), .B(p_unit_i_2_n3), .Z(
        p_unit_i_2_N6) );
  OAI211_X1 p_unit_i_2_U9 ( .C1(p_unit_i_2_int_ps0_1_), .C2(
        p_unit_i_2_int_ps1_1_), .A(p_unit_i_2_int_ps0_0_), .B(
        p_unit_i_2_int_ps1_0_), .ZN(p_unit_i_2_n10) );
  INV_X1 p_unit_i_2_U8 ( .A(p_unit_i_2_n10), .ZN(p_unit_i_2_n17) );
  AOI21_X1 p_unit_i_2_U7 ( .B1(p_unit_i_2_int_ps0_1_), .B2(
        p_unit_i_2_int_ps1_1_), .A(p_unit_i_2_n17), .ZN(p_unit_i_2_n8) );
  AND3_X1 p_unit_i_2_U6 ( .A1(o_data_relu[6]), .A2(p_unit_i_2_n15), .A3(
        o_data_relu[4]), .ZN(p_unit_i_2_n14) );
  AOI21_X1 p_unit_i_2_U5 ( .B1(o_data_relu[5]), .B2(o_data_relu[7]), .A(
        p_unit_i_2_n14), .ZN(p_unit_i_2_n13) );
  INV_X1 p_unit_i_2_U4 ( .A(p_unit_i_2_n13), .ZN(p_unit_i_2_n12) );
  NAND2_X1 p_unit_i_2_U3 ( .A1(o_data_relu[6]), .A2(o_data_relu[4]), .ZN(
        p_unit_i_2_n1) );
  XNOR2_X1 p_unit_i_2_U2 ( .A(p_unit_i_2_n1), .B(p_unit_i_2_n15), .ZN(
        p_unit_i_2_N3) );
  XOR2_X1 p_unit_i_2_U22 ( .A(o_data_relu[4]), .B(o_data_relu[6]), .Z(
        p_unit_i_2_N2) );
  XOR2_X1 p_unit_i_2_U21 ( .A(o_data_relu[7]), .B(o_data_relu[5]), .Z(
        p_unit_i_2_n15) );
  XOR2_X1 p_unit_i_2_U19 ( .A(p_unit_i_2_int_ps1_0_), .B(p_unit_i_2_int_ps0_0_), .Z(p_unit_i_2_N5) );
  XOR2_X1 p_unit_i_2_U16 ( .A(p_unit_i_2_int_ps1_2_), .B(p_unit_i_2_int_ps0_2_), .Z(p_unit_i_2_n9) );
  DFFR_X1 p_unit_i_2_o_data_reg_1_ ( .D(p_unit_i_2_N6), .CK(p_unit_i_2_net2975), .RN(p_unit_i_2_n11), .Q(int_o_data_p[5]) );
  DFFR_X1 p_unit_i_2_o_data_reg_2_ ( .D(p_unit_i_2_N7), .CK(p_unit_i_2_net2975), .RN(p_unit_i_2_n11), .Q(int_o_data_p[6]) );
  DFFR_X1 p_unit_i_2_o_data_reg_3_ ( .D(p_unit_i_2_n4), .CK(p_unit_i_2_net2975), .RN(p_unit_i_2_n11), .Q(int_o_data_p[7]) );
  DFFR_X1 p_unit_i_2_o_data_reg_0_ ( .D(p_unit_i_2_N5), .CK(p_unit_i_2_net2975), .RN(p_unit_i_2_n11), .Q(int_o_data_p[4]) );
  DFFR_X1 p_unit_i_2_int_ps1_reg_0_ ( .D(p_unit_i_2_int_ps0_0_), .CK(
        p_unit_i_2_net2975), .RN(p_unit_i_2_n11), .Q(p_unit_i_2_int_ps1_0_) );
  DFFR_X1 p_unit_i_2_int_ps1_reg_1_ ( .D(p_unit_i_2_int_ps0_1_), .CK(
        p_unit_i_2_net2975), .RN(p_unit_i_2_n11), .Q(p_unit_i_2_int_ps1_1_) );
  DFFR_X1 p_unit_i_2_int_ps1_reg_2_ ( .D(p_unit_i_2_int_ps0_2_), .CK(
        p_unit_i_2_net2975), .RN(p_unit_i_2_n11), .Q(p_unit_i_2_int_ps1_2_), 
        .QN(p_unit_i_2_n7) );
  DFFR_X1 p_unit_i_2_int_ps0_reg_0_ ( .D(p_unit_i_2_N2), .CK(
        p_unit_i_2_net2975), .RN(p_unit_i_2_n11), .Q(p_unit_i_2_int_ps0_0_) );
  DFFR_X1 p_unit_i_2_int_ps0_reg_1_ ( .D(p_unit_i_2_N3), .CK(
        p_unit_i_2_net2975), .RN(p_unit_i_2_n11), .Q(p_unit_i_2_int_ps0_1_) );
  DFFR_X1 p_unit_i_2_int_ps0_reg_2_ ( .D(p_unit_i_2_n12), .CK(
        p_unit_i_2_net2975), .RN(p_unit_i_2_n11), .Q(p_unit_i_2_int_ps0_2_), 
        .QN(p_unit_i_2_n5) );
  CLKGATETST_X1 p_unit_i_2_clk_gate_o_data_reg_latch ( .CK(ck), .E(
        ps_ctrl_en_p), .SE(1'b0), .GCK(p_unit_i_2_net2975) );
  INV_X1 p_unit_i_3_U18 ( .A(n48), .ZN(p_unit_i_3_n11) );
  INV_X1 p_unit_i_3_U17 ( .A(p_unit_i_3_n8), .ZN(p_unit_i_3_n16) );
  NOR2_X1 p_unit_i_3_U15 ( .A1(p_unit_i_3_int_ps0_2_), .A2(p_unit_i_3_n16), 
        .ZN(p_unit_i_3_n6) );
  OAI22_X1 p_unit_i_3_U14 ( .A1(p_unit_i_3_n8), .A2(p_unit_i_3_n5), .B1(
        p_unit_i_3_n6), .B2(p_unit_i_3_n7), .ZN(p_unit_i_3_n4) );
  XNOR2_X1 p_unit_i_3_U13 ( .A(p_unit_i_3_n8), .B(p_unit_i_3_n9), .ZN(
        p_unit_i_3_N7) );
  XNOR2_X1 p_unit_i_3_U12 ( .A(p_unit_i_3_int_ps1_1_), .B(
        p_unit_i_3_int_ps0_1_), .ZN(p_unit_i_3_n3) );
  NAND2_X1 p_unit_i_3_U11 ( .A1(p_unit_i_3_int_ps0_0_), .A2(
        p_unit_i_3_int_ps1_0_), .ZN(p_unit_i_3_n2) );
  XOR2_X1 p_unit_i_3_U10 ( .A(p_unit_i_3_n2), .B(p_unit_i_3_n3), .Z(
        p_unit_i_3_N6) );
  OAI211_X1 p_unit_i_3_U9 ( .C1(p_unit_i_3_int_ps0_1_), .C2(
        p_unit_i_3_int_ps1_1_), .A(p_unit_i_3_int_ps0_0_), .B(
        p_unit_i_3_int_ps1_0_), .ZN(p_unit_i_3_n10) );
  INV_X1 p_unit_i_3_U8 ( .A(p_unit_i_3_n10), .ZN(p_unit_i_3_n17) );
  AOI21_X1 p_unit_i_3_U7 ( .B1(p_unit_i_3_int_ps0_1_), .B2(
        p_unit_i_3_int_ps1_1_), .A(p_unit_i_3_n17), .ZN(p_unit_i_3_n8) );
  AND3_X1 p_unit_i_3_U6 ( .A1(o_data_relu[2]), .A2(p_unit_i_3_n15), .A3(
        o_data_relu[0]), .ZN(p_unit_i_3_n14) );
  AOI21_X1 p_unit_i_3_U5 ( .B1(o_data_relu[1]), .B2(o_data_relu[3]), .A(
        p_unit_i_3_n14), .ZN(p_unit_i_3_n13) );
  INV_X1 p_unit_i_3_U4 ( .A(p_unit_i_3_n13), .ZN(p_unit_i_3_n12) );
  NAND2_X1 p_unit_i_3_U3 ( .A1(o_data_relu[2]), .A2(o_data_relu[0]), .ZN(
        p_unit_i_3_n1) );
  XNOR2_X1 p_unit_i_3_U2 ( .A(p_unit_i_3_n1), .B(p_unit_i_3_n15), .ZN(
        p_unit_i_3_N3) );
  XOR2_X1 p_unit_i_3_U22 ( .A(o_data_relu[0]), .B(o_data_relu[2]), .Z(
        p_unit_i_3_N2) );
  XOR2_X1 p_unit_i_3_U21 ( .A(o_data_relu[3]), .B(o_data_relu[1]), .Z(
        p_unit_i_3_n15) );
  XOR2_X1 p_unit_i_3_U19 ( .A(p_unit_i_3_int_ps1_0_), .B(p_unit_i_3_int_ps0_0_), .Z(p_unit_i_3_N5) );
  XOR2_X1 p_unit_i_3_U16 ( .A(p_unit_i_3_int_ps1_2_), .B(p_unit_i_3_int_ps0_2_), .Z(p_unit_i_3_n9) );
  DFFR_X1 p_unit_i_3_o_data_reg_1_ ( .D(p_unit_i_3_N6), .CK(p_unit_i_3_net2957), .RN(p_unit_i_3_n11), .Q(int_o_data_p[1]) );
  DFFR_X1 p_unit_i_3_o_data_reg_2_ ( .D(p_unit_i_3_N7), .CK(p_unit_i_3_net2957), .RN(p_unit_i_3_n11), .Q(int_o_data_p[2]) );
  DFFR_X1 p_unit_i_3_o_data_reg_3_ ( .D(p_unit_i_3_n4), .CK(p_unit_i_3_net2957), .RN(p_unit_i_3_n11), .Q(int_o_data_p[3]) );
  DFFR_X1 p_unit_i_3_o_data_reg_0_ ( .D(p_unit_i_3_N5), .CK(p_unit_i_3_net2957), .RN(p_unit_i_3_n11), .Q(int_o_data_p[0]) );
  DFFR_X1 p_unit_i_3_int_ps1_reg_0_ ( .D(p_unit_i_3_int_ps0_0_), .CK(
        p_unit_i_3_net2957), .RN(p_unit_i_3_n11), .Q(p_unit_i_3_int_ps1_0_) );
  DFFR_X1 p_unit_i_3_int_ps1_reg_1_ ( .D(p_unit_i_3_int_ps0_1_), .CK(
        p_unit_i_3_net2957), .RN(p_unit_i_3_n11), .Q(p_unit_i_3_int_ps1_1_) );
  DFFR_X1 p_unit_i_3_int_ps1_reg_2_ ( .D(p_unit_i_3_int_ps0_2_), .CK(
        p_unit_i_3_net2957), .RN(p_unit_i_3_n11), .Q(p_unit_i_3_int_ps1_2_), 
        .QN(p_unit_i_3_n7) );
  DFFR_X1 p_unit_i_3_int_ps0_reg_0_ ( .D(p_unit_i_3_N2), .CK(
        p_unit_i_3_net2957), .RN(p_unit_i_3_n11), .Q(p_unit_i_3_int_ps0_0_) );
  DFFR_X1 p_unit_i_3_int_ps0_reg_1_ ( .D(p_unit_i_3_N3), .CK(
        p_unit_i_3_net2957), .RN(p_unit_i_3_n11), .Q(p_unit_i_3_int_ps0_1_) );
  DFFR_X1 p_unit_i_3_int_ps0_reg_2_ ( .D(p_unit_i_3_n12), .CK(
        p_unit_i_3_net2957), .RN(p_unit_i_3_n11), .Q(p_unit_i_3_int_ps0_2_), 
        .QN(p_unit_i_3_n5) );
  CLKGATETST_X1 p_unit_i_3_clk_gate_o_data_reg_latch ( .CK(ck), .E(
        ps_ctrl_en_p), .SE(1'b0), .GCK(p_unit_i_3_net2957) );
  INV_X1 round_i_0_U5 ( .A(int_o_data_p[14]), .ZN(round_i_0_n2) );
  OAI21_X1 round_i_0_U4 ( .B1(int_o_data_p[13]), .B2(round_i_0_n2), .A(
        round_i_0_n3), .ZN(o_data[6]) );
  NAND2_X1 round_i_0_U3 ( .A1(int_o_data_p[13]), .A2(int_o_data_p[14]), .ZN(
        round_i_0_n1) );
  XNOR2_X1 round_i_0_U2 ( .A(int_o_data_p[15]), .B(round_i_0_n1), .ZN(
        o_data[7]) );
  NAND3_X1 round_i_0_U6 ( .A1(int_o_data_p[13]), .A2(round_i_0_n2), .A3(
        int_o_data_p[12]), .ZN(round_i_0_n3) );
  INV_X1 round_i_1_U5 ( .A(int_o_data_p[10]), .ZN(round_i_1_n2) );
  OAI21_X1 round_i_1_U4 ( .B1(int_o_data_p[9]), .B2(round_i_1_n2), .A(
        round_i_1_n4), .ZN(o_data[4]) );
  NAND2_X1 round_i_1_U3 ( .A1(int_o_data_p[9]), .A2(int_o_data_p[10]), .ZN(
        round_i_1_n1) );
  XNOR2_X1 round_i_1_U2 ( .A(int_o_data_p[11]), .B(round_i_1_n1), .ZN(
        o_data[5]) );
  NAND3_X1 round_i_1_U6 ( .A1(int_o_data_p[9]), .A2(round_i_1_n2), .A3(
        int_o_data_p[8]), .ZN(round_i_1_n4) );
  INV_X1 round_i_2_U5 ( .A(int_o_data_p[6]), .ZN(round_i_2_n2) );
  OAI21_X1 round_i_2_U4 ( .B1(int_o_data_p[5]), .B2(round_i_2_n2), .A(
        round_i_2_n4), .ZN(o_data[2]) );
  NAND2_X1 round_i_2_U3 ( .A1(int_o_data_p[5]), .A2(int_o_data_p[6]), .ZN(
        round_i_2_n1) );
  XNOR2_X1 round_i_2_U2 ( .A(int_o_data_p[7]), .B(round_i_2_n1), .ZN(o_data[3]) );
  NAND3_X1 round_i_2_U6 ( .A1(int_o_data_p[5]), .A2(round_i_2_n2), .A3(
        int_o_data_p[4]), .ZN(round_i_2_n4) );
  INV_X1 round_i_3_U5 ( .A(int_o_data_p[2]), .ZN(round_i_3_n2) );
  OAI21_X1 round_i_3_U4 ( .B1(int_o_data_p[1]), .B2(round_i_3_n2), .A(
        round_i_3_n4), .ZN(o_data[0]) );
  NAND2_X1 round_i_3_U3 ( .A1(int_o_data_p[1]), .A2(int_o_data_p[2]), .ZN(
        round_i_3_n1) );
  XNOR2_X1 round_i_3_U2 ( .A(int_o_data_p[3]), .B(round_i_3_n1), .ZN(o_data[1]) );
  NAND3_X1 round_i_3_U6 ( .A1(int_o_data_p[1]), .A2(round_i_3_n2), .A3(
        int_o_data_p[0]), .ZN(round_i_3_n4) );
  INV_X1 hmode_cnt_inst_U14 ( .A(n48), .ZN(hmode_cnt_inst_n12) );
  AOI21_X1 hmode_cnt_inst_U13 ( .B1(hmode_cnt_inst_n10), .B2(hmode_cnt_inst_n7), .A(hmode_cnt_inst_N10), .ZN(hmode_cnt_inst_n8) );
  NAND4_X1 hmode_cnt_inst_U12 ( .A1(hmode_cnt_inst_n10), .A2(int_hmode_cnt[1]), 
        .A3(int_hmode_cnt[0]), .A4(hmode_cnt_inst_n5), .ZN(hmode_cnt_inst_n9)
         );
  OAI21_X1 hmode_cnt_inst_U11 ( .B1(hmode_cnt_inst_n8), .B2(hmode_cnt_inst_n5), 
        .A(hmode_cnt_inst_n9), .ZN(hmode_cnt_inst_N12) );
  XNOR2_X1 hmode_cnt_inst_U10 ( .A(int_hmode_cnt[0]), .B(int_hmode_cnt[1]), 
        .ZN(hmode_cnt_inst_n11) );
  AND2_X1 hmode_cnt_inst_U9 ( .A1(hmode_cnt_inst_n10), .A2(hmode_cnt_inst_n6), 
        .ZN(hmode_cnt_inst_N10) );
  NOR2_X1 hmode_cnt_inst_U8 ( .A1(s_tc_hmode), .A2(1'b0), .ZN(
        hmode_cnt_inst_n10) );
  XOR2_X1 hmode_cnt_inst_U7 ( .A(int_hmode_cnt[1]), .B(arv_k[1]), .Z(
        hmode_cnt_inst_n4) );
  XOR2_X1 hmode_cnt_inst_U6 ( .A(int_hmode_cnt[0]), .B(arv_k[0]), .Z(
        hmode_cnt_inst_n2) );
  XOR2_X1 hmode_cnt_inst_U5 ( .A(int_hmode_cnt[2]), .B(arv_k[2]), .Z(
        hmode_cnt_inst_n1) );
  NOR3_X1 hmode_cnt_inst_U4 ( .A1(hmode_cnt_inst_n1), .A2(hmode_cnt_inst_n2), 
        .A3(hmode_cnt_inst_n4), .ZN(s_tc_hmode) );
  DFFR_X1 hmode_cnt_inst_cnt_out_reg_2_ ( .D(hmode_cnt_inst_N12), .CK(
        hmode_cnt_inst_net2939), .RN(hmode_cnt_inst_n12), .Q(int_hmode_cnt[2]), 
        .QN(hmode_cnt_inst_n5) );
  SDFFR_X1 hmode_cnt_inst_cnt_out_reg_1_ ( .D(hmode_cnt_inst_n10), .SI(1'b0), 
        .SE(hmode_cnt_inst_n11), .CK(hmode_cnt_inst_net2939), .RN(
        hmode_cnt_inst_n12), .Q(int_hmode_cnt[1]), .QN(hmode_cnt_inst_n7) );
  DFFR_X1 hmode_cnt_inst_cnt_out_reg_0_ ( .D(hmode_cnt_inst_N10), .CK(
        hmode_cnt_inst_net2939), .RN(hmode_cnt_inst_n12), .Q(int_hmode_cnt[0]), 
        .QN(hmode_cnt_inst_n6) );
  CLKGATETST_X1 hmode_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        int_en_hmode), .SE(1'b0), .GCK(hmode_cnt_inst_net2939) );
  INV_X1 vmode_cnt_inst_U14 ( .A(n47), .ZN(vmode_cnt_inst_n12) );
  AOI21_X1 vmode_cnt_inst_U13 ( .B1(vmode_cnt_inst_n10), .B2(vmode_cnt_inst_n7), .A(vmode_cnt_inst_N10), .ZN(vmode_cnt_inst_n8) );
  NAND4_X1 vmode_cnt_inst_U12 ( .A1(vmode_cnt_inst_n10), .A2(
        vmode_cnt_inst_q_1_), .A3(vmode_cnt_inst_q_0_), .A4(vmode_cnt_inst_n5), 
        .ZN(vmode_cnt_inst_n9) );
  OAI21_X1 vmode_cnt_inst_U11 ( .B1(vmode_cnt_inst_n8), .B2(vmode_cnt_inst_n5), 
        .A(vmode_cnt_inst_n9), .ZN(vmode_cnt_inst_N12) );
  XNOR2_X1 vmode_cnt_inst_U10 ( .A(vmode_cnt_inst_q_0_), .B(
        vmode_cnt_inst_q_1_), .ZN(vmode_cnt_inst_n11) );
  AND2_X1 vmode_cnt_inst_U9 ( .A1(vmode_cnt_inst_n10), .A2(vmode_cnt_inst_n6), 
        .ZN(vmode_cnt_inst_N10) );
  NOR2_X1 vmode_cnt_inst_U8 ( .A1(s_tc_vmode), .A2(1'b0), .ZN(
        vmode_cnt_inst_n10) );
  XOR2_X1 vmode_cnt_inst_U7 ( .A(vmode_cnt_inst_q_1_), .B(arv_k[1]), .Z(
        vmode_cnt_inst_n4) );
  XOR2_X1 vmode_cnt_inst_U6 ( .A(vmode_cnt_inst_q_0_), .B(arv_k[0]), .Z(
        vmode_cnt_inst_n2) );
  XOR2_X1 vmode_cnt_inst_U5 ( .A(vmode_cnt_inst_q_2_), .B(arv_k[2]), .Z(
        vmode_cnt_inst_n1) );
  NOR3_X1 vmode_cnt_inst_U4 ( .A1(vmode_cnt_inst_n1), .A2(vmode_cnt_inst_n2), 
        .A3(vmode_cnt_inst_n4), .ZN(s_tc_vmode) );
  DFFR_X1 vmode_cnt_inst_cnt_out_reg_2_ ( .D(vmode_cnt_inst_N12), .CK(
        vmode_cnt_inst_net2921), .RN(vmode_cnt_inst_n12), .Q(
        vmode_cnt_inst_q_2_), .QN(vmode_cnt_inst_n5) );
  SDFFR_X1 vmode_cnt_inst_cnt_out_reg_1_ ( .D(vmode_cnt_inst_n10), .SI(1'b0), 
        .SE(vmode_cnt_inst_n11), .CK(vmode_cnt_inst_net2921), .RN(
        vmode_cnt_inst_n12), .Q(vmode_cnt_inst_q_1_), .QN(vmode_cnt_inst_n7)
         );
  DFFR_X1 vmode_cnt_inst_cnt_out_reg_0_ ( .D(vmode_cnt_inst_N10), .CK(
        vmode_cnt_inst_net2921), .RN(vmode_cnt_inst_n12), .Q(
        vmode_cnt_inst_q_0_), .QN(vmode_cnt_inst_n6) );
  CLKGATETST_X1 vmode_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        int_en_vmode), .SE(1'b0), .GCK(vmode_cnt_inst_net2921) );
  INV_X1 res_cnt_inst_U14 ( .A(n47), .ZN(res_cnt_inst_n2) );
  XNOR2_X1 res_cnt_inst_U13 ( .A(res_cnt_inst_q_0_), .B(res_cnt_inst_q_1_), 
        .ZN(res_cnt_inst_n11) );
  AND2_X1 res_cnt_inst_U12 ( .A1(res_cnt_inst_n10), .A2(res_cnt_inst_n1), .ZN(
        res_cnt_inst_N10) );
  AOI21_X1 res_cnt_inst_U11 ( .B1(res_cnt_inst_n10), .B2(res_cnt_inst_n7), .A(
        res_cnt_inst_N10), .ZN(res_cnt_inst_n8) );
  NAND4_X1 res_cnt_inst_U10 ( .A1(res_cnt_inst_n10), .A2(res_cnt_inst_q_1_), 
        .A3(res_cnt_inst_q_0_), .A4(res_cnt_inst_n5), .ZN(res_cnt_inst_n9) );
  OAI21_X1 res_cnt_inst_U9 ( .B1(res_cnt_inst_n8), .B2(res_cnt_inst_n5), .A(
        res_cnt_inst_n9), .ZN(res_cnt_inst_N12) );
  XNOR2_X1 res_cnt_inst_U8 ( .A(res_cnt_inst_q_1_), .B(int_arv_res[1]), .ZN(
        res_cnt_inst_n14) );
  XNOR2_X1 res_cnt_inst_U7 ( .A(res_cnt_inst_q_0_), .B(int_arv_res[0]), .ZN(
        res_cnt_inst_n13) );
  XNOR2_X1 res_cnt_inst_U6 ( .A(res_cnt_inst_q_2_), .B(int_arv_res[2]), .ZN(
        res_cnt_inst_n12) );
  AND3_X1 res_cnt_inst_U5 ( .A1(res_cnt_inst_n12), .A2(res_cnt_inst_n13), .A3(
        res_cnt_inst_n14), .ZN(s_tc_res) );
  NOR2_X1 res_cnt_inst_U4 ( .A1(s_tc_res), .A2(1'b0), .ZN(res_cnt_inst_n10) );
  DFFR_X1 res_cnt_inst_cnt_out_reg_2_ ( .D(res_cnt_inst_N12), .CK(
        res_cnt_inst_net2903), .RN(res_cnt_inst_n2), .Q(res_cnt_inst_q_2_), 
        .QN(res_cnt_inst_n5) );
  SDFFR_X1 res_cnt_inst_cnt_out_reg_1_ ( .D(res_cnt_inst_n10), .SI(1'b0), .SE(
        res_cnt_inst_n11), .CK(res_cnt_inst_net2903), .RN(res_cnt_inst_n2), 
        .Q(res_cnt_inst_q_1_), .QN(res_cnt_inst_n7) );
  DFFR_X1 res_cnt_inst_cnt_out_reg_0_ ( .D(res_cnt_inst_N10), .CK(
        res_cnt_inst_net2903), .RN(res_cnt_inst_n2), .Q(res_cnt_inst_q_0_), 
        .QN(res_cnt_inst_n1) );
  CLKGATETST_X1 res_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        ctrl_wr_pipe), .SE(1'b0), .GCK(res_cnt_inst_net2903) );
  INV_X1 i_data_npu_cnt_inst_U14 ( .A(n47), .ZN(i_data_npu_cnt_inst_n12) );
  AOI21_X1 i_data_npu_cnt_inst_U13 ( .B1(i_data_npu_cnt_inst_n10), .B2(
        i_data_npu_cnt_inst_n7), .A(i_data_npu_cnt_inst_N10), .ZN(
        i_data_npu_cnt_inst_n8) );
  NAND4_X1 i_data_npu_cnt_inst_U12 ( .A1(i_data_npu_cnt_inst_n10), .A2(
        int_npu_ptr[1]), .A3(int_npu_ptr[0]), .A4(i_data_npu_cnt_inst_n5), 
        .ZN(i_data_npu_cnt_inst_n9) );
  OAI21_X1 i_data_npu_cnt_inst_U11 ( .B1(i_data_npu_cnt_inst_n8), .B2(
        i_data_npu_cnt_inst_n5), .A(i_data_npu_cnt_inst_n9), .ZN(
        i_data_npu_cnt_inst_N12) );
  XOR2_X1 i_data_npu_cnt_inst_U10 ( .A(int_npu_ptr[1]), .B(1'b1), .Z(
        i_data_npu_cnt_inst_n6) );
  XOR2_X1 i_data_npu_cnt_inst_U9 ( .A(int_npu_ptr[0]), .B(1'b1), .Z(
        i_data_npu_cnt_inst_n4) );
  XOR2_X1 i_data_npu_cnt_inst_U8 ( .A(int_npu_ptr[2]), .B(1'b1), .Z(
        i_data_npu_cnt_inst_n2) );
  NOR3_X1 i_data_npu_cnt_inst_U7 ( .A1(i_data_npu_cnt_inst_n2), .A2(
        i_data_npu_cnt_inst_n4), .A3(i_data_npu_cnt_inst_n6), .ZN(s_tc_npu_ptr) );
  XNOR2_X1 i_data_npu_cnt_inst_U6 ( .A(int_npu_ptr[0]), .B(int_npu_ptr[1]), 
        .ZN(i_data_npu_cnt_inst_n11) );
  AND2_X1 i_data_npu_cnt_inst_U5 ( .A1(i_data_npu_cnt_inst_n10), .A2(
        i_data_npu_cnt_inst_n1), .ZN(i_data_npu_cnt_inst_N10) );
  NOR2_X1 i_data_npu_cnt_inst_U4 ( .A1(s_tc_npu_ptr), .A2(1'b0), .ZN(
        i_data_npu_cnt_inst_n10) );
  DFFR_X1 i_data_npu_cnt_inst_cnt_out_reg_2_ ( .D(i_data_npu_cnt_inst_N12), 
        .CK(i_data_npu_cnt_inst_net2885), .RN(i_data_npu_cnt_inst_n12), .Q(
        int_npu_ptr[2]), .QN(i_data_npu_cnt_inst_n5) );
  SDFFR_X1 i_data_npu_cnt_inst_cnt_out_reg_1_ ( .D(i_data_npu_cnt_inst_n10), 
        .SI(1'b0), .SE(i_data_npu_cnt_inst_n11), .CK(
        i_data_npu_cnt_inst_net2885), .RN(i_data_npu_cnt_inst_n12), .Q(
        int_npu_ptr[1]), .QN(i_data_npu_cnt_inst_n7) );
  DFFR_X1 i_data_npu_cnt_inst_cnt_out_reg_0_ ( .D(i_data_npu_cnt_inst_N10), 
        .CK(i_data_npu_cnt_inst_net2885), .RN(i_data_npu_cnt_inst_n12), .Q(
        int_npu_ptr[0]), .QN(i_data_npu_cnt_inst_n1) );
  CLKGATETST_X1 i_data_npu_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        int_en_npu_ptr), .SE(1'b0), .GCK(i_data_npu_cnt_inst_net2885) );
  INV_X1 i_data_tilev_cnt_inst_U16 ( .A(n47), .ZN(i_data_tilev_cnt_inst_n3) );
  INV_X1 i_data_tilev_cnt_inst_U15 ( .A(arv_i_tile[0]), .ZN(
        i_data_tilev_cnt_inst_n8) );
  NOR2_X1 i_data_tilev_cnt_inst_U14 ( .A1(1'b0), .A2(
        i_data_tilev_cnt_inst_q_0_), .ZN(i_data_tilev_cnt_inst_n13) );
  OAI211_X1 i_data_tilev_cnt_inst_U13 ( .C1(arv_i_tile[0]), .C2(
        i_data_tilev_cnt_inst_n12), .A(int_en_tilev_ptr), .B(
        i_data_tilev_cnt_inst_n13), .ZN(i_data_tilev_cnt_inst_n11) );
  OAI21_X1 i_data_tilev_cnt_inst_U12 ( .B1(int_en_tilev_ptr), .B2(
        i_data_tilev_cnt_inst_n2), .A(i_data_tilev_cnt_inst_n11), .ZN(
        i_data_tilev_cnt_inst_n17) );
  OAI21_X1 i_data_tilev_cnt_inst_U11 ( .B1(i_data_tilev_cnt_inst_n8), .B2(
        arv_i_tile[1]), .A(i_data_tilev_cnt_inst_n1), .ZN(
        i_data_tilev_cnt_inst_n9) );
  AND2_X1 i_data_tilev_cnt_inst_U10 ( .A1(int_en_tilev_ptr), .A2(
        i_data_tilev_cnt_inst_q_0_), .ZN(i_data_tilev_cnt_inst_n5) );
  XNOR2_X1 i_data_tilev_cnt_inst_U9 ( .A(i_data_tilev_cnt_inst_n2), .B(
        arv_i_tile[0]), .ZN(i_data_tilev_cnt_inst_n14) );
  NOR2_X1 i_data_tilev_cnt_inst_U8 ( .A1(i_data_tilev_cnt_inst_n12), .A2(
        i_data_tilev_cnt_inst_n14), .ZN(int_d_tc[2]) );
  INV_X1 i_data_tilev_cnt_inst_U7 ( .A(i_data_tilev_cnt_inst_n9), .ZN(
        i_data_tilev_cnt_inst_n6) );
  AOI21_X1 i_data_tilev_cnt_inst_U6 ( .B1(arv_i_tile[1]), .B2(
        i_data_tilev_cnt_inst_n8), .A(i_data_tilev_cnt_inst_q_0_), .ZN(
        i_data_tilev_cnt_inst_n7) );
  AOI22_X1 i_data_tilev_cnt_inst_U5 ( .A1(i_data_tilev_cnt_inst_n5), .A2(
        i_data_tilev_cnt_inst_n6), .B1(i_data_tilev_cnt_inst_n7), .B2(
        i_data_tilev_cnt_inst_q_1_), .ZN(i_data_tilev_cnt_inst_n4) );
  OAI22_X1 i_data_tilev_cnt_inst_U4 ( .A1(int_en_tilev_ptr), .A2(
        i_data_tilev_cnt_inst_n1), .B1(1'b0), .B2(i_data_tilev_cnt_inst_n4), 
        .ZN(i_data_tilev_cnt_inst_n15) );
  XNOR2_X1 i_data_tilev_cnt_inst_U3 ( .A(arv_i_tile[1]), .B(
        i_data_tilev_cnt_inst_n1), .ZN(i_data_tilev_cnt_inst_n12) );
  DFFR_X1 i_data_tilev_cnt_inst_cnt_out_reg_1_ ( .D(i_data_tilev_cnt_inst_n15), 
        .CK(ck), .RN(i_data_tilev_cnt_inst_n3), .Q(i_data_tilev_cnt_inst_q_1_), 
        .QN(i_data_tilev_cnt_inst_n1) );
  DFFR_X1 i_data_tilev_cnt_inst_cnt_out_reg_0_ ( .D(i_data_tilev_cnt_inst_n17), 
        .CK(ck), .RN(i_data_tilev_cnt_inst_n3), .Q(i_data_tilev_cnt_inst_q_0_), 
        .QN(i_data_tilev_cnt_inst_n2) );
  INV_X1 i_data_tileh_cnt_inst_U16 ( .A(n48), .ZN(i_data_tileh_cnt_inst_n1) );
  INV_X1 i_data_tileh_cnt_inst_U15 ( .A(arv_i_tile[0]), .ZN(
        i_data_tileh_cnt_inst_n8) );
  OAI21_X1 i_data_tileh_cnt_inst_U14 ( .B1(i_data_tileh_cnt_inst_n8), .B2(
        arv_i_tile[1]), .A(i_data_tileh_cnt_inst_n6), .ZN(
        i_data_tileh_cnt_inst_n21) );
  AND2_X1 i_data_tileh_cnt_inst_U13 ( .A1(n59), .A2(i_data_ev_odd_n), .ZN(
        i_data_tileh_cnt_inst_n23) );
  NOR2_X1 i_data_tileh_cnt_inst_U12 ( .A1(1'b0), .A2(i_data_ev_odd_n), .ZN(
        i_data_tileh_cnt_inst_n18) );
  OAI211_X1 i_data_tileh_cnt_inst_U11 ( .C1(arv_i_tile[0]), .C2(
        i_data_tileh_cnt_inst_n19), .A(n59), .B(i_data_tileh_cnt_inst_n18), 
        .ZN(i_data_tileh_cnt_inst_n20) );
  OAI21_X1 i_data_tileh_cnt_inst_U10 ( .B1(n59), .B2(i_data_tileh_cnt_inst_n2), 
        .A(i_data_tileh_cnt_inst_n20), .ZN(i_data_tileh_cnt_inst_n10) );
  XNOR2_X1 i_data_tileh_cnt_inst_U9 ( .A(i_data_tileh_cnt_inst_n2), .B(
        arv_i_tile[0]), .ZN(i_data_tileh_cnt_inst_n17) );
  NOR2_X1 i_data_tileh_cnt_inst_U8 ( .A1(i_data_tileh_cnt_inst_n19), .A2(
        i_data_tileh_cnt_inst_n17), .ZN(int_d_tc[1]) );
  INV_X1 i_data_tileh_cnt_inst_U7 ( .A(i_data_tileh_cnt_inst_n21), .ZN(
        i_data_tileh_cnt_inst_n3) );
  AOI21_X1 i_data_tileh_cnt_inst_U6 ( .B1(arv_i_tile[1]), .B2(
        i_data_tileh_cnt_inst_n8), .A(i_data_ev_odd_n), .ZN(
        i_data_tileh_cnt_inst_n22) );
  AOI22_X1 i_data_tileh_cnt_inst_U5 ( .A1(i_data_tileh_cnt_inst_n23), .A2(
        i_data_tileh_cnt_inst_n3), .B1(i_data_tileh_cnt_inst_n22), .B2(
        int_tileh_ptr_1_), .ZN(i_data_tileh_cnt_inst_n24) );
  OAI22_X1 i_data_tileh_cnt_inst_U4 ( .A1(n59), .A2(i_data_tileh_cnt_inst_n6), 
        .B1(1'b0), .B2(i_data_tileh_cnt_inst_n24), .ZN(
        i_data_tileh_cnt_inst_n16) );
  XNOR2_X1 i_data_tileh_cnt_inst_U3 ( .A(arv_i_tile[1]), .B(
        i_data_tileh_cnt_inst_n6), .ZN(i_data_tileh_cnt_inst_n19) );
  DFFR_X1 i_data_tileh_cnt_inst_cnt_out_reg_1_ ( .D(i_data_tileh_cnt_inst_n16), 
        .CK(ck), .RN(i_data_tileh_cnt_inst_n1), .Q(int_tileh_ptr_1_), .QN(
        i_data_tileh_cnt_inst_n6) );
  DFFR_X1 i_data_tileh_cnt_inst_cnt_out_reg_0_ ( .D(i_data_tileh_cnt_inst_n10), 
        .CK(ck), .RN(i_data_tileh_cnt_inst_n1), .Q(i_data_ev_odd_n), .QN(
        i_data_tileh_cnt_inst_n2) );
  INV_X1 ifmaps_cnt_inst_U14 ( .A(n46), .ZN(ifmaps_cnt_inst_n12) );
  AOI21_X1 ifmaps_cnt_inst_U13 ( .B1(ifmaps_cnt_inst_n10), .B2(
        ifmaps_cnt_inst_n7), .A(ifmaps_cnt_inst_N10), .ZN(ifmaps_cnt_inst_n8)
         );
  NAND4_X1 ifmaps_cnt_inst_U12 ( .A1(ifmaps_cnt_inst_n10), .A2(
        int_ifmaps_ptr[1]), .A3(int_ifmaps_ptr[0]), .A4(ifmaps_cnt_inst_n5), 
        .ZN(ifmaps_cnt_inst_n9) );
  OAI21_X1 ifmaps_cnt_inst_U11 ( .B1(ifmaps_cnt_inst_n8), .B2(
        ifmaps_cnt_inst_n5), .A(ifmaps_cnt_inst_n9), .ZN(ifmaps_cnt_inst_N12)
         );
  XNOR2_X1 ifmaps_cnt_inst_U10 ( .A(int_ifmaps_ptr[0]), .B(int_ifmaps_ptr[1]), 
        .ZN(ifmaps_cnt_inst_n11) );
  AND2_X1 ifmaps_cnt_inst_U9 ( .A1(ifmaps_cnt_inst_n10), .A2(
        ifmaps_cnt_inst_n6), .ZN(ifmaps_cnt_inst_N10) );
  NOR2_X1 ifmaps_cnt_inst_U8 ( .A1(s_tc_ifmaps), .A2(1'b0), .ZN(
        ifmaps_cnt_inst_n10) );
  XOR2_X1 ifmaps_cnt_inst_U7 ( .A(int_ifmaps_ptr[1]), .B(arv_ifmaps[1]), .Z(
        ifmaps_cnt_inst_n4) );
  XOR2_X1 ifmaps_cnt_inst_U6 ( .A(int_ifmaps_ptr[0]), .B(arv_ifmaps[0]), .Z(
        ifmaps_cnt_inst_n2) );
  XOR2_X1 ifmaps_cnt_inst_U5 ( .A(int_ifmaps_ptr[2]), .B(arv_ifmaps[2]), .Z(
        ifmaps_cnt_inst_n1) );
  NOR3_X1 ifmaps_cnt_inst_U4 ( .A1(ifmaps_cnt_inst_n1), .A2(ifmaps_cnt_inst_n2), .A3(ifmaps_cnt_inst_n4), .ZN(s_tc_ifmaps) );
  DFFR_X1 ifmaps_cnt_inst_cnt_out_reg_2_ ( .D(ifmaps_cnt_inst_N12), .CK(
        ifmaps_cnt_inst_net2867), .RN(ifmaps_cnt_inst_n12), .Q(
        int_ifmaps_ptr[2]), .QN(ifmaps_cnt_inst_n5) );
  SDFFR_X1 ifmaps_cnt_inst_cnt_out_reg_1_ ( .D(ifmaps_cnt_inst_n10), .SI(1'b0), 
        .SE(ifmaps_cnt_inst_n11), .CK(ifmaps_cnt_inst_net2867), .RN(
        ifmaps_cnt_inst_n12), .Q(int_ifmaps_ptr[1]), .QN(ifmaps_cnt_inst_n7)
         );
  DFFR_X1 ifmaps_cnt_inst_cnt_out_reg_0_ ( .D(ifmaps_cnt_inst_N10), .CK(
        ifmaps_cnt_inst_net2867), .RN(ifmaps_cnt_inst_n12), .Q(
        int_ifmaps_ptr[0]), .QN(ifmaps_cnt_inst_n6) );
  CLKGATETST_X1 ifmaps_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        ctrl_en_npu), .SE(1'b0), .GCK(ifmaps_cnt_inst_net2867) );
  INV_X1 ofmaps_cnt_inst_U17 ( .A(n47), .ZN(ofmaps_cnt_inst_n2) );
  XNOR2_X1 ofmaps_cnt_inst_U16 ( .A(ofmaps_cnt_inst_q_0_), .B(
        ofmaps_cnt_inst_q_1_), .ZN(ofmaps_cnt_inst_n15) );
  XNOR2_X1 ofmaps_cnt_inst_U15 ( .A(ofmaps_cnt_inst_q_3_), .B(arv_ofmaps[3]), 
        .ZN(ofmaps_cnt_inst_n18) );
  XNOR2_X1 ofmaps_cnt_inst_U14 ( .A(ofmaps_cnt_inst_q_2_), .B(arv_ofmaps[2]), 
        .ZN(ofmaps_cnt_inst_n17) );
  AND4_X1 ofmaps_cnt_inst_U13 ( .A1(ofmaps_cnt_inst_n16), .A2(
        ofmaps_cnt_inst_n17), .A3(ofmaps_cnt_inst_n18), .A4(
        ofmaps_cnt_inst_n19), .ZN(int_d_tc[0]) );
  INV_X1 ofmaps_cnt_inst_U12 ( .A(ofmaps_cnt_inst_n14), .ZN(ofmaps_cnt_inst_n4) );
  AOI21_X1 ofmaps_cnt_inst_U11 ( .B1(ofmaps_cnt_inst_n13), .B2(
        ofmaps_cnt_inst_n8), .A(ofmaps_cnt_inst_n4), .ZN(ofmaps_cnt_inst_n10)
         );
  OR3_X1 ofmaps_cnt_inst_U10 ( .A1(ofmaps_cnt_inst_n8), .A2(
        ofmaps_cnt_inst_q_3_), .A3(ofmaps_cnt_inst_n12), .ZN(
        ofmaps_cnt_inst_n11) );
  OAI21_X1 ofmaps_cnt_inst_U9 ( .B1(ofmaps_cnt_inst_n10), .B2(
        ofmaps_cnt_inst_n5), .A(ofmaps_cnt_inst_n11), .ZN(ofmaps_cnt_inst_N14)
         );
  AND2_X1 ofmaps_cnt_inst_U8 ( .A1(ofmaps_cnt_inst_n13), .A2(
        ofmaps_cnt_inst_n1), .ZN(ofmaps_cnt_inst_N11) );
  XNOR2_X1 ofmaps_cnt_inst_U7 ( .A(ofmaps_cnt_inst_q_0_), .B(arv_ofmaps[0]), 
        .ZN(ofmaps_cnt_inst_n19) );
  OAI22_X1 ofmaps_cnt_inst_U6 ( .A1(ofmaps_cnt_inst_n14), .A2(
        ofmaps_cnt_inst_n8), .B1(ofmaps_cnt_inst_q_2_), .B2(
        ofmaps_cnt_inst_n12), .ZN(ofmaps_cnt_inst_N13) );
  AOI21_X1 ofmaps_cnt_inst_U5 ( .B1(ofmaps_cnt_inst_n9), .B2(
        ofmaps_cnt_inst_n13), .A(ofmaps_cnt_inst_N11), .ZN(ofmaps_cnt_inst_n14) );
  NOR2_X1 ofmaps_cnt_inst_U4 ( .A1(int_d_tc[0]), .A2(1'b0), .ZN(
        ofmaps_cnt_inst_n13) );
  XOR2_X1 ofmaps_cnt_inst_U20 ( .A(ofmaps_cnt_inst_n9), .B(arv_ofmaps[1]), .Z(
        ofmaps_cnt_inst_n16) );
  NAND3_X1 ofmaps_cnt_inst_U19 ( .A1(ofmaps_cnt_inst_q_1_), .A2(
        ofmaps_cnt_inst_q_0_), .A3(ofmaps_cnt_inst_n13), .ZN(
        ofmaps_cnt_inst_n12) );
  DFFR_X1 ofmaps_cnt_inst_cnt_out_reg_3_ ( .D(ofmaps_cnt_inst_N14), .CK(
        ofmaps_cnt_inst_net2849), .RN(ofmaps_cnt_inst_n2), .Q(
        ofmaps_cnt_inst_q_3_), .QN(ofmaps_cnt_inst_n5) );
  DFFR_X1 ofmaps_cnt_inst_cnt_out_reg_2_ ( .D(ofmaps_cnt_inst_N13), .CK(
        ofmaps_cnt_inst_net2849), .RN(ofmaps_cnt_inst_n2), .Q(
        ofmaps_cnt_inst_q_2_), .QN(ofmaps_cnt_inst_n8) );
  SDFFR_X1 ofmaps_cnt_inst_cnt_out_reg_1_ ( .D(ofmaps_cnt_inst_n13), .SI(1'b0), 
        .SE(ofmaps_cnt_inst_n15), .CK(ofmaps_cnt_inst_net2849), .RN(
        ofmaps_cnt_inst_n2), .Q(ofmaps_cnt_inst_q_1_), .QN(ofmaps_cnt_inst_n9)
         );
  DFFR_X1 ofmaps_cnt_inst_cnt_out_reg_0_ ( .D(ofmaps_cnt_inst_N11), .CK(
        ofmaps_cnt_inst_net2849), .RN(ofmaps_cnt_inst_n2), .Q(
        ofmaps_cnt_inst_q_0_), .QN(ofmaps_cnt_inst_n1) );
  CLKGATETST_X1 ofmaps_cnt_inst_clk_gate_cnt_out_reg_latch ( .CK(ck), .E(
        int_en_ofmaps_ptr), .SE(1'b0), .GCK(ofmaps_cnt_inst_net2849) );
  CLKBUF_X1 i_weight_addr_gen_inst_U66 ( .A(i_weight_addr[15]), .Z(
        i_weight_addr_gen_inst_n8) );
  INV_X1 i_weight_addr_gen_inst_U65 ( .A(i_weight_addr_gen_inst_n6), .ZN(
        i_weight_addr_gen_inst_n7) );
  OR2_X1 i_weight_addr_gen_inst_U64 ( .A1(s_tc_res), .A2(ctrl_en_hmode), .ZN(
        i_weight_addr_gen_inst_N95) );
  OR2_X1 i_weight_addr_gen_inst_U63 ( .A1(int_c_i_en_weight_addr), .A2(1'b0), 
        .ZN(i_weight_addr_gen_inst_N58) );
  AOI22_X1 i_weight_addr_gen_inst_U62 ( .A1(i_weight_addr_gen_inst_N41), .A2(
        i_weight_addr_gen_inst_n45), .B1(i_weight_addr_gen_inst_N25), .B2(
        i_weight_addr_gen_inst_n46), .ZN(i_weight_addr_gen_inst_n44) );
  INV_X1 i_weight_addr_gen_inst_U61 ( .A(i_weight_addr_gen_inst_n44), .ZN(
        i_weight_addr_gen_inst_n29) );
  INV_X1 i_weight_addr_gen_inst_U60 ( .A(int_c_i_en_weight_addr), .ZN(
        i_weight_addr_gen_inst_n64) );
  INV_X1 i_weight_addr_gen_inst_U59 ( .A(s_tc_res), .ZN(
        i_weight_addr_gen_inst_n63) );
  AOI22_X1 i_weight_addr_gen_inst_U58 ( .A1(i_weight_addr_gen_inst_N26), .A2(
        i_weight_addr_gen_inst_n45), .B1(i_weight_addr_gen_inst_N10), .B2(
        i_weight_addr_gen_inst_n46), .ZN(i_weight_addr_gen_inst_n61) );
  INV_X1 i_weight_addr_gen_inst_U57 ( .A(i_weight_addr_gen_inst_n61), .ZN(
        i_weight_addr_gen_inst_n62) );
  AOI22_X1 i_weight_addr_gen_inst_U56 ( .A1(i_weight_addr_gen_inst_N27), .A2(
        i_weight_addr_gen_inst_n45), .B1(i_weight_addr_gen_inst_N11), .B2(
        i_weight_addr_gen_inst_n46), .ZN(i_weight_addr_gen_inst_n60) );
  INV_X1 i_weight_addr_gen_inst_U55 ( .A(i_weight_addr_gen_inst_n60), .ZN(
        i_weight_addr_gen_inst_n43) );
  AOI22_X1 i_weight_addr_gen_inst_U54 ( .A1(i_weight_addr_gen_inst_N28), .A2(
        i_weight_addr_gen_inst_n45), .B1(i_weight_addr_gen_inst_N12), .B2(
        i_weight_addr_gen_inst_n46), .ZN(i_weight_addr_gen_inst_n59) );
  INV_X1 i_weight_addr_gen_inst_U53 ( .A(i_weight_addr_gen_inst_n59), .ZN(
        i_weight_addr_gen_inst_n42) );
  AOI22_X1 i_weight_addr_gen_inst_U52 ( .A1(i_weight_addr_gen_inst_N29), .A2(
        i_weight_addr_gen_inst_n45), .B1(i_weight_addr_gen_inst_N13), .B2(
        i_weight_addr_gen_inst_n46), .ZN(i_weight_addr_gen_inst_n58) );
  INV_X1 i_weight_addr_gen_inst_U51 ( .A(i_weight_addr_gen_inst_n58), .ZN(
        i_weight_addr_gen_inst_n41) );
  AOI22_X1 i_weight_addr_gen_inst_U50 ( .A1(i_weight_addr_gen_inst_N30), .A2(
        i_weight_addr_gen_inst_n45), .B1(i_weight_addr_gen_inst_N14), .B2(
        i_weight_addr_gen_inst_n46), .ZN(i_weight_addr_gen_inst_n57) );
  INV_X1 i_weight_addr_gen_inst_U49 ( .A(i_weight_addr_gen_inst_n57), .ZN(
        i_weight_addr_gen_inst_n40) );
  AOI22_X1 i_weight_addr_gen_inst_U48 ( .A1(i_weight_addr_gen_inst_N31), .A2(
        i_weight_addr_gen_inst_n45), .B1(i_weight_addr_gen_inst_N15), .B2(
        i_weight_addr_gen_inst_n46), .ZN(i_weight_addr_gen_inst_n56) );
  INV_X1 i_weight_addr_gen_inst_U47 ( .A(i_weight_addr_gen_inst_n56), .ZN(
        i_weight_addr_gen_inst_n39) );
  AOI22_X1 i_weight_addr_gen_inst_U46 ( .A1(i_weight_addr_gen_inst_N32), .A2(
        i_weight_addr_gen_inst_n45), .B1(i_weight_addr_gen_inst_N16), .B2(
        i_weight_addr_gen_inst_n46), .ZN(i_weight_addr_gen_inst_n55) );
  INV_X1 i_weight_addr_gen_inst_U45 ( .A(i_weight_addr_gen_inst_n55), .ZN(
        i_weight_addr_gen_inst_n38) );
  AOI22_X1 i_weight_addr_gen_inst_U44 ( .A1(i_weight_addr_gen_inst_N33), .A2(
        i_weight_addr_gen_inst_n45), .B1(i_weight_addr_gen_inst_N17), .B2(
        i_weight_addr_gen_inst_n46), .ZN(i_weight_addr_gen_inst_n54) );
  INV_X1 i_weight_addr_gen_inst_U43 ( .A(i_weight_addr_gen_inst_n54), .ZN(
        i_weight_addr_gen_inst_n37) );
  AOI22_X1 i_weight_addr_gen_inst_U42 ( .A1(i_weight_addr_gen_inst_N34), .A2(
        i_weight_addr_gen_inst_n45), .B1(i_weight_addr_gen_inst_N18), .B2(
        i_weight_addr_gen_inst_n46), .ZN(i_weight_addr_gen_inst_n53) );
  INV_X1 i_weight_addr_gen_inst_U41 ( .A(i_weight_addr_gen_inst_n53), .ZN(
        i_weight_addr_gen_inst_n36) );
  AOI22_X1 i_weight_addr_gen_inst_U40 ( .A1(i_weight_addr_gen_inst_N35), .A2(
        i_weight_addr_gen_inst_n45), .B1(i_weight_addr_gen_inst_N19), .B2(
        i_weight_addr_gen_inst_n46), .ZN(i_weight_addr_gen_inst_n52) );
  INV_X1 i_weight_addr_gen_inst_U39 ( .A(i_weight_addr_gen_inst_n52), .ZN(
        i_weight_addr_gen_inst_n35) );
  AOI22_X1 i_weight_addr_gen_inst_U38 ( .A1(i_weight_addr_gen_inst_N36), .A2(
        i_weight_addr_gen_inst_n45), .B1(i_weight_addr_gen_inst_N20), .B2(
        i_weight_addr_gen_inst_n46), .ZN(i_weight_addr_gen_inst_n51) );
  INV_X1 i_weight_addr_gen_inst_U37 ( .A(i_weight_addr_gen_inst_n51), .ZN(
        i_weight_addr_gen_inst_n34) );
  AOI22_X1 i_weight_addr_gen_inst_U36 ( .A1(i_weight_addr_gen_inst_N37), .A2(
        i_weight_addr_gen_inst_n45), .B1(i_weight_addr_gen_inst_N21), .B2(
        i_weight_addr_gen_inst_n46), .ZN(i_weight_addr_gen_inst_n50) );
  INV_X1 i_weight_addr_gen_inst_U35 ( .A(i_weight_addr_gen_inst_n50), .ZN(
        i_weight_addr_gen_inst_n33) );
  AOI22_X1 i_weight_addr_gen_inst_U34 ( .A1(i_weight_addr_gen_inst_N38), .A2(
        i_weight_addr_gen_inst_n45), .B1(i_weight_addr_gen_inst_N22), .B2(
        i_weight_addr_gen_inst_n46), .ZN(i_weight_addr_gen_inst_n49) );
  INV_X1 i_weight_addr_gen_inst_U33 ( .A(i_weight_addr_gen_inst_n49), .ZN(
        i_weight_addr_gen_inst_n32) );
  AOI22_X1 i_weight_addr_gen_inst_U32 ( .A1(i_weight_addr_gen_inst_N39), .A2(
        i_weight_addr_gen_inst_n45), .B1(i_weight_addr_gen_inst_N23), .B2(
        i_weight_addr_gen_inst_n46), .ZN(i_weight_addr_gen_inst_n48) );
  INV_X1 i_weight_addr_gen_inst_U31 ( .A(i_weight_addr_gen_inst_n48), .ZN(
        i_weight_addr_gen_inst_n31) );
  AOI22_X1 i_weight_addr_gen_inst_U30 ( .A1(i_weight_addr_gen_inst_N40), .A2(
        i_weight_addr_gen_inst_n45), .B1(i_weight_addr_gen_inst_N24), .B2(
        i_weight_addr_gen_inst_n46), .ZN(i_weight_addr_gen_inst_n47) );
  INV_X1 i_weight_addr_gen_inst_U29 ( .A(i_weight_addr_gen_inst_n47), .ZN(
        i_weight_addr_gen_inst_n30) );
  INV_X1 i_weight_addr_gen_inst_U28 ( .A(n46), .ZN(i_weight_addr_gen_inst_n28)
         );
  BUF_X1 i_weight_addr_gen_inst_U27 ( .A(i_weight_addr_gen_inst_n28), .Z(
        i_weight_addr_gen_inst_n27) );
  BUF_X1 i_weight_addr_gen_inst_U26 ( .A(i_weight_addr_gen_inst_n28), .Z(
        i_weight_addr_gen_inst_n24) );
  BUF_X1 i_weight_addr_gen_inst_U25 ( .A(i_weight_addr_gen_inst_n28), .Z(
        i_weight_addr_gen_inst_n26) );
  NOR2_X2 i_weight_addr_gen_inst_U24 ( .A1(int_c_i_en_weight_addr), .A2(1'b0), 
        .ZN(i_weight_addr_gen_inst_n45) );
  NOR2_X2 i_weight_addr_gen_inst_U22 ( .A1(i_weight_addr_gen_inst_n64), .A2(
        1'b0), .ZN(i_weight_addr_gen_inst_n46) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_14_ ( .D(
        i_weight_addr_gen_inst_n30), .CK(i_weight_addr_gen_inst_net2826), .RN(
        i_weight_addr_gen_inst_n24), .Q(
        i_weight_addr_gen_inst_int_base_addr_14_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_13_ ( .D(
        i_weight_addr_gen_inst_n31), .CK(i_weight_addr_gen_inst_net2826), .RN(
        i_weight_addr_gen_inst_n24), .Q(
        i_weight_addr_gen_inst_int_base_addr_13_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_12_ ( .D(
        i_weight_addr_gen_inst_n32), .CK(i_weight_addr_gen_inst_net2826), .RN(
        i_weight_addr_gen_inst_n24), .Q(
        i_weight_addr_gen_inst_int_base_addr_12_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_11_ ( .D(
        i_weight_addr_gen_inst_n33), .CK(i_weight_addr_gen_inst_net2826), .RN(
        i_weight_addr_gen_inst_n24), .Q(
        i_weight_addr_gen_inst_int_base_addr_11_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_10_ ( .D(
        i_weight_addr_gen_inst_n34), .CK(i_weight_addr_gen_inst_net2826), .RN(
        i_weight_addr_gen_inst_n24), .Q(
        i_weight_addr_gen_inst_int_base_addr_10_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_9_ ( .D(
        i_weight_addr_gen_inst_n35), .CK(i_weight_addr_gen_inst_net2826), .RN(
        i_weight_addr_gen_inst_n24), .Q(
        i_weight_addr_gen_inst_int_base_addr_9_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_8_ ( .D(
        i_weight_addr_gen_inst_n36), .CK(i_weight_addr_gen_inst_net2826), .RN(
        i_weight_addr_gen_inst_n24), .Q(
        i_weight_addr_gen_inst_int_base_addr_8_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_7_ ( .D(
        i_weight_addr_gen_inst_n37), .CK(i_weight_addr_gen_inst_net2826), .RN(
        i_weight_addr_gen_inst_n24), .Q(
        i_weight_addr_gen_inst_int_base_addr_7_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_6_ ( .D(
        i_weight_addr_gen_inst_n38), .CK(i_weight_addr_gen_inst_net2826), .RN(
        i_weight_addr_gen_inst_n24), .Q(
        i_weight_addr_gen_inst_int_base_addr_6_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_5_ ( .D(
        i_weight_addr_gen_inst_n39), .CK(i_weight_addr_gen_inst_net2826), .RN(
        i_weight_addr_gen_inst_n24), .Q(
        i_weight_addr_gen_inst_int_base_addr_5_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_4_ ( .D(
        i_weight_addr_gen_inst_n40), .CK(i_weight_addr_gen_inst_net2826), .RN(
        i_weight_addr_gen_inst_n24), .Q(
        i_weight_addr_gen_inst_int_base_addr_4_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_3_ ( .D(
        i_weight_addr_gen_inst_n41), .CK(i_weight_addr_gen_inst_net2826), .RN(
        i_weight_addr_gen_inst_n24), .Q(
        i_weight_addr_gen_inst_int_base_addr_3_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_2_ ( .D(
        i_weight_addr_gen_inst_n42), .CK(i_weight_addr_gen_inst_net2826), .RN(
        i_weight_addr_gen_inst_n26), .Q(
        i_weight_addr_gen_inst_int_base_addr_2_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_1_ ( .D(
        i_weight_addr_gen_inst_n43), .CK(i_weight_addr_gen_inst_net2826), .RN(
        i_weight_addr_gen_inst_n26), .Q(
        i_weight_addr_gen_inst_int_base_addr_1_) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_0_ ( .D(
        i_weight_addr_gen_inst_n62), .CK(i_weight_addr_gen_inst_net2826), .RN(
        i_weight_addr_gen_inst_n26), .Q(
        i_weight_addr_gen_inst_int_base_addr_0_), .QN(
        i_weight_addr_gen_inst_n6) );
  DFFR_X1 i_weight_addr_gen_inst_int_base_addr_reg_15_ ( .D(
        i_weight_addr_gen_inst_n29), .CK(i_weight_addr_gen_inst_net2826), .RN(
        i_weight_addr_gen_inst_n26), .Q(
        i_weight_addr_gen_inst_int_base_addr_15_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_15_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n63), .SE(i_weight_addr_gen_inst_N94), .CK(
        i_weight_addr_gen_inst_net2832), .RN(i_weight_addr_gen_inst_n26), .Q(
        i_weight_addr_gen_inst_int_offs_addr_15_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_14_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n63), .SE(i_weight_addr_gen_inst_N93), .CK(
        i_weight_addr_gen_inst_net2832), .RN(i_weight_addr_gen_inst_n26), .Q(
        i_weight_addr_gen_inst_int_offs_addr_14_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_13_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n63), .SE(i_weight_addr_gen_inst_N92), .CK(
        i_weight_addr_gen_inst_net2832), .RN(i_weight_addr_gen_inst_n26), .Q(
        i_weight_addr_gen_inst_int_offs_addr_13_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_12_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n63), .SE(i_weight_addr_gen_inst_N91), .CK(
        i_weight_addr_gen_inst_net2832), .RN(i_weight_addr_gen_inst_n26), .Q(
        i_weight_addr_gen_inst_int_offs_addr_12_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_11_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n63), .SE(i_weight_addr_gen_inst_N90), .CK(
        i_weight_addr_gen_inst_net2832), .RN(i_weight_addr_gen_inst_n26), .Q(
        i_weight_addr_gen_inst_int_offs_addr_11_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_10_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n63), .SE(i_weight_addr_gen_inst_N89), .CK(
        i_weight_addr_gen_inst_net2832), .RN(i_weight_addr_gen_inst_n26), .Q(
        i_weight_addr_gen_inst_int_offs_addr_10_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_9_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n63), .SE(i_weight_addr_gen_inst_N88), .CK(
        i_weight_addr_gen_inst_net2832), .RN(i_weight_addr_gen_inst_n26), .Q(
        i_weight_addr_gen_inst_int_offs_addr_9_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_8_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n63), .SE(i_weight_addr_gen_inst_N87), .CK(
        i_weight_addr_gen_inst_net2832), .RN(i_weight_addr_gen_inst_n26), .Q(
        i_weight_addr_gen_inst_int_offs_addr_8_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_7_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n63), .SE(i_weight_addr_gen_inst_N86), .CK(
        i_weight_addr_gen_inst_net2832), .RN(i_weight_addr_gen_inst_n26), .Q(
        i_weight_addr_gen_inst_int_offs_addr_7_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_6_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n63), .SE(i_weight_addr_gen_inst_N85), .CK(
        i_weight_addr_gen_inst_net2832), .RN(i_weight_addr_gen_inst_n27), .Q(
        i_weight_addr_gen_inst_int_offs_addr_6_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_5_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n63), .SE(i_weight_addr_gen_inst_N84), .CK(
        i_weight_addr_gen_inst_net2832), .RN(i_weight_addr_gen_inst_n27), .Q(
        i_weight_addr_gen_inst_int_offs_addr_5_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_4_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n63), .SE(i_weight_addr_gen_inst_N83), .CK(
        i_weight_addr_gen_inst_net2832), .RN(i_weight_addr_gen_inst_n27), .Q(
        i_weight_addr_gen_inst_int_offs_addr_4_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_3_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n63), .SE(i_weight_addr_gen_inst_N82), .CK(
        i_weight_addr_gen_inst_net2832), .RN(i_weight_addr_gen_inst_n27), .Q(
        i_weight_addr_gen_inst_int_offs_addr_3_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_2_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n63), .SE(i_weight_addr_gen_inst_N81), .CK(
        i_weight_addr_gen_inst_net2832), .RN(i_weight_addr_gen_inst_n27), .Q(
        i_weight_addr_gen_inst_int_offs_addr_2_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_1_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n63), .SE(i_weight_addr_gen_inst_N80), .CK(
        i_weight_addr_gen_inst_net2832), .RN(i_weight_addr_gen_inst_n27), .Q(
        i_weight_addr_gen_inst_int_offs_addr_1_) );
  SDFFR_X1 i_weight_addr_gen_inst_int_offs_addr_reg_0_ ( .D(1'b0), .SI(
        i_weight_addr_gen_inst_n63), .SE(i_weight_addr_gen_inst_N79), .CK(
        i_weight_addr_gen_inst_net2832), .RN(i_weight_addr_gen_inst_n27), .Q(
        i_weight_addr_gen_inst_n5) );
  CLKGATETST_X1 i_weight_addr_gen_inst_clk_gate_int_base_addr_reg_latch ( .CK(
        ck), .E(i_weight_addr_gen_inst_N58), .SE(1'b0), .GCK(
        i_weight_addr_gen_inst_net2826) );
  CLKGATETST_X1 i_weight_addr_gen_inst_clk_gate_int_offs_addr_reg_latch ( .CK(
        ck), .E(i_weight_addr_gen_inst_N95), .SE(1'b0), .GCK(
        i_weight_addr_gen_inst_net2832) );
  XOR2_X1 i_weight_addr_gen_inst_add_61_U2 ( .A(1'b1), .B(
        i_weight_addr_gen_inst_n5), .Z(i_weight_addr_gen_inst_N79) );
  AND2_X1 i_weight_addr_gen_inst_add_61_U1 ( .A1(1'b1), .A2(
        i_weight_addr_gen_inst_n5), .ZN(i_weight_addr_gen_inst_add_61_n1) );
  FA_X1 i_weight_addr_gen_inst_add_61_U1_1 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_1_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_61_n1), .CO(
        i_weight_addr_gen_inst_add_61_carry[2]), .S(i_weight_addr_gen_inst_N80) );
  FA_X1 i_weight_addr_gen_inst_add_61_U1_2 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_2_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_61_carry[2]), .CO(
        i_weight_addr_gen_inst_add_61_carry[3]), .S(i_weight_addr_gen_inst_N81) );
  FA_X1 i_weight_addr_gen_inst_add_61_U1_3 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_3_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_61_carry[3]), .CO(
        i_weight_addr_gen_inst_add_61_carry[4]), .S(i_weight_addr_gen_inst_N82) );
  FA_X1 i_weight_addr_gen_inst_add_61_U1_4 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_4_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_61_carry[4]), .CO(
        i_weight_addr_gen_inst_add_61_carry[5]), .S(i_weight_addr_gen_inst_N83) );
  FA_X1 i_weight_addr_gen_inst_add_61_U1_5 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_5_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_61_carry[5]), .CO(
        i_weight_addr_gen_inst_add_61_carry[6]), .S(i_weight_addr_gen_inst_N84) );
  FA_X1 i_weight_addr_gen_inst_add_61_U1_6 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_6_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_61_carry[6]), .CO(
        i_weight_addr_gen_inst_add_61_carry[7]), .S(i_weight_addr_gen_inst_N85) );
  FA_X1 i_weight_addr_gen_inst_add_61_U1_7 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_7_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_61_carry[7]), .CO(
        i_weight_addr_gen_inst_add_61_carry[8]), .S(i_weight_addr_gen_inst_N86) );
  FA_X1 i_weight_addr_gen_inst_add_61_U1_8 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_8_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_61_carry[8]), .CO(
        i_weight_addr_gen_inst_add_61_carry[9]), .S(i_weight_addr_gen_inst_N87) );
  FA_X1 i_weight_addr_gen_inst_add_61_U1_9 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_9_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_61_carry[9]), .CO(
        i_weight_addr_gen_inst_add_61_carry[10]), .S(
        i_weight_addr_gen_inst_N88) );
  FA_X1 i_weight_addr_gen_inst_add_61_U1_10 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_10_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_61_carry[10]), .CO(
        i_weight_addr_gen_inst_add_61_carry[11]), .S(
        i_weight_addr_gen_inst_N89) );
  FA_X1 i_weight_addr_gen_inst_add_61_U1_11 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_11_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_61_carry[11]), .CO(
        i_weight_addr_gen_inst_add_61_carry[12]), .S(
        i_weight_addr_gen_inst_N90) );
  FA_X1 i_weight_addr_gen_inst_add_61_U1_12 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_12_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_61_carry[12]), .CO(
        i_weight_addr_gen_inst_add_61_carry[13]), .S(
        i_weight_addr_gen_inst_N91) );
  FA_X1 i_weight_addr_gen_inst_add_61_U1_13 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_13_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_61_carry[13]), .CO(
        i_weight_addr_gen_inst_add_61_carry[14]), .S(
        i_weight_addr_gen_inst_N92) );
  FA_X1 i_weight_addr_gen_inst_add_61_U1_14 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_14_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_61_carry[14]), .CO(
        i_weight_addr_gen_inst_add_61_carry[15]), .S(
        i_weight_addr_gen_inst_N93) );
  FA_X1 i_weight_addr_gen_inst_add_61_U1_15 ( .A(
        i_weight_addr_gen_inst_int_offs_addr_15_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_61_carry[15]), .S(
        i_weight_addr_gen_inst_N94) );
  AND2_X1 i_weight_addr_gen_inst_add_46_U2 ( .A1(1'b0), .A2(
        i_weight_addr_gen_inst_int_base_addr_0_), .ZN(
        i_weight_addr_gen_inst_add_46_n2) );
  XOR2_X1 i_weight_addr_gen_inst_add_46_U1 ( .A(1'b0), .B(
        i_weight_addr_gen_inst_int_base_addr_0_), .Z(
        i_weight_addr_gen_inst_N26) );
  FA_X1 i_weight_addr_gen_inst_add_46_U1_1 ( .A(
        i_weight_addr_gen_inst_int_base_addr_1_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_46_n2), .CO(
        i_weight_addr_gen_inst_add_46_carry[2]), .S(i_weight_addr_gen_inst_N27) );
  FA_X1 i_weight_addr_gen_inst_add_46_U1_2 ( .A(
        i_weight_addr_gen_inst_int_base_addr_2_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_46_carry[2]), .CO(
        i_weight_addr_gen_inst_add_46_carry[3]), .S(i_weight_addr_gen_inst_N28) );
  FA_X1 i_weight_addr_gen_inst_add_46_U1_3 ( .A(
        i_weight_addr_gen_inst_int_base_addr_3_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_46_carry[3]), .CO(
        i_weight_addr_gen_inst_add_46_carry[4]), .S(i_weight_addr_gen_inst_N29) );
  FA_X1 i_weight_addr_gen_inst_add_46_U1_4 ( .A(
        i_weight_addr_gen_inst_int_base_addr_4_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_46_carry[4]), .CO(
        i_weight_addr_gen_inst_add_46_carry[5]), .S(i_weight_addr_gen_inst_N30) );
  FA_X1 i_weight_addr_gen_inst_add_46_U1_5 ( .A(
        i_weight_addr_gen_inst_int_base_addr_5_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_46_carry[5]), .CO(
        i_weight_addr_gen_inst_add_46_carry[6]), .S(i_weight_addr_gen_inst_N31) );
  FA_X1 i_weight_addr_gen_inst_add_46_U1_6 ( .A(
        i_weight_addr_gen_inst_int_base_addr_6_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_46_carry[6]), .CO(
        i_weight_addr_gen_inst_add_46_carry[7]), .S(i_weight_addr_gen_inst_N32) );
  FA_X1 i_weight_addr_gen_inst_add_46_U1_7 ( .A(
        i_weight_addr_gen_inst_int_base_addr_7_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_46_carry[7]), .CO(
        i_weight_addr_gen_inst_add_46_carry[8]), .S(i_weight_addr_gen_inst_N33) );
  FA_X1 i_weight_addr_gen_inst_add_46_U1_8 ( .A(
        i_weight_addr_gen_inst_int_base_addr_8_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_46_carry[8]), .CO(
        i_weight_addr_gen_inst_add_46_carry[9]), .S(i_weight_addr_gen_inst_N34) );
  FA_X1 i_weight_addr_gen_inst_add_46_U1_9 ( .A(
        i_weight_addr_gen_inst_int_base_addr_9_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_46_carry[9]), .CO(
        i_weight_addr_gen_inst_add_46_carry[10]), .S(
        i_weight_addr_gen_inst_N35) );
  FA_X1 i_weight_addr_gen_inst_add_46_U1_10 ( .A(
        i_weight_addr_gen_inst_int_base_addr_10_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_46_carry[10]), .CO(
        i_weight_addr_gen_inst_add_46_carry[11]), .S(
        i_weight_addr_gen_inst_N36) );
  FA_X1 i_weight_addr_gen_inst_add_46_U1_11 ( .A(
        i_weight_addr_gen_inst_int_base_addr_11_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_46_carry[11]), .CO(
        i_weight_addr_gen_inst_add_46_carry[12]), .S(
        i_weight_addr_gen_inst_N37) );
  FA_X1 i_weight_addr_gen_inst_add_46_U1_12 ( .A(
        i_weight_addr_gen_inst_int_base_addr_12_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_46_carry[12]), .CO(
        i_weight_addr_gen_inst_add_46_carry[13]), .S(
        i_weight_addr_gen_inst_N38) );
  FA_X1 i_weight_addr_gen_inst_add_46_U1_13 ( .A(
        i_weight_addr_gen_inst_int_base_addr_13_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_46_carry[13]), .CO(
        i_weight_addr_gen_inst_add_46_carry[14]), .S(
        i_weight_addr_gen_inst_N39) );
  FA_X1 i_weight_addr_gen_inst_add_46_U1_14 ( .A(
        i_weight_addr_gen_inst_int_base_addr_14_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_46_carry[14]), .CO(
        i_weight_addr_gen_inst_add_46_carry[15]), .S(
        i_weight_addr_gen_inst_N40) );
  FA_X1 i_weight_addr_gen_inst_add_46_U1_15 ( .A(
        i_weight_addr_gen_inst_int_base_addr_15_), .B(1'b0), .CI(
        i_weight_addr_gen_inst_add_46_carry[15]), .S(
        i_weight_addr_gen_inst_N41) );
  AND2_X1 i_weight_addr_gen_inst_add_44_U2 ( .A1(1'b0), .A2(i_weight_addr[0]), 
        .ZN(i_weight_addr_gen_inst_add_44_n2) );
  XOR2_X1 i_weight_addr_gen_inst_add_44_U1 ( .A(1'b0), .B(i_weight_addr[0]), 
        .Z(i_weight_addr_gen_inst_N10) );
  FA_X1 i_weight_addr_gen_inst_add_44_U1_1 ( .A(i_weight_addr[1]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_44_n2), .CO(
        i_weight_addr_gen_inst_add_44_carry[2]), .S(i_weight_addr_gen_inst_N11) );
  FA_X1 i_weight_addr_gen_inst_add_44_U1_2 ( .A(i_weight_addr[2]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_44_carry[2]), .CO(
        i_weight_addr_gen_inst_add_44_carry[3]), .S(i_weight_addr_gen_inst_N12) );
  FA_X1 i_weight_addr_gen_inst_add_44_U1_3 ( .A(i_weight_addr[3]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_44_carry[3]), .CO(
        i_weight_addr_gen_inst_add_44_carry[4]), .S(i_weight_addr_gen_inst_N13) );
  FA_X1 i_weight_addr_gen_inst_add_44_U1_4 ( .A(i_weight_addr[4]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_44_carry[4]), .CO(
        i_weight_addr_gen_inst_add_44_carry[5]), .S(i_weight_addr_gen_inst_N14) );
  FA_X1 i_weight_addr_gen_inst_add_44_U1_5 ( .A(i_weight_addr[5]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_44_carry[5]), .CO(
        i_weight_addr_gen_inst_add_44_carry[6]), .S(i_weight_addr_gen_inst_N15) );
  FA_X1 i_weight_addr_gen_inst_add_44_U1_6 ( .A(i_weight_addr[6]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_44_carry[6]), .CO(
        i_weight_addr_gen_inst_add_44_carry[7]), .S(i_weight_addr_gen_inst_N16) );
  FA_X1 i_weight_addr_gen_inst_add_44_U1_7 ( .A(i_weight_addr[7]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_44_carry[7]), .CO(
        i_weight_addr_gen_inst_add_44_carry[8]), .S(i_weight_addr_gen_inst_N17) );
  FA_X1 i_weight_addr_gen_inst_add_44_U1_8 ( .A(i_weight_addr[8]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_44_carry[8]), .CO(
        i_weight_addr_gen_inst_add_44_carry[9]), .S(i_weight_addr_gen_inst_N18) );
  FA_X1 i_weight_addr_gen_inst_add_44_U1_9 ( .A(i_weight_addr[9]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_44_carry[9]), .CO(
        i_weight_addr_gen_inst_add_44_carry[10]), .S(
        i_weight_addr_gen_inst_N19) );
  FA_X1 i_weight_addr_gen_inst_add_44_U1_10 ( .A(i_weight_addr[10]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_44_carry[10]), .CO(
        i_weight_addr_gen_inst_add_44_carry[11]), .S(
        i_weight_addr_gen_inst_N20) );
  FA_X1 i_weight_addr_gen_inst_add_44_U1_11 ( .A(i_weight_addr[11]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_44_carry[11]), .CO(
        i_weight_addr_gen_inst_add_44_carry[12]), .S(
        i_weight_addr_gen_inst_N21) );
  FA_X1 i_weight_addr_gen_inst_add_44_U1_12 ( .A(i_weight_addr[12]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_44_carry[12]), .CO(
        i_weight_addr_gen_inst_add_44_carry[13]), .S(
        i_weight_addr_gen_inst_N22) );
  FA_X1 i_weight_addr_gen_inst_add_44_U1_13 ( .A(i_weight_addr[13]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_44_carry[13]), .CO(
        i_weight_addr_gen_inst_add_44_carry[14]), .S(
        i_weight_addr_gen_inst_N23) );
  FA_X1 i_weight_addr_gen_inst_add_44_U1_14 ( .A(i_weight_addr[14]), .B(1'b0), 
        .CI(i_weight_addr_gen_inst_add_44_carry[14]), .CO(
        i_weight_addr_gen_inst_add_44_carry[15]), .S(
        i_weight_addr_gen_inst_N24) );
  FA_X1 i_weight_addr_gen_inst_add_44_U1_15 ( .A(i_weight_addr_gen_inst_n8), 
        .B(1'b0), .CI(i_weight_addr_gen_inst_add_44_carry[15]), .S(
        i_weight_addr_gen_inst_N25) );
  XOR2_X1 i_weight_addr_gen_inst_add_32_U49 ( .A(i_weight_addr_gen_inst_n5), 
        .B(i_weight_addr_gen_inst_n7), .Z(i_weight_addr[0]) );
  AND2_X1 i_weight_addr_gen_inst_add_32_U48 ( .A1(i_weight_addr_gen_inst_n5), 
        .A2(i_weight_addr_gen_inst_n7), .ZN(i_weight_addr_gen_inst_add_32_n33)
         );
  NAND3_X1 i_weight_addr_gen_inst_add_32_U47 ( .A1(
        i_weight_addr_gen_inst_add_32_n30), .A2(
        i_weight_addr_gen_inst_add_32_n31), .A3(
        i_weight_addr_gen_inst_add_32_n32), .ZN(
        i_weight_addr_gen_inst_add_32_carry_13_) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U46 ( .A1(
        i_weight_addr_gen_inst_int_base_addr_12_), .A2(
        i_weight_addr_gen_inst_int_offs_addr_12_), .ZN(
        i_weight_addr_gen_inst_add_32_n32) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U45 ( .A1(
        i_weight_addr_gen_inst_add_32_n18), .A2(
        i_weight_addr_gen_inst_int_offs_addr_12_), .ZN(
        i_weight_addr_gen_inst_add_32_n31) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U44 ( .A1(
        i_weight_addr_gen_inst_add_32_n19), .A2(
        i_weight_addr_gen_inst_int_base_addr_12_), .ZN(
        i_weight_addr_gen_inst_add_32_n30) );
  XOR2_X1 i_weight_addr_gen_inst_add_32_U43 ( .A(
        i_weight_addr_gen_inst_add_32_carry_12_), .B(
        i_weight_addr_gen_inst_add_32_n29), .Z(i_weight_addr[12]) );
  XOR2_X1 i_weight_addr_gen_inst_add_32_U42 ( .A(
        i_weight_addr_gen_inst_int_base_addr_12_), .B(
        i_weight_addr_gen_inst_int_offs_addr_12_), .Z(
        i_weight_addr_gen_inst_add_32_n29) );
  XNOR2_X1 i_weight_addr_gen_inst_add_32_U41 ( .A(
        i_weight_addr_gen_inst_int_base_addr_15_), .B(
        i_weight_addr_gen_inst_int_offs_addr_15_), .ZN(
        i_weight_addr_gen_inst_add_32_n28) );
  XNOR2_X1 i_weight_addr_gen_inst_add_32_U40 ( .A(
        i_weight_addr_gen_inst_add_32_carry_15_), .B(
        i_weight_addr_gen_inst_add_32_n28), .ZN(i_weight_addr[15]) );
  NAND3_X1 i_weight_addr_gen_inst_add_32_U39 ( .A1(
        i_weight_addr_gen_inst_add_32_n25), .A2(
        i_weight_addr_gen_inst_add_32_n26), .A3(
        i_weight_addr_gen_inst_add_32_n27), .ZN(
        i_weight_addr_gen_inst_add_32_carry_12_) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U38 ( .A1(
        i_weight_addr_gen_inst_int_base_addr_11_), .A2(
        i_weight_addr_gen_inst_int_offs_addr_11_), .ZN(
        i_weight_addr_gen_inst_add_32_n27) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U37 ( .A1(
        i_weight_addr_gen_inst_add_32_carry_11_), .A2(
        i_weight_addr_gen_inst_int_offs_addr_11_), .ZN(
        i_weight_addr_gen_inst_add_32_n26) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U36 ( .A1(
        i_weight_addr_gen_inst_add_32_carry_11_), .A2(
        i_weight_addr_gen_inst_int_base_addr_11_), .ZN(
        i_weight_addr_gen_inst_add_32_n25) );
  XOR2_X1 i_weight_addr_gen_inst_add_32_U35 ( .A(
        i_weight_addr_gen_inst_add_32_carry_11_), .B(
        i_weight_addr_gen_inst_add_32_n24), .Z(i_weight_addr[11]) );
  XOR2_X1 i_weight_addr_gen_inst_add_32_U34 ( .A(
        i_weight_addr_gen_inst_int_base_addr_11_), .B(
        i_weight_addr_gen_inst_int_offs_addr_11_), .Z(
        i_weight_addr_gen_inst_add_32_n24) );
  NAND3_X1 i_weight_addr_gen_inst_add_32_U33 ( .A1(
        i_weight_addr_gen_inst_add_32_n21), .A2(
        i_weight_addr_gen_inst_add_32_n22), .A3(
        i_weight_addr_gen_inst_add_32_n23), .ZN(
        i_weight_addr_gen_inst_add_32_carry_9_) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U32 ( .A1(
        i_weight_addr_gen_inst_int_base_addr_8_), .A2(
        i_weight_addr_gen_inst_int_offs_addr_8_), .ZN(
        i_weight_addr_gen_inst_add_32_n23) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U31 ( .A1(
        i_weight_addr_gen_inst_add_32_carry_8_), .A2(
        i_weight_addr_gen_inst_int_offs_addr_8_), .ZN(
        i_weight_addr_gen_inst_add_32_n22) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U30 ( .A1(
        i_weight_addr_gen_inst_add_32_carry_8_), .A2(
        i_weight_addr_gen_inst_int_base_addr_8_), .ZN(
        i_weight_addr_gen_inst_add_32_n21) );
  XOR2_X1 i_weight_addr_gen_inst_add_32_U29 ( .A(
        i_weight_addr_gen_inst_add_32_carry_8_), .B(
        i_weight_addr_gen_inst_add_32_n20), .Z(i_weight_addr[8]) );
  XOR2_X1 i_weight_addr_gen_inst_add_32_U28 ( .A(
        i_weight_addr_gen_inst_int_base_addr_8_), .B(
        i_weight_addr_gen_inst_int_offs_addr_8_), .Z(
        i_weight_addr_gen_inst_add_32_n20) );
  NAND3_X1 i_weight_addr_gen_inst_add_32_U27 ( .A1(
        i_weight_addr_gen_inst_add_32_n25), .A2(
        i_weight_addr_gen_inst_add_32_n26), .A3(
        i_weight_addr_gen_inst_add_32_n27), .ZN(
        i_weight_addr_gen_inst_add_32_n19) );
  NAND3_X1 i_weight_addr_gen_inst_add_32_U26 ( .A1(
        i_weight_addr_gen_inst_add_32_n25), .A2(
        i_weight_addr_gen_inst_add_32_n26), .A3(
        i_weight_addr_gen_inst_add_32_n27), .ZN(
        i_weight_addr_gen_inst_add_32_n18) );
  NAND3_X1 i_weight_addr_gen_inst_add_32_U25 ( .A1(
        i_weight_addr_gen_inst_add_32_n15), .A2(
        i_weight_addr_gen_inst_add_32_n16), .A3(
        i_weight_addr_gen_inst_add_32_n17), .ZN(
        i_weight_addr_gen_inst_add_32_carry_8_) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U24 ( .A1(
        i_weight_addr_gen_inst_int_base_addr_7_), .A2(
        i_weight_addr_gen_inst_int_offs_addr_7_), .ZN(
        i_weight_addr_gen_inst_add_32_n17) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U23 ( .A1(
        i_weight_addr_gen_inst_add_32_carry_7_), .A2(
        i_weight_addr_gen_inst_int_offs_addr_7_), .ZN(
        i_weight_addr_gen_inst_add_32_n16) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U22 ( .A1(
        i_weight_addr_gen_inst_add_32_carry_7_), .A2(
        i_weight_addr_gen_inst_int_base_addr_7_), .ZN(
        i_weight_addr_gen_inst_add_32_n15) );
  XOR2_X1 i_weight_addr_gen_inst_add_32_U21 ( .A(
        i_weight_addr_gen_inst_add_32_carry_7_), .B(
        i_weight_addr_gen_inst_add_32_n14), .Z(i_weight_addr[7]) );
  XOR2_X1 i_weight_addr_gen_inst_add_32_U20 ( .A(
        i_weight_addr_gen_inst_int_base_addr_7_), .B(
        i_weight_addr_gen_inst_int_offs_addr_7_), .Z(
        i_weight_addr_gen_inst_add_32_n14) );
  NAND3_X1 i_weight_addr_gen_inst_add_32_U19 ( .A1(
        i_weight_addr_gen_inst_add_32_n11), .A2(
        i_weight_addr_gen_inst_add_32_n12), .A3(
        i_weight_addr_gen_inst_add_32_n13), .ZN(
        i_weight_addr_gen_inst_add_32_carry_15_) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U18 ( .A1(
        i_weight_addr_gen_inst_int_base_addr_14_), .A2(
        i_weight_addr_gen_inst_int_offs_addr_14_), .ZN(
        i_weight_addr_gen_inst_add_32_n13) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U17 ( .A1(
        i_weight_addr_gen_inst_add_32_carry_14_), .A2(
        i_weight_addr_gen_inst_int_offs_addr_14_), .ZN(
        i_weight_addr_gen_inst_add_32_n12) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U16 ( .A1(
        i_weight_addr_gen_inst_add_32_carry_14_), .A2(
        i_weight_addr_gen_inst_int_base_addr_14_), .ZN(
        i_weight_addr_gen_inst_add_32_n11) );
  XOR2_X1 i_weight_addr_gen_inst_add_32_U15 ( .A(
        i_weight_addr_gen_inst_add_32_n1), .B(
        i_weight_addr_gen_inst_add_32_n10), .Z(i_weight_addr[14]) );
  XOR2_X1 i_weight_addr_gen_inst_add_32_U14 ( .A(
        i_weight_addr_gen_inst_int_base_addr_14_), .B(
        i_weight_addr_gen_inst_int_offs_addr_14_), .Z(
        i_weight_addr_gen_inst_add_32_n10) );
  NAND3_X1 i_weight_addr_gen_inst_add_32_U13 ( .A1(
        i_weight_addr_gen_inst_add_32_n7), .A2(
        i_weight_addr_gen_inst_add_32_n8), .A3(
        i_weight_addr_gen_inst_add_32_n9), .ZN(
        i_weight_addr_gen_inst_add_32_carry_14_) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U12 ( .A1(
        i_weight_addr_gen_inst_int_base_addr_13_), .A2(
        i_weight_addr_gen_inst_int_offs_addr_13_), .ZN(
        i_weight_addr_gen_inst_add_32_n9) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U11 ( .A1(
        i_weight_addr_gen_inst_add_32_carry_13_), .A2(
        i_weight_addr_gen_inst_int_offs_addr_13_), .ZN(
        i_weight_addr_gen_inst_add_32_n8) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U10 ( .A1(
        i_weight_addr_gen_inst_add_32_carry_13_), .A2(
        i_weight_addr_gen_inst_int_base_addr_13_), .ZN(
        i_weight_addr_gen_inst_add_32_n7) );
  XOR2_X1 i_weight_addr_gen_inst_add_32_U9 ( .A(
        i_weight_addr_gen_inst_add_32_carry_13_), .B(
        i_weight_addr_gen_inst_add_32_n6), .Z(i_weight_addr[13]) );
  XOR2_X1 i_weight_addr_gen_inst_add_32_U8 ( .A(
        i_weight_addr_gen_inst_int_base_addr_13_), .B(
        i_weight_addr_gen_inst_int_offs_addr_13_), .Z(
        i_weight_addr_gen_inst_add_32_n6) );
  NAND3_X1 i_weight_addr_gen_inst_add_32_U7 ( .A1(
        i_weight_addr_gen_inst_add_32_n3), .A2(
        i_weight_addr_gen_inst_add_32_n4), .A3(
        i_weight_addr_gen_inst_add_32_n5), .ZN(
        i_weight_addr_gen_inst_add_32_carry_7_) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U6 ( .A1(
        i_weight_addr_gen_inst_int_base_addr_6_), .A2(
        i_weight_addr_gen_inst_int_offs_addr_6_), .ZN(
        i_weight_addr_gen_inst_add_32_n5) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U5 ( .A1(
        i_weight_addr_gen_inst_add_32_carry_6_), .A2(
        i_weight_addr_gen_inst_int_offs_addr_6_), .ZN(
        i_weight_addr_gen_inst_add_32_n4) );
  NAND2_X1 i_weight_addr_gen_inst_add_32_U4 ( .A1(
        i_weight_addr_gen_inst_add_32_carry_6_), .A2(
        i_weight_addr_gen_inst_int_base_addr_6_), .ZN(
        i_weight_addr_gen_inst_add_32_n3) );
  XOR2_X1 i_weight_addr_gen_inst_add_32_U3 ( .A(
        i_weight_addr_gen_inst_add_32_carry_6_), .B(
        i_weight_addr_gen_inst_add_32_n2), .Z(i_weight_addr[6]) );
  XOR2_X1 i_weight_addr_gen_inst_add_32_U2 ( .A(
        i_weight_addr_gen_inst_int_base_addr_6_), .B(
        i_weight_addr_gen_inst_int_offs_addr_6_), .Z(
        i_weight_addr_gen_inst_add_32_n2) );
  CLKBUF_X1 i_weight_addr_gen_inst_add_32_U1 ( .A(
        i_weight_addr_gen_inst_add_32_carry_14_), .Z(
        i_weight_addr_gen_inst_add_32_n1) );
  FA_X1 i_weight_addr_gen_inst_add_32_U1_1 ( .A(
        i_weight_addr_gen_inst_int_base_addr_1_), .B(
        i_weight_addr_gen_inst_int_offs_addr_1_), .CI(
        i_weight_addr_gen_inst_add_32_n33), .CO(
        i_weight_addr_gen_inst_add_32_carry_2_), .S(i_weight_addr[1]) );
  FA_X1 i_weight_addr_gen_inst_add_32_U1_2 ( .A(
        i_weight_addr_gen_inst_int_base_addr_2_), .B(
        i_weight_addr_gen_inst_int_offs_addr_2_), .CI(
        i_weight_addr_gen_inst_add_32_carry_2_), .CO(
        i_weight_addr_gen_inst_add_32_carry_3_), .S(i_weight_addr[2]) );
  FA_X1 i_weight_addr_gen_inst_add_32_U1_3 ( .A(
        i_weight_addr_gen_inst_int_base_addr_3_), .B(
        i_weight_addr_gen_inst_int_offs_addr_3_), .CI(
        i_weight_addr_gen_inst_add_32_carry_3_), .CO(
        i_weight_addr_gen_inst_add_32_carry_4_), .S(i_weight_addr[3]) );
  FA_X1 i_weight_addr_gen_inst_add_32_U1_4 ( .A(
        i_weight_addr_gen_inst_int_base_addr_4_), .B(
        i_weight_addr_gen_inst_int_offs_addr_4_), .CI(
        i_weight_addr_gen_inst_add_32_carry_4_), .CO(
        i_weight_addr_gen_inst_add_32_carry_5_), .S(i_weight_addr[4]) );
  FA_X1 i_weight_addr_gen_inst_add_32_U1_5 ( .A(
        i_weight_addr_gen_inst_int_base_addr_5_), .B(
        i_weight_addr_gen_inst_int_offs_addr_5_), .CI(
        i_weight_addr_gen_inst_add_32_carry_5_), .CO(
        i_weight_addr_gen_inst_add_32_carry_6_), .S(i_weight_addr[5]) );
  FA_X1 i_weight_addr_gen_inst_add_32_U1_9 ( .A(
        i_weight_addr_gen_inst_int_base_addr_9_), .B(
        i_weight_addr_gen_inst_int_offs_addr_9_), .CI(
        i_weight_addr_gen_inst_add_32_carry_9_), .CO(
        i_weight_addr_gen_inst_add_32_carry_10_), .S(i_weight_addr[9]) );
  FA_X1 i_weight_addr_gen_inst_add_32_U1_10 ( .A(
        i_weight_addr_gen_inst_int_base_addr_10_), .B(
        i_weight_addr_gen_inst_int_offs_addr_10_), .CI(
        i_weight_addr_gen_inst_add_32_carry_10_), .CO(
        i_weight_addr_gen_inst_add_32_carry_11_), .S(i_weight_addr[10]) );
  INV_X1 i_data_even_addr_gen_inst_U44 ( .A(n47), .ZN(
        i_data_even_addr_gen_inst_n6) );
  INV_X1 i_data_even_addr_gen_inst_U43 ( .A(n47), .ZN(
        i_data_even_addr_gen_inst_n5) );
  AOI22_X1 i_data_even_addr_gen_inst_U42 ( .A1(i_data_even_addr_gen_inst_N29), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N19), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n32)
         );
  INV_X1 i_data_even_addr_gen_inst_U41 ( .A(i_data_even_addr_gen_inst_n32), 
        .ZN(i_data_even_addr_gen_inst_n7) );
  OR2_X1 i_data_even_addr_gen_inst_U40 ( .A1(n59), .A2(ctrl_ldh_v_n), .ZN(
        i_data_even_addr_gen_inst_N65) );
  AOI22_X1 i_data_even_addr_gen_inst_U39 ( .A1(i_data_even_addr_gen_inst_N20), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N10), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n43)
         );
  INV_X1 i_data_even_addr_gen_inst_U38 ( .A(i_data_even_addr_gen_inst_n43), 
        .ZN(i_data_even_addr_gen_inst_n26) );
  AOI22_X1 i_data_even_addr_gen_inst_U37 ( .A1(i_data_even_addr_gen_inst_N21), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N11), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n42)
         );
  INV_X1 i_data_even_addr_gen_inst_U36 ( .A(i_data_even_addr_gen_inst_n42), 
        .ZN(i_data_even_addr_gen_inst_n25) );
  AOI22_X1 i_data_even_addr_gen_inst_U35 ( .A1(i_data_even_addr_gen_inst_N22), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N12), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n41)
         );
  INV_X1 i_data_even_addr_gen_inst_U34 ( .A(i_data_even_addr_gen_inst_n41), 
        .ZN(i_data_even_addr_gen_inst_n24) );
  AOI22_X1 i_data_even_addr_gen_inst_U33 ( .A1(i_data_even_addr_gen_inst_N23), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N13), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n40)
         );
  INV_X1 i_data_even_addr_gen_inst_U32 ( .A(i_data_even_addr_gen_inst_n40), 
        .ZN(i_data_even_addr_gen_inst_n23) );
  AOI22_X1 i_data_even_addr_gen_inst_U31 ( .A1(i_data_even_addr_gen_inst_N24), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N14), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n39)
         );
  INV_X1 i_data_even_addr_gen_inst_U30 ( .A(i_data_even_addr_gen_inst_n39), 
        .ZN(i_data_even_addr_gen_inst_n22) );
  AOI22_X1 i_data_even_addr_gen_inst_U29 ( .A1(i_data_even_addr_gen_inst_N25), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N15), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n38)
         );
  INV_X1 i_data_even_addr_gen_inst_U28 ( .A(i_data_even_addr_gen_inst_n38), 
        .ZN(i_data_even_addr_gen_inst_n21) );
  AOI22_X1 i_data_even_addr_gen_inst_U27 ( .A1(i_data_even_addr_gen_inst_N26), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N16), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n37)
         );
  INV_X1 i_data_even_addr_gen_inst_U26 ( .A(i_data_even_addr_gen_inst_n37), 
        .ZN(i_data_even_addr_gen_inst_n20) );
  AOI22_X1 i_data_even_addr_gen_inst_U25 ( .A1(i_data_even_addr_gen_inst_N27), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N17), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n36)
         );
  INV_X1 i_data_even_addr_gen_inst_U24 ( .A(i_data_even_addr_gen_inst_n36), 
        .ZN(i_data_even_addr_gen_inst_n18) );
  AOI22_X1 i_data_even_addr_gen_inst_U23 ( .A1(i_data_even_addr_gen_inst_N28), 
        .A2(i_data_even_addr_gen_inst_n33), .B1(i_data_even_addr_gen_inst_N18), 
        .B2(i_data_even_addr_gen_inst_n34), .ZN(i_data_even_addr_gen_inst_n35)
         );
  INV_X1 i_data_even_addr_gen_inst_U22 ( .A(i_data_even_addr_gen_inst_n35), 
        .ZN(i_data_even_addr_gen_inst_n8) );
  OR2_X1 i_data_even_addr_gen_inst_U21 ( .A1(int_c_i_en_even), .A2(
        int_en_ofmaps_ptr), .ZN(i_data_even_addr_gen_inst_N40) );
  INV_X1 i_data_even_addr_gen_inst_U20 ( .A(int_c_i_en_even), .ZN(
        i_data_even_addr_gen_inst_n27) );
  NOR2_X1 i_data_even_addr_gen_inst_U19 ( .A1(i_data_even_addr_gen_inst_n27), 
        .A2(int_en_ofmaps_ptr), .ZN(i_data_even_addr_gen_inst_n34) );
  NOR2_X1 i_data_even_addr_gen_inst_U18 ( .A1(int_c_i_en_even), .A2(
        int_en_ofmaps_ptr), .ZN(i_data_even_addr_gen_inst_n33) );
  INV_X1 i_data_even_addr_gen_inst_U16 ( .A(n59), .ZN(
        i_data_even_addr_gen_inst_n28) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_8_ ( .D(
        i_data_even_addr_gen_inst_n8), .CK(i_data_even_addr_gen_inst_net2803), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_8_) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_7_ ( .D(
        i_data_even_addr_gen_inst_n18), .CK(i_data_even_addr_gen_inst_net2803), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_7_) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_6_ ( .D(
        i_data_even_addr_gen_inst_n20), .CK(i_data_even_addr_gen_inst_net2803), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_6_) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_5_ ( .D(
        i_data_even_addr_gen_inst_n21), .CK(i_data_even_addr_gen_inst_net2803), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_5_) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_4_ ( .D(
        i_data_even_addr_gen_inst_n22), .CK(i_data_even_addr_gen_inst_net2803), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_4_) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_3_ ( .D(
        i_data_even_addr_gen_inst_n23), .CK(i_data_even_addr_gen_inst_net2803), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_3_) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_2_ ( .D(
        i_data_even_addr_gen_inst_n24), .CK(i_data_even_addr_gen_inst_net2803), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_2_) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_1_ ( .D(
        i_data_even_addr_gen_inst_n25), .CK(i_data_even_addr_gen_inst_net2803), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_1_) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_0_ ( .D(
        i_data_even_addr_gen_inst_n26), .CK(i_data_even_addr_gen_inst_net2803), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_0_) );
  DFFR_X1 i_data_even_addr_gen_inst_int_base_addr_reg_9_ ( .D(
        i_data_even_addr_gen_inst_n7), .CK(i_data_even_addr_gen_inst_net2803), 
        .RN(i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_base_addr_9_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_9_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n28), .SE(i_data_even_addr_gen_inst_N64), 
        .CK(i_data_even_addr_gen_inst_net2809), .RN(
        i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_9_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_8_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n28), .SE(i_data_even_addr_gen_inst_N63), 
        .CK(i_data_even_addr_gen_inst_net2809), .RN(
        i_data_even_addr_gen_inst_n5), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_8_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_7_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n28), .SE(i_data_even_addr_gen_inst_N62), 
        .CK(i_data_even_addr_gen_inst_net2809), .RN(
        i_data_even_addr_gen_inst_n6), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_7_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_6_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n28), .SE(i_data_even_addr_gen_inst_N61), 
        .CK(i_data_even_addr_gen_inst_net2809), .RN(
        i_data_even_addr_gen_inst_n6), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_6_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_5_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n28), .SE(i_data_even_addr_gen_inst_N60), 
        .CK(i_data_even_addr_gen_inst_net2809), .RN(
        i_data_even_addr_gen_inst_n6), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_5_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_4_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n28), .SE(i_data_even_addr_gen_inst_N59), 
        .CK(i_data_even_addr_gen_inst_net2809), .RN(
        i_data_even_addr_gen_inst_n6), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_4_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_3_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n28), .SE(i_data_even_addr_gen_inst_N58), 
        .CK(i_data_even_addr_gen_inst_net2809), .RN(
        i_data_even_addr_gen_inst_n6), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_3_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_2_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n28), .SE(i_data_even_addr_gen_inst_N57), 
        .CK(i_data_even_addr_gen_inst_net2809), .RN(
        i_data_even_addr_gen_inst_n6), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_2_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_1_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n28), .SE(i_data_even_addr_gen_inst_N56), 
        .CK(i_data_even_addr_gen_inst_net2809), .RN(
        i_data_even_addr_gen_inst_n6), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_1_) );
  SDFFR_X1 i_data_even_addr_gen_inst_int_offs_addr_reg_0_ ( .D(1'b0), .SI(
        i_data_even_addr_gen_inst_n28), .SE(i_data_even_addr_gen_inst_N55), 
        .CK(i_data_even_addr_gen_inst_net2809), .RN(
        i_data_even_addr_gen_inst_n6), .Q(
        i_data_even_addr_gen_inst_int_offs_addr_0_) );
  CLKGATETST_X1 i_data_even_addr_gen_inst_clk_gate_int_base_addr_reg_latch ( 
        .CK(ck), .E(i_data_even_addr_gen_inst_N40), .SE(1'b0), .GCK(
        i_data_even_addr_gen_inst_net2803) );
  CLKGATETST_X1 i_data_even_addr_gen_inst_clk_gate_int_offs_addr_reg_latch ( 
        .CK(ck), .E(i_data_even_addr_gen_inst_N65), .SE(1'b0), .GCK(
        i_data_even_addr_gen_inst_net2809) );
  XOR2_X1 i_data_even_addr_gen_inst_add_61_U2 ( .A(1'b1), .B(
        i_data_even_addr_gen_inst_int_offs_addr_0_), .Z(
        i_data_even_addr_gen_inst_N55) );
  AND2_X1 i_data_even_addr_gen_inst_add_61_U1 ( .A1(1'b1), .A2(
        i_data_even_addr_gen_inst_int_offs_addr_0_), .ZN(
        i_data_even_addr_gen_inst_add_61_n1) );
  FA_X1 i_data_even_addr_gen_inst_add_61_U1_1 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_1_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_61_n1), .CO(
        i_data_even_addr_gen_inst_add_61_carry[2]), .S(
        i_data_even_addr_gen_inst_N56) );
  FA_X1 i_data_even_addr_gen_inst_add_61_U1_2 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_2_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_61_carry[2]), .CO(
        i_data_even_addr_gen_inst_add_61_carry[3]), .S(
        i_data_even_addr_gen_inst_N57) );
  FA_X1 i_data_even_addr_gen_inst_add_61_U1_3 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_3_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_61_carry[3]), .CO(
        i_data_even_addr_gen_inst_add_61_carry[4]), .S(
        i_data_even_addr_gen_inst_N58) );
  FA_X1 i_data_even_addr_gen_inst_add_61_U1_4 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_4_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_61_carry[4]), .CO(
        i_data_even_addr_gen_inst_add_61_carry[5]), .S(
        i_data_even_addr_gen_inst_N59) );
  FA_X1 i_data_even_addr_gen_inst_add_61_U1_5 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_5_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_61_carry[5]), .CO(
        i_data_even_addr_gen_inst_add_61_carry[6]), .S(
        i_data_even_addr_gen_inst_N60) );
  FA_X1 i_data_even_addr_gen_inst_add_61_U1_6 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_6_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_61_carry[6]), .CO(
        i_data_even_addr_gen_inst_add_61_carry[7]), .S(
        i_data_even_addr_gen_inst_N61) );
  FA_X1 i_data_even_addr_gen_inst_add_61_U1_7 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_7_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_61_carry[7]), .CO(
        i_data_even_addr_gen_inst_add_61_carry[8]), .S(
        i_data_even_addr_gen_inst_N62) );
  FA_X1 i_data_even_addr_gen_inst_add_61_U1_8 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_8_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_61_carry[8]), .CO(
        i_data_even_addr_gen_inst_add_61_carry[9]), .S(
        i_data_even_addr_gen_inst_N63) );
  FA_X1 i_data_even_addr_gen_inst_add_61_U1_9 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_9_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_61_carry[9]), .S(
        i_data_even_addr_gen_inst_N64) );
  AND2_X1 i_data_even_addr_gen_inst_add_46_U2 ( .A1(1'b1), .A2(
        i_data_even_addr_gen_inst_int_base_addr_0_), .ZN(
        i_data_even_addr_gen_inst_add_46_n2) );
  XOR2_X1 i_data_even_addr_gen_inst_add_46_U1 ( .A(1'b1), .B(
        i_data_even_addr_gen_inst_int_base_addr_0_), .Z(
        i_data_even_addr_gen_inst_N20) );
  FA_X1 i_data_even_addr_gen_inst_add_46_U1_1 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_1_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_46_n2), .CO(
        i_data_even_addr_gen_inst_add_46_carry[2]), .S(
        i_data_even_addr_gen_inst_N21) );
  FA_X1 i_data_even_addr_gen_inst_add_46_U1_2 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_2_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_46_carry[2]), .CO(
        i_data_even_addr_gen_inst_add_46_carry[3]), .S(
        i_data_even_addr_gen_inst_N22) );
  FA_X1 i_data_even_addr_gen_inst_add_46_U1_3 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_3_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_46_carry[3]), .CO(
        i_data_even_addr_gen_inst_add_46_carry[4]), .S(
        i_data_even_addr_gen_inst_N23) );
  FA_X1 i_data_even_addr_gen_inst_add_46_U1_4 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_4_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_46_carry[4]), .CO(
        i_data_even_addr_gen_inst_add_46_carry[5]), .S(
        i_data_even_addr_gen_inst_N24) );
  FA_X1 i_data_even_addr_gen_inst_add_46_U1_5 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_5_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_46_carry[5]), .CO(
        i_data_even_addr_gen_inst_add_46_carry[6]), .S(
        i_data_even_addr_gen_inst_N25) );
  FA_X1 i_data_even_addr_gen_inst_add_46_U1_6 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_6_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_46_carry[6]), .CO(
        i_data_even_addr_gen_inst_add_46_carry[7]), .S(
        i_data_even_addr_gen_inst_N26) );
  FA_X1 i_data_even_addr_gen_inst_add_46_U1_7 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_7_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_46_carry[7]), .CO(
        i_data_even_addr_gen_inst_add_46_carry[8]), .S(
        i_data_even_addr_gen_inst_N27) );
  FA_X1 i_data_even_addr_gen_inst_add_46_U1_8 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_8_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_46_carry[8]), .CO(
        i_data_even_addr_gen_inst_add_46_carry[9]), .S(
        i_data_even_addr_gen_inst_N28) );
  FA_X1 i_data_even_addr_gen_inst_add_46_U1_9 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_9_), .B(1'b0), .CI(
        i_data_even_addr_gen_inst_add_46_carry[9]), .S(
        i_data_even_addr_gen_inst_N29) );
  AND2_X1 i_data_even_addr_gen_inst_add_44_U2 ( .A1(1'b1), .A2(
        i_data_even_addr[0]), .ZN(i_data_even_addr_gen_inst_add_44_n2) );
  XOR2_X1 i_data_even_addr_gen_inst_add_44_U1 ( .A(1'b1), .B(
        i_data_even_addr[0]), .Z(i_data_even_addr_gen_inst_N10) );
  FA_X1 i_data_even_addr_gen_inst_add_44_U1_1 ( .A(i_data_even_addr[1]), .B(
        1'b0), .CI(i_data_even_addr_gen_inst_add_44_n2), .CO(
        i_data_even_addr_gen_inst_add_44_carry[2]), .S(
        i_data_even_addr_gen_inst_N11) );
  FA_X1 i_data_even_addr_gen_inst_add_44_U1_2 ( .A(i_data_even_addr[2]), .B(
        1'b0), .CI(i_data_even_addr_gen_inst_add_44_carry[2]), .CO(
        i_data_even_addr_gen_inst_add_44_carry[3]), .S(
        i_data_even_addr_gen_inst_N12) );
  FA_X1 i_data_even_addr_gen_inst_add_44_U1_3 ( .A(i_data_even_addr[3]), .B(
        1'b0), .CI(i_data_even_addr_gen_inst_add_44_carry[3]), .CO(
        i_data_even_addr_gen_inst_add_44_carry[4]), .S(
        i_data_even_addr_gen_inst_N13) );
  FA_X1 i_data_even_addr_gen_inst_add_44_U1_4 ( .A(i_data_even_addr[4]), .B(
        1'b0), .CI(i_data_even_addr_gen_inst_add_44_carry[4]), .CO(
        i_data_even_addr_gen_inst_add_44_carry[5]), .S(
        i_data_even_addr_gen_inst_N14) );
  FA_X1 i_data_even_addr_gen_inst_add_44_U1_5 ( .A(i_data_even_addr[5]), .B(
        1'b0), .CI(i_data_even_addr_gen_inst_add_44_carry[5]), .CO(
        i_data_even_addr_gen_inst_add_44_carry[6]), .S(
        i_data_even_addr_gen_inst_N15) );
  FA_X1 i_data_even_addr_gen_inst_add_44_U1_6 ( .A(i_data_even_addr[6]), .B(
        1'b0), .CI(i_data_even_addr_gen_inst_add_44_carry[6]), .CO(
        i_data_even_addr_gen_inst_add_44_carry[7]), .S(
        i_data_even_addr_gen_inst_N16) );
  FA_X1 i_data_even_addr_gen_inst_add_44_U1_7 ( .A(i_data_even_addr[7]), .B(
        1'b0), .CI(i_data_even_addr_gen_inst_add_44_carry[7]), .CO(
        i_data_even_addr_gen_inst_add_44_carry[8]), .S(
        i_data_even_addr_gen_inst_N17) );
  FA_X1 i_data_even_addr_gen_inst_add_44_U1_8 ( .A(i_data_even_addr[8]), .B(
        1'b0), .CI(i_data_even_addr_gen_inst_add_44_carry[8]), .CO(
        i_data_even_addr_gen_inst_add_44_carry[9]), .S(
        i_data_even_addr_gen_inst_N18) );
  FA_X1 i_data_even_addr_gen_inst_add_44_U1_9 ( .A(i_data_even_addr[9]), .B(
        1'b0), .CI(i_data_even_addr_gen_inst_add_44_carry[9]), .S(
        i_data_even_addr_gen_inst_N19) );
  AND2_X1 i_data_even_addr_gen_inst_add_32_U2 ( .A1(
        i_data_even_addr_gen_inst_int_offs_addr_0_), .A2(
        i_data_even_addr_gen_inst_int_base_addr_0_), .ZN(
        i_data_even_addr_gen_inst_add_32_n2) );
  XOR2_X1 i_data_even_addr_gen_inst_add_32_U1 ( .A(
        i_data_even_addr_gen_inst_int_offs_addr_0_), .B(
        i_data_even_addr_gen_inst_int_base_addr_0_), .Z(i_data_even_addr[0])
         );
  FA_X1 i_data_even_addr_gen_inst_add_32_U1_1 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_1_), .B(
        i_data_even_addr_gen_inst_int_offs_addr_1_), .CI(
        i_data_even_addr_gen_inst_add_32_n2), .CO(
        i_data_even_addr_gen_inst_add_32_carry[2]), .S(i_data_even_addr[1]) );
  FA_X1 i_data_even_addr_gen_inst_add_32_U1_2 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_2_), .B(
        i_data_even_addr_gen_inst_int_offs_addr_2_), .CI(
        i_data_even_addr_gen_inst_add_32_carry[2]), .CO(
        i_data_even_addr_gen_inst_add_32_carry[3]), .S(i_data_even_addr[2]) );
  FA_X1 i_data_even_addr_gen_inst_add_32_U1_3 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_3_), .B(
        i_data_even_addr_gen_inst_int_offs_addr_3_), .CI(
        i_data_even_addr_gen_inst_add_32_carry[3]), .CO(
        i_data_even_addr_gen_inst_add_32_carry[4]), .S(i_data_even_addr[3]) );
  FA_X1 i_data_even_addr_gen_inst_add_32_U1_4 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_4_), .B(
        i_data_even_addr_gen_inst_int_offs_addr_4_), .CI(
        i_data_even_addr_gen_inst_add_32_carry[4]), .CO(
        i_data_even_addr_gen_inst_add_32_carry[5]), .S(i_data_even_addr[4]) );
  FA_X1 i_data_even_addr_gen_inst_add_32_U1_5 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_5_), .B(
        i_data_even_addr_gen_inst_int_offs_addr_5_), .CI(
        i_data_even_addr_gen_inst_add_32_carry[5]), .CO(
        i_data_even_addr_gen_inst_add_32_carry[6]), .S(i_data_even_addr[5]) );
  FA_X1 i_data_even_addr_gen_inst_add_32_U1_6 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_6_), .B(
        i_data_even_addr_gen_inst_int_offs_addr_6_), .CI(
        i_data_even_addr_gen_inst_add_32_carry[6]), .CO(
        i_data_even_addr_gen_inst_add_32_carry[7]), .S(i_data_even_addr[6]) );
  FA_X1 i_data_even_addr_gen_inst_add_32_U1_7 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_7_), .B(
        i_data_even_addr_gen_inst_int_offs_addr_7_), .CI(
        i_data_even_addr_gen_inst_add_32_carry[7]), .CO(
        i_data_even_addr_gen_inst_add_32_carry[8]), .S(i_data_even_addr[7]) );
  FA_X1 i_data_even_addr_gen_inst_add_32_U1_8 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_8_), .B(
        i_data_even_addr_gen_inst_int_offs_addr_8_), .CI(
        i_data_even_addr_gen_inst_add_32_carry[8]), .CO(
        i_data_even_addr_gen_inst_add_32_carry[9]), .S(i_data_even_addr[8]) );
  FA_X1 i_data_even_addr_gen_inst_add_32_U1_9 ( .A(
        i_data_even_addr_gen_inst_int_base_addr_9_), .B(
        i_data_even_addr_gen_inst_int_offs_addr_9_), .CI(
        i_data_even_addr_gen_inst_add_32_carry[9]), .S(i_data_even_addr[9]) );
  INV_X1 i_data_odd_addr_gen_inst_U44 ( .A(n46), .ZN(
        i_data_odd_addr_gen_inst_n6) );
  INV_X1 i_data_odd_addr_gen_inst_U43 ( .A(n46), .ZN(
        i_data_odd_addr_gen_inst_n5) );
  AOI22_X1 i_data_odd_addr_gen_inst_U42 ( .A1(i_data_odd_addr_gen_inst_N29), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N19), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n32)
         );
  INV_X1 i_data_odd_addr_gen_inst_U41 ( .A(i_data_odd_addr_gen_inst_n32), .ZN(
        i_data_odd_addr_gen_inst_n7) );
  OR2_X1 i_data_odd_addr_gen_inst_U40 ( .A1(n59), .A2(ctrl_ldh_v_n), .ZN(
        i_data_odd_addr_gen_inst_N65) );
  AOI22_X1 i_data_odd_addr_gen_inst_U39 ( .A1(i_data_odd_addr_gen_inst_N20), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N10), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n43)
         );
  INV_X1 i_data_odd_addr_gen_inst_U38 ( .A(i_data_odd_addr_gen_inst_n43), .ZN(
        i_data_odd_addr_gen_inst_n26) );
  AOI22_X1 i_data_odd_addr_gen_inst_U37 ( .A1(i_data_odd_addr_gen_inst_N21), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N11), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n42)
         );
  INV_X1 i_data_odd_addr_gen_inst_U36 ( .A(i_data_odd_addr_gen_inst_n42), .ZN(
        i_data_odd_addr_gen_inst_n25) );
  AOI22_X1 i_data_odd_addr_gen_inst_U35 ( .A1(i_data_odd_addr_gen_inst_N22), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N12), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n41)
         );
  INV_X1 i_data_odd_addr_gen_inst_U34 ( .A(i_data_odd_addr_gen_inst_n41), .ZN(
        i_data_odd_addr_gen_inst_n24) );
  AOI22_X1 i_data_odd_addr_gen_inst_U33 ( .A1(i_data_odd_addr_gen_inst_N23), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N13), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n40)
         );
  INV_X1 i_data_odd_addr_gen_inst_U32 ( .A(i_data_odd_addr_gen_inst_n40), .ZN(
        i_data_odd_addr_gen_inst_n23) );
  AOI22_X1 i_data_odd_addr_gen_inst_U31 ( .A1(i_data_odd_addr_gen_inst_N24), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N14), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n39)
         );
  INV_X1 i_data_odd_addr_gen_inst_U30 ( .A(i_data_odd_addr_gen_inst_n39), .ZN(
        i_data_odd_addr_gen_inst_n22) );
  AOI22_X1 i_data_odd_addr_gen_inst_U29 ( .A1(i_data_odd_addr_gen_inst_N25), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N15), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n38)
         );
  INV_X1 i_data_odd_addr_gen_inst_U28 ( .A(i_data_odd_addr_gen_inst_n38), .ZN(
        i_data_odd_addr_gen_inst_n21) );
  AOI22_X1 i_data_odd_addr_gen_inst_U27 ( .A1(i_data_odd_addr_gen_inst_N26), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N16), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n37)
         );
  INV_X1 i_data_odd_addr_gen_inst_U26 ( .A(i_data_odd_addr_gen_inst_n37), .ZN(
        i_data_odd_addr_gen_inst_n20) );
  AOI22_X1 i_data_odd_addr_gen_inst_U25 ( .A1(i_data_odd_addr_gen_inst_N27), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N17), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n36)
         );
  INV_X1 i_data_odd_addr_gen_inst_U24 ( .A(i_data_odd_addr_gen_inst_n36), .ZN(
        i_data_odd_addr_gen_inst_n18) );
  AOI22_X1 i_data_odd_addr_gen_inst_U23 ( .A1(i_data_odd_addr_gen_inst_N28), 
        .A2(i_data_odd_addr_gen_inst_n33), .B1(i_data_odd_addr_gen_inst_N18), 
        .B2(i_data_odd_addr_gen_inst_n34), .ZN(i_data_odd_addr_gen_inst_n35)
         );
  INV_X1 i_data_odd_addr_gen_inst_U22 ( .A(i_data_odd_addr_gen_inst_n35), .ZN(
        i_data_odd_addr_gen_inst_n8) );
  OR2_X1 i_data_odd_addr_gen_inst_U21 ( .A1(int_c_i_en_odd), .A2(
        int_en_ofmaps_ptr), .ZN(i_data_odd_addr_gen_inst_N40) );
  INV_X1 i_data_odd_addr_gen_inst_U20 ( .A(int_c_i_en_odd), .ZN(
        i_data_odd_addr_gen_inst_n27) );
  NOR2_X1 i_data_odd_addr_gen_inst_U19 ( .A1(i_data_odd_addr_gen_inst_n27), 
        .A2(int_en_ofmaps_ptr), .ZN(i_data_odd_addr_gen_inst_n34) );
  NOR2_X1 i_data_odd_addr_gen_inst_U18 ( .A1(int_c_i_en_odd), .A2(
        int_en_ofmaps_ptr), .ZN(i_data_odd_addr_gen_inst_n33) );
  INV_X1 i_data_odd_addr_gen_inst_U16 ( .A(n59), .ZN(
        i_data_odd_addr_gen_inst_n28) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_8_ ( .D(
        i_data_odd_addr_gen_inst_n8), .CK(i_data_odd_addr_gen_inst_net2780), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_8_) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_7_ ( .D(
        i_data_odd_addr_gen_inst_n18), .CK(i_data_odd_addr_gen_inst_net2780), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_7_) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_6_ ( .D(
        i_data_odd_addr_gen_inst_n20), .CK(i_data_odd_addr_gen_inst_net2780), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_6_) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_5_ ( .D(
        i_data_odd_addr_gen_inst_n21), .CK(i_data_odd_addr_gen_inst_net2780), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_5_) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_4_ ( .D(
        i_data_odd_addr_gen_inst_n22), .CK(i_data_odd_addr_gen_inst_net2780), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_4_) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_3_ ( .D(
        i_data_odd_addr_gen_inst_n23), .CK(i_data_odd_addr_gen_inst_net2780), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_3_) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_2_ ( .D(
        i_data_odd_addr_gen_inst_n24), .CK(i_data_odd_addr_gen_inst_net2780), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_2_) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_1_ ( .D(
        i_data_odd_addr_gen_inst_n25), .CK(i_data_odd_addr_gen_inst_net2780), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_1_) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_0_ ( .D(
        i_data_odd_addr_gen_inst_n26), .CK(i_data_odd_addr_gen_inst_net2780), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_0_) );
  DFFR_X1 i_data_odd_addr_gen_inst_int_base_addr_reg_9_ ( .D(
        i_data_odd_addr_gen_inst_n7), .CK(i_data_odd_addr_gen_inst_net2780), 
        .RN(i_data_odd_addr_gen_inst_n5), .Q(
        i_data_odd_addr_gen_inst_int_base_addr_9_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_9_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n28), .SE(i_data_odd_addr_gen_inst_N64), .CK(
        i_data_odd_addr_gen_inst_net2786), .RN(i_data_odd_addr_gen_inst_n5), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_9_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_8_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n28), .SE(i_data_odd_addr_gen_inst_N63), .CK(
        i_data_odd_addr_gen_inst_net2786), .RN(i_data_odd_addr_gen_inst_n5), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_8_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_7_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n28), .SE(i_data_odd_addr_gen_inst_N62), .CK(
        i_data_odd_addr_gen_inst_net2786), .RN(i_data_odd_addr_gen_inst_n6), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_7_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_6_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n28), .SE(i_data_odd_addr_gen_inst_N61), .CK(
        i_data_odd_addr_gen_inst_net2786), .RN(i_data_odd_addr_gen_inst_n6), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_6_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_5_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n28), .SE(i_data_odd_addr_gen_inst_N60), .CK(
        i_data_odd_addr_gen_inst_net2786), .RN(i_data_odd_addr_gen_inst_n6), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_5_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_4_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n28), .SE(i_data_odd_addr_gen_inst_N59), .CK(
        i_data_odd_addr_gen_inst_net2786), .RN(i_data_odd_addr_gen_inst_n6), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_4_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_3_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n28), .SE(i_data_odd_addr_gen_inst_N58), .CK(
        i_data_odd_addr_gen_inst_net2786), .RN(i_data_odd_addr_gen_inst_n6), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_3_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_2_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n28), .SE(i_data_odd_addr_gen_inst_N57), .CK(
        i_data_odd_addr_gen_inst_net2786), .RN(i_data_odd_addr_gen_inst_n6), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_2_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_1_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n28), .SE(i_data_odd_addr_gen_inst_N56), .CK(
        i_data_odd_addr_gen_inst_net2786), .RN(i_data_odd_addr_gen_inst_n6), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_1_) );
  SDFFR_X1 i_data_odd_addr_gen_inst_int_offs_addr_reg_0_ ( .D(1'b0), .SI(
        i_data_odd_addr_gen_inst_n28), .SE(i_data_odd_addr_gen_inst_N55), .CK(
        i_data_odd_addr_gen_inst_net2786), .RN(i_data_odd_addr_gen_inst_n6), 
        .Q(i_data_odd_addr_gen_inst_int_offs_addr_0_) );
  CLKGATETST_X1 i_data_odd_addr_gen_inst_clk_gate_int_base_addr_reg_latch ( 
        .CK(ck), .E(i_data_odd_addr_gen_inst_N40), .SE(1'b0), .GCK(
        i_data_odd_addr_gen_inst_net2780) );
  CLKGATETST_X1 i_data_odd_addr_gen_inst_clk_gate_int_offs_addr_reg_latch ( 
        .CK(ck), .E(i_data_odd_addr_gen_inst_N65), .SE(1'b0), .GCK(
        i_data_odd_addr_gen_inst_net2786) );
  XOR2_X1 i_data_odd_addr_gen_inst_add_61_U2 ( .A(1'b1), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_0_), .Z(
        i_data_odd_addr_gen_inst_N55) );
  AND2_X1 i_data_odd_addr_gen_inst_add_61_U1 ( .A1(1'b1), .A2(
        i_data_odd_addr_gen_inst_int_offs_addr_0_), .ZN(
        i_data_odd_addr_gen_inst_add_61_n1) );
  FA_X1 i_data_odd_addr_gen_inst_add_61_U1_1 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_1_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_61_n1), .CO(
        i_data_odd_addr_gen_inst_add_61_carry[2]), .S(
        i_data_odd_addr_gen_inst_N56) );
  FA_X1 i_data_odd_addr_gen_inst_add_61_U1_2 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_2_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_61_carry[2]), .CO(
        i_data_odd_addr_gen_inst_add_61_carry[3]), .S(
        i_data_odd_addr_gen_inst_N57) );
  FA_X1 i_data_odd_addr_gen_inst_add_61_U1_3 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_3_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_61_carry[3]), .CO(
        i_data_odd_addr_gen_inst_add_61_carry[4]), .S(
        i_data_odd_addr_gen_inst_N58) );
  FA_X1 i_data_odd_addr_gen_inst_add_61_U1_4 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_4_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_61_carry[4]), .CO(
        i_data_odd_addr_gen_inst_add_61_carry[5]), .S(
        i_data_odd_addr_gen_inst_N59) );
  FA_X1 i_data_odd_addr_gen_inst_add_61_U1_5 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_5_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_61_carry[5]), .CO(
        i_data_odd_addr_gen_inst_add_61_carry[6]), .S(
        i_data_odd_addr_gen_inst_N60) );
  FA_X1 i_data_odd_addr_gen_inst_add_61_U1_6 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_6_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_61_carry[6]), .CO(
        i_data_odd_addr_gen_inst_add_61_carry[7]), .S(
        i_data_odd_addr_gen_inst_N61) );
  FA_X1 i_data_odd_addr_gen_inst_add_61_U1_7 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_7_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_61_carry[7]), .CO(
        i_data_odd_addr_gen_inst_add_61_carry[8]), .S(
        i_data_odd_addr_gen_inst_N62) );
  FA_X1 i_data_odd_addr_gen_inst_add_61_U1_8 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_8_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_61_carry[8]), .CO(
        i_data_odd_addr_gen_inst_add_61_carry[9]), .S(
        i_data_odd_addr_gen_inst_N63) );
  FA_X1 i_data_odd_addr_gen_inst_add_61_U1_9 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_9_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_61_carry[9]), .S(
        i_data_odd_addr_gen_inst_N64) );
  AND2_X1 i_data_odd_addr_gen_inst_add_46_U2 ( .A1(1'b1), .A2(
        i_data_odd_addr_gen_inst_int_base_addr_0_), .ZN(
        i_data_odd_addr_gen_inst_add_46_n2) );
  XOR2_X1 i_data_odd_addr_gen_inst_add_46_U1 ( .A(1'b1), .B(
        i_data_odd_addr_gen_inst_int_base_addr_0_), .Z(
        i_data_odd_addr_gen_inst_N20) );
  FA_X1 i_data_odd_addr_gen_inst_add_46_U1_1 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_1_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_46_n2), .CO(
        i_data_odd_addr_gen_inst_add_46_carry[2]), .S(
        i_data_odd_addr_gen_inst_N21) );
  FA_X1 i_data_odd_addr_gen_inst_add_46_U1_2 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_2_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_46_carry[2]), .CO(
        i_data_odd_addr_gen_inst_add_46_carry[3]), .S(
        i_data_odd_addr_gen_inst_N22) );
  FA_X1 i_data_odd_addr_gen_inst_add_46_U1_3 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_3_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_46_carry[3]), .CO(
        i_data_odd_addr_gen_inst_add_46_carry[4]), .S(
        i_data_odd_addr_gen_inst_N23) );
  FA_X1 i_data_odd_addr_gen_inst_add_46_U1_4 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_4_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_46_carry[4]), .CO(
        i_data_odd_addr_gen_inst_add_46_carry[5]), .S(
        i_data_odd_addr_gen_inst_N24) );
  FA_X1 i_data_odd_addr_gen_inst_add_46_U1_5 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_5_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_46_carry[5]), .CO(
        i_data_odd_addr_gen_inst_add_46_carry[6]), .S(
        i_data_odd_addr_gen_inst_N25) );
  FA_X1 i_data_odd_addr_gen_inst_add_46_U1_6 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_6_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_46_carry[6]), .CO(
        i_data_odd_addr_gen_inst_add_46_carry[7]), .S(
        i_data_odd_addr_gen_inst_N26) );
  FA_X1 i_data_odd_addr_gen_inst_add_46_U1_7 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_7_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_46_carry[7]), .CO(
        i_data_odd_addr_gen_inst_add_46_carry[8]), .S(
        i_data_odd_addr_gen_inst_N27) );
  FA_X1 i_data_odd_addr_gen_inst_add_46_U1_8 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_8_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_46_carry[8]), .CO(
        i_data_odd_addr_gen_inst_add_46_carry[9]), .S(
        i_data_odd_addr_gen_inst_N28) );
  FA_X1 i_data_odd_addr_gen_inst_add_46_U1_9 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_9_), .B(1'b0), .CI(
        i_data_odd_addr_gen_inst_add_46_carry[9]), .S(
        i_data_odd_addr_gen_inst_N29) );
  AND2_X1 i_data_odd_addr_gen_inst_add_44_U2 ( .A1(1'b1), .A2(
        i_data_odd_addr[0]), .ZN(i_data_odd_addr_gen_inst_add_44_n2) );
  XOR2_X1 i_data_odd_addr_gen_inst_add_44_U1 ( .A(1'b1), .B(i_data_odd_addr[0]), .Z(i_data_odd_addr_gen_inst_N10) );
  FA_X1 i_data_odd_addr_gen_inst_add_44_U1_1 ( .A(i_data_odd_addr[1]), .B(1'b0), .CI(i_data_odd_addr_gen_inst_add_44_n2), .CO(
        i_data_odd_addr_gen_inst_add_44_carry[2]), .S(
        i_data_odd_addr_gen_inst_N11) );
  FA_X1 i_data_odd_addr_gen_inst_add_44_U1_2 ( .A(i_data_odd_addr[2]), .B(1'b0), .CI(i_data_odd_addr_gen_inst_add_44_carry[2]), .CO(
        i_data_odd_addr_gen_inst_add_44_carry[3]), .S(
        i_data_odd_addr_gen_inst_N12) );
  FA_X1 i_data_odd_addr_gen_inst_add_44_U1_3 ( .A(i_data_odd_addr[3]), .B(1'b0), .CI(i_data_odd_addr_gen_inst_add_44_carry[3]), .CO(
        i_data_odd_addr_gen_inst_add_44_carry[4]), .S(
        i_data_odd_addr_gen_inst_N13) );
  FA_X1 i_data_odd_addr_gen_inst_add_44_U1_4 ( .A(i_data_odd_addr[4]), .B(1'b0), .CI(i_data_odd_addr_gen_inst_add_44_carry[4]), .CO(
        i_data_odd_addr_gen_inst_add_44_carry[5]), .S(
        i_data_odd_addr_gen_inst_N14) );
  FA_X1 i_data_odd_addr_gen_inst_add_44_U1_5 ( .A(i_data_odd_addr[5]), .B(1'b0), .CI(i_data_odd_addr_gen_inst_add_44_carry[5]), .CO(
        i_data_odd_addr_gen_inst_add_44_carry[6]), .S(
        i_data_odd_addr_gen_inst_N15) );
  FA_X1 i_data_odd_addr_gen_inst_add_44_U1_6 ( .A(i_data_odd_addr[6]), .B(1'b0), .CI(i_data_odd_addr_gen_inst_add_44_carry[6]), .CO(
        i_data_odd_addr_gen_inst_add_44_carry[7]), .S(
        i_data_odd_addr_gen_inst_N16) );
  FA_X1 i_data_odd_addr_gen_inst_add_44_U1_7 ( .A(i_data_odd_addr[7]), .B(1'b0), .CI(i_data_odd_addr_gen_inst_add_44_carry[7]), .CO(
        i_data_odd_addr_gen_inst_add_44_carry[8]), .S(
        i_data_odd_addr_gen_inst_N17) );
  FA_X1 i_data_odd_addr_gen_inst_add_44_U1_8 ( .A(i_data_odd_addr[8]), .B(1'b0), .CI(i_data_odd_addr_gen_inst_add_44_carry[8]), .CO(
        i_data_odd_addr_gen_inst_add_44_carry[9]), .S(
        i_data_odd_addr_gen_inst_N18) );
  FA_X1 i_data_odd_addr_gen_inst_add_44_U1_9 ( .A(i_data_odd_addr[9]), .B(1'b0), .CI(i_data_odd_addr_gen_inst_add_44_carry[9]), .S(
        i_data_odd_addr_gen_inst_N19) );
  AND2_X1 i_data_odd_addr_gen_inst_add_32_U2 ( .A1(
        i_data_odd_addr_gen_inst_int_offs_addr_0_), .A2(
        i_data_odd_addr_gen_inst_int_base_addr_0_), .ZN(
        i_data_odd_addr_gen_inst_add_32_n2) );
  XOR2_X1 i_data_odd_addr_gen_inst_add_32_U1 ( .A(
        i_data_odd_addr_gen_inst_int_offs_addr_0_), .B(
        i_data_odd_addr_gen_inst_int_base_addr_0_), .Z(i_data_odd_addr[0]) );
  FA_X1 i_data_odd_addr_gen_inst_add_32_U1_1 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_1_), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_1_), .CI(
        i_data_odd_addr_gen_inst_add_32_n2), .CO(
        i_data_odd_addr_gen_inst_add_32_carry[2]), .S(i_data_odd_addr[1]) );
  FA_X1 i_data_odd_addr_gen_inst_add_32_U1_2 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_2_), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_2_), .CI(
        i_data_odd_addr_gen_inst_add_32_carry[2]), .CO(
        i_data_odd_addr_gen_inst_add_32_carry[3]), .S(i_data_odd_addr[2]) );
  FA_X1 i_data_odd_addr_gen_inst_add_32_U1_3 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_3_), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_3_), .CI(
        i_data_odd_addr_gen_inst_add_32_carry[3]), .CO(
        i_data_odd_addr_gen_inst_add_32_carry[4]), .S(i_data_odd_addr[3]) );
  FA_X1 i_data_odd_addr_gen_inst_add_32_U1_4 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_4_), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_4_), .CI(
        i_data_odd_addr_gen_inst_add_32_carry[4]), .CO(
        i_data_odd_addr_gen_inst_add_32_carry[5]), .S(i_data_odd_addr[4]) );
  FA_X1 i_data_odd_addr_gen_inst_add_32_U1_5 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_5_), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_5_), .CI(
        i_data_odd_addr_gen_inst_add_32_carry[5]), .CO(
        i_data_odd_addr_gen_inst_add_32_carry[6]), .S(i_data_odd_addr[5]) );
  FA_X1 i_data_odd_addr_gen_inst_add_32_U1_6 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_6_), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_6_), .CI(
        i_data_odd_addr_gen_inst_add_32_carry[6]), .CO(
        i_data_odd_addr_gen_inst_add_32_carry[7]), .S(i_data_odd_addr[6]) );
  FA_X1 i_data_odd_addr_gen_inst_add_32_U1_7 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_7_), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_7_), .CI(
        i_data_odd_addr_gen_inst_add_32_carry[7]), .CO(
        i_data_odd_addr_gen_inst_add_32_carry[8]), .S(i_data_odd_addr[7]) );
  FA_X1 i_data_odd_addr_gen_inst_add_32_U1_8 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_8_), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_8_), .CI(
        i_data_odd_addr_gen_inst_add_32_carry[8]), .CO(
        i_data_odd_addr_gen_inst_add_32_carry[9]), .S(i_data_odd_addr[8]) );
  FA_X1 i_data_odd_addr_gen_inst_add_32_U1_9 ( .A(
        i_data_odd_addr_gen_inst_int_base_addr_9_), .B(
        i_data_odd_addr_gen_inst_int_offs_addr_9_), .CI(
        i_data_odd_addr_gen_inst_add_32_carry[9]), .S(i_data_odd_addr[9]) );
  CLKGATETST_X1 clk_gate_int_q_tc_reg_latch ( .CK(ck), .E(s_tc_res), .SE(1'b0), 
        .GCK(net2747) );
  CLKGATETST_X1 clk_gate_int_o_data_odd_offs_addr_reg_latch ( .CK(ck), .E(N123), .SE(1'b0), .GCK(net2753) );
  CLKGATETST_X1 clk_gate_int_o_data_even_base_addr_reg_latch ( .CK(ck), .E(
        N124), .SE(1'b0), .GCK(net2758) );
  CLKGATETST_X1 clk_gate_int_o_data_even_offs_addr_reg_latch ( .CK(ck), .E(
        N125), .SE(1'b0), .GCK(net2763) );
  XOR2_X1 add_554_U2 ( .A(int_o_data_odd_offs_addr[0]), .B(
        int_o_data_odd_base_addr[0]), .Z(o_data_odd_addr[0]) );
  AND2_X1 add_554_U1 ( .A1(int_o_data_odd_offs_addr[0]), .A2(
        int_o_data_odd_base_addr[0]), .ZN(add_554_n1) );
  FA_X1 add_554_U1_1 ( .A(int_o_data_odd_base_addr[1]), .B(
        int_o_data_odd_offs_addr[1]), .CI(add_554_n1), .CO(add_554_carry[2]), 
        .S(o_data_odd_addr[1]) );
  FA_X1 add_554_U1_2 ( .A(int_o_data_odd_base_addr[2]), .B(
        int_o_data_odd_offs_addr[2]), .CI(add_554_carry[2]), .CO(
        add_554_carry[3]), .S(o_data_odd_addr[2]) );
  FA_X1 add_554_U1_3 ( .A(int_o_data_odd_base_addr[3]), .B(
        int_o_data_odd_offs_addr[3]), .CI(add_554_carry[3]), .CO(
        add_554_carry[4]), .S(o_data_odd_addr[3]) );
  FA_X1 add_554_U1_4 ( .A(int_o_data_odd_base_addr[4]), .B(
        int_o_data_odd_offs_addr[4]), .CI(add_554_carry[4]), .CO(
        add_554_carry[5]), .S(o_data_odd_addr[4]) );
  FA_X1 add_554_U1_5 ( .A(int_o_data_odd_base_addr[5]), .B(
        int_o_data_odd_offs_addr[5]), .CI(add_554_carry[5]), .CO(
        add_554_carry[6]), .S(o_data_odd_addr[5]) );
  FA_X1 add_554_U1_6 ( .A(int_o_data_odd_base_addr[6]), .B(
        int_o_data_odd_offs_addr[6]), .CI(add_554_carry[6]), .CO(
        add_554_carry[7]), .S(o_data_odd_addr[6]) );
  FA_X1 add_554_U1_7 ( .A(int_o_data_odd_base_addr[7]), .B(
        int_o_data_odd_offs_addr[7]), .CI(add_554_carry[7]), .CO(
        add_554_carry[8]), .S(o_data_odd_addr[7]) );
  FA_X1 add_554_U1_8 ( .A(int_o_data_odd_base_addr[8]), .B(
        int_o_data_odd_offs_addr[8]), .CI(add_554_carry[8]), .CO(
        add_554_carry[9]), .S(o_data_odd_addr[8]) );
  FA_X1 add_554_U1_9 ( .A(int_o_data_odd_base_addr[9]), .B(
        int_o_data_odd_offs_addr[9]), .CI(add_554_carry[9]), .S(
        o_data_odd_addr[9]) );
  XOR2_X1 add_553_U2 ( .A(int_o_data_even_offs_addr[0]), .B(
        int_o_data_even_base_addr[0]), .Z(o_data_even_addr[0]) );
  AND2_X1 add_553_U1 ( .A1(int_o_data_even_offs_addr[0]), .A2(
        int_o_data_even_base_addr[0]), .ZN(add_553_n1) );
  FA_X1 add_553_U1_1 ( .A(int_o_data_even_base_addr[1]), .B(
        int_o_data_even_offs_addr[1]), .CI(add_553_n1), .CO(add_553_carry[2]), 
        .S(o_data_even_addr[1]) );
  FA_X1 add_553_U1_2 ( .A(int_o_data_even_base_addr[2]), .B(
        int_o_data_even_offs_addr[2]), .CI(add_553_carry[2]), .CO(
        add_553_carry[3]), .S(o_data_even_addr[2]) );
  FA_X1 add_553_U1_3 ( .A(int_o_data_even_base_addr[3]), .B(
        int_o_data_even_offs_addr[3]), .CI(add_553_carry[3]), .CO(
        add_553_carry[4]), .S(o_data_even_addr[3]) );
  FA_X1 add_553_U1_4 ( .A(int_o_data_even_base_addr[4]), .B(
        int_o_data_even_offs_addr[4]), .CI(add_553_carry[4]), .CO(
        add_553_carry[5]), .S(o_data_even_addr[4]) );
  FA_X1 add_553_U1_5 ( .A(int_o_data_even_base_addr[5]), .B(
        int_o_data_even_offs_addr[5]), .CI(add_553_carry[5]), .CO(
        add_553_carry[6]), .S(o_data_even_addr[5]) );
  FA_X1 add_553_U1_6 ( .A(int_o_data_even_base_addr[6]), .B(
        int_o_data_even_offs_addr[6]), .CI(add_553_carry[6]), .CO(
        add_553_carry[7]), .S(o_data_even_addr[6]) );
  FA_X1 add_553_U1_7 ( .A(int_o_data_even_base_addr[7]), .B(
        int_o_data_even_offs_addr[7]), .CI(add_553_carry[7]), .CO(
        add_553_carry[8]), .S(o_data_even_addr[7]) );
  FA_X1 add_553_U1_8 ( .A(int_o_data_even_base_addr[8]), .B(
        int_o_data_even_offs_addr[8]), .CI(add_553_carry[8]), .CO(
        add_553_carry[9]), .S(o_data_even_addr[8]) );
  FA_X1 add_553_U1_9 ( .A(int_o_data_even_base_addr[9]), .B(
        int_o_data_even_offs_addr[9]), .CI(add_553_carry[9]), .S(
        o_data_even_addr[9]) );
  XOR2_X1 add_539_U2 ( .A(add_539_carry[9]), .B(int_o_data_odd_base_addr[9]), 
        .Z(N59) );
  INV_X1 add_539_U1 ( .A(int_o_data_odd_base_addr[0]), .ZN(N50) );
  HA_X1 add_539_U1_1_1 ( .A(int_o_data_odd_base_addr[1]), .B(
        int_o_data_odd_base_addr[0]), .CO(add_539_carry[2]), .S(N51) );
  HA_X1 add_539_U1_1_2 ( .A(int_o_data_odd_base_addr[2]), .B(add_539_carry[2]), 
        .CO(add_539_carry[3]), .S(N52) );
  HA_X1 add_539_U1_1_3 ( .A(int_o_data_odd_base_addr[3]), .B(add_539_carry[3]), 
        .CO(add_539_carry[4]), .S(N53) );
  HA_X1 add_539_U1_1_4 ( .A(int_o_data_odd_base_addr[4]), .B(add_539_carry[4]), 
        .CO(add_539_carry[5]), .S(N54) );
  HA_X1 add_539_U1_1_5 ( .A(int_o_data_odd_base_addr[5]), .B(add_539_carry[5]), 
        .CO(add_539_carry[6]), .S(N55) );
  HA_X1 add_539_U1_1_6 ( .A(int_o_data_odd_base_addr[6]), .B(add_539_carry[6]), 
        .CO(add_539_carry[7]), .S(N56) );
  HA_X1 add_539_U1_1_7 ( .A(int_o_data_odd_base_addr[7]), .B(add_539_carry[7]), 
        .CO(add_539_carry[8]), .S(N57) );
  HA_X1 add_539_U1_1_8 ( .A(int_o_data_odd_base_addr[8]), .B(add_539_carry[8]), 
        .CO(add_539_carry[9]), .S(N58) );
  XOR2_X1 add_538_U2 ( .A(add_538_carry[9]), .B(int_o_data_even_base_addr[9]), 
        .Z(N49) );
  INV_X1 add_538_U1 ( .A(int_o_data_even_base_addr[0]), .ZN(N40) );
  HA_X1 add_538_U1_1_1 ( .A(int_o_data_even_base_addr[1]), .B(
        int_o_data_even_base_addr[0]), .CO(add_538_carry[2]), .S(N41) );
  HA_X1 add_538_U1_1_2 ( .A(int_o_data_even_base_addr[2]), .B(add_538_carry[2]), .CO(add_538_carry[3]), .S(N42) );
  HA_X1 add_538_U1_1_3 ( .A(int_o_data_even_base_addr[3]), .B(add_538_carry[3]), .CO(add_538_carry[4]), .S(N43) );
  HA_X1 add_538_U1_1_4 ( .A(int_o_data_even_base_addr[4]), .B(add_538_carry[4]), .CO(add_538_carry[5]), .S(N44) );
  HA_X1 add_538_U1_1_5 ( .A(int_o_data_even_base_addr[5]), .B(add_538_carry[5]), .CO(add_538_carry[6]), .S(N45) );
  HA_X1 add_538_U1_1_6 ( .A(int_o_data_even_base_addr[6]), .B(add_538_carry[6]), .CO(add_538_carry[7]), .S(N46) );
  HA_X1 add_538_U1_1_7 ( .A(int_o_data_even_base_addr[7]), .B(add_538_carry[7]), .CO(add_538_carry[8]), .S(N47) );
  HA_X1 add_538_U1_1_8 ( .A(int_o_data_even_base_addr[8]), .B(add_538_carry[8]), .CO(add_538_carry[9]), .S(N48) );
endmodule

